PK   �i;Y�K�e�5  E�    cirkitFile.json�}[��6��_I�_v�T�x�����x���m7z\FB
I���ʨ������_Jq�T��8��E�,��`�2D����!yί������a�Zw?w�������0w��u�K���������a�z�i]�p�����b�O]�X}��z�6eU���u]_�Y��E����e���}�ÏwW��W]��P����/ݺX���i��k]xY�B�N�(�BUVW���6�C�z��z����?B��[+��S���S��U����������!�Gͬo����L�	&���?�����L����Z�WB��o��_��.�����,�^�EӊrfNӆӴb5�D�d�^2Q/��WL�+&�w�D�ʡ^�z!D���m����0J��wz�+�`��s�'5��p�r�6���i�j�g��\/�ժp�	=e\��a�N.���2^q�f�p��4�YM�\ӽ.E^*��|U4�*��5�+Si�µ�H�XM+NӞ�tn4S^8�Z[�w�^H��D��k����6�G9M3��:7$�X�a�9�k���s�a��9��n�s�a�����4L�&���?�ğe��2�g���L�Y&�,��?�ğc��1���sL�9&���d��1����L�y&�<��?�ğ��� ʫ�T=�}��+�n�:�M�6T��i�����ߐXa��H��q�0��a�Դ�j�RB܌q��s�v������cp�r�#��8M��2ѽ�i��4��WP=[��s�W���t��Au�2��y_�N5F�9�+թ�h�b�%el��0�)B�]���.z�C��V�Q8�u�*�L+���h��A����t��*!-��,�Bߘ���0G�a9�r�5����k�l�+�wQ�h�4��]i�^I۹a���ۤ�YC�`���q��&r#:	'9|Sp�;��Z��o��w��O��q�a�5��L什�z�
ozWh��L��bs�5a�_.�B��A!7Q��X��P�:EPa0Κ�en�#��3�=�$B��4oC�:�Pa4͚�dn�R�oˮ�5]�;ӄeW���a�_V����!$U�+��d-˳7��Pa4͚d�ؖbl^�f�$	Pa�y(e�?�3�(��s�R��UYBzj�}\���^Tm��^d7ehЄ�VQz�`��Ec�fL��U���|��(�� 3FӬM�b�]����;'��3#)��,�*��)߯)�J��A��V�gīWWMր��S����\sz�5I��I���q7�FR�\k:�5�.(�j:i�W��tvAs�]Cj�?�R���sy�^�3c��Ή�tn�B\�s��9��JN�9q��Yjd�����א��<�Iݬ��mV��%��M���0S5�8&��`sU#ت�j`�����/X`#囐C؏+���'����/������ڏ+���'���/��+\a����'��	�|ې<�k��4�~\�V>��o���p����ڏ+���'����=�+�b�g����'��	�|qt�7a?w,�M�3=W5���g��&lg0�V%s�鱽���Fa��A�	D��(��x��3=W5����p�;�������{v7��#��у  �rB���N'��	�v����nh�y`�[DQ�EL�׻@�`�� ;��"
��,b"��Z{���Q�E`�&/�:�%��(��,� ���y���)vI�E`X�D����K	��E�E`X�D�����L�A���aE`!�/�:�[$�>�Q�E`��/�Y ulL�A�*�}7XX�D8����H��-� �(�"&�����@�96R.]b�"&  W��w��n�(�=?��`�郗`�[;"�= �#	�I�ǈ-� �(�"�2<0��I�ǈ-� �(�"&�e���1b~�`v6��#��у ��l�`g�;��"
��,b"��Z;�$���Q�E`��I�8����1�Z1�;|W�X�;����B�1��	ν��j�/Jք��n˶h�Ţ��Vt��Eu"2,�z62l��PO����a��E��ȅn�V�V�c�Zξާ��MPEc;sM��0F�9m��oc�C����q�f&i������4!�jP�*
BET~�{&3P���w�pLԴ� ����P�0���^�����Wh�!����`X`@,0(�K��A�ĠX�(��I����u2K�%��b�A� X����X��E�GM�z�U�w���$'G�T�����h��F�(v�H���ŦW�Ȱ�d��_��i�j��M�=o:��m�h8dv(vm���IN�y��B�=H�!�YQ��X���33h�X�1c�ƌ�3�Xl0c�����.6̊�`Pl0(6[�-��b�A�Š�bPl1(�[�-��b�A�à�aP�0(v;���b�A�à�cP�1(�{�=��,���BT�ډ�:�������?����?��F��F���D�d���QԼ���BMOy�MB�4y�KBMyڟ@��xڝ@M�x�aC��x�_CM�x�%A͕x�#AM{x��S�~e����nO��W��hF��[ʪ�eC����8]�R��P#����'����/Tj{�T��7�lI"���/Ԉ���9=\j�P#�v }��x	� By�P#���W��x{��j{��j{�Դ�gj�=g�"��93�3�Y��>ߠ��9����9�j��z���9}�E�*sZ/Ԍ0��#��.g �<-g�FĔ+�y�fO9=�S���n�9MN�o��$�'j���#85i��!����4/�T)^.�ʑ��9R?�F�׋�m ���n���^d���SZ$t��Nh����Nhi��q*8U��3n~~~8U��AB�I?�T��Μ��3���-:N�
�t氌�3Nhi��q"8U��3����"p�@K���S���-��8��C��:v�\�Zc�k'�X:s���v��>~Ɏ�� ��"p�@Kg�����4H�8�*�ss�Ei30�:ʞr���d	��d��ƹʮ�+����-����:����f@�<Y��a>��ȝ�D�7�m%���E��9��܉�% {ÜgQz<Y��a���ȝ�n�7̅%��E��E��܉<( {�iQ�<Y��a���ȝȘ�7̝%��E��Q��܉�* {ÜjQ<Y��a~��ȝ���7̵%,��E��]��܉|-��*0�Z��Oye�_��܉�. {��kQ<Y��a���ȝ��7�Bڕn��~&�a	J�D�<Y��a��(�	�$�t��0�ZBn4Y��a��(
�,��0��U�N���_�Ҧ��"��]E�D���a��(K
h<��%w";�,��0�Z�OOio��*r'�ɀ��E�W�d����׮"w"���0�Z�-4�_��J�D�<٬�߼Z%�9�B����t�j&��Q�*�,�cP� ����BE��慚4���k��M��	P���ͺ~�0GM�§"!T���P1*B�A�x�
�:x1��
~��`����`X`@,0(�K��A�ĠXbP,1(�K�%��b�A� X��+��
�b�A� XaP�1(�k�5hE�A�ƠXcP�1(�k���b�A���؀6v���b�A�Š�bPl1(�[�-�?�A�Š�bPl1(v;���b�A�à؁�l;���b�A�Ǡ�cP�1(�gQLN�§r�N�(|*g�DN�§r�F�(|*gmDN�r�
9
��Y��	P�T΢�� �O�,��	P�T��n�(|*g�6z zϟ"�� �` |��� @���H�(�Q���H�( 2�?E�'@�����)=
���O��	P d@K��(�&@�S9�j>��z!'@�S9�r>��z!'@�S9�j>��Rj>��/j>��P����P��dx�,J� 
���F0@h�:� M&t�[���-:� Mh��TH���
�4H�D4U��3�)@4U��AB'���-������-:� Mh�+� Mhi�Љ(h�@Kg�e�(h�@K��N$@ASZ:��$@ASZ$t"
�*���3 
�*�� �	P�T��� ���-:� M�9�9��D p�H�	�Ov�S	P0�ƹʮ�+����-����:����D8Y��a>��ȝJ���7�m'��E��9��ܩ({Ügq"8Y��a���ȝJ���7̅'��E��E��ܩ({�iq"8Y��a���ȝJ���7̝'��E��Q��ܩ({Üjq"8Y��a~��ȝJ���7̵'��E��]��ܩ(��*0�Z�Nye�_��ܩ({��kq"8Y��a���ȝJ���7�Bڕn�]�J�Nڕ.�]ǿ�{ۄH�'��7̿v�S	P0�����D p�H{��kW�;� co�-N'��7̿v�S	P0�����D p�H{��kW�;� co�-N'��7̿v�S	P0�����D p�H{��kW�;� co�-N'��7̿v�S	Pd߼Z�&@�S9���� �O���@k�(|*o%��.����q�~X��}'���/�u����^t����a�n���~`��#��w��,Y�ʴLLZ�8�h�ța�l��JI�N>	b�5VӆѴ�5]1�V<f2QC��������L�*b�9��3�1B�i�h��&�����9�p� I��AD�� 1}23�Ö�`���EYMg�b8�L�Đ�P�Y��Z�1�f@��ɰ���t"yjuF��	�Z��v�k�����G��h;���Vg���j������ս��TYmst.x:�K��%g8ϯ"��mgW������řKTv.!�>d�<5b�DF�<��\۴���s ��u�mh�
�v/bHF��*�9��t�s�M2�ήӈ1*Mg�i����ь�Jˬ��4Y�xn�M���ۇҜ��sZ]N˹��h�9u�b<��Ӽ����,Vh� D��8�$�a��đtB�}�WLg�%1���M����qN��>�~�ڇ��M�����bw?��`�ߝd����9B����K��U�=�p�<�p�<� �y�������`�) ��a�I�ș �#�� �#�	!'܃B R�� �ǆ'9�"���9�����,��H��d�����������������z����(��D���$���$��1%��i�I>ˡ%���%�K2�00O2O�g>ǁ&������8��s�=�<���8��s�=��̣O���<=����|��#_N���p��1�E�8�s>>}������O��&��U�>;N��u��|Z=<o�Mw�������6���e{��׋��>0����Y_1�A{��'�,:"ǁ�eJ��=�~�E�\|
.@�c�v�%�����Pp�(�H�\$J�H�E��"QƃeιI=M��e�h��8�\�J.N%���S�ũbO�\��Ĥ���J���*��m��7X�~���Q���r�����"y3�pꭥ�^愃����8G��y"{�io�D�X[��8βw����;�����;�k�8n����;��8n�+_���(���D�E��"�r�h�H�\$Z.-���D�E��"�r��Ht\$:.���D�E�c;��Ht\$:.=���D�E��"�s��O �t���H�O؀x��!ޏ�zC�7�#r�6�:|D�w��!^���ev��k����h�P����%�;�����'>+�n�o��������z��) >š:
��#ݱ��ŝ^2�F�X�}����*���7��u�?�<y����7��;�"�<y����W&�k�O��m�D�`�_��q&���O�D�`ɛ���R&�K�D�`�͌豞�$���f��n�'��w���ݭ��9r�Rȝ�>oiQO]���"r��	ee�$r'�E�PF=�#^ً�eV�ԅ�yy�C{.A^&��>P�#���.r�O�k���M|l@��/�� u�&^˧rG�c����"�;2���"��6�Gb��X���DL�Ƚ�=T�	=��"
��,b�^�q�V��3��Q�E`���k=�����"[DQ�Eܾ`j=�苣�"[DQ�E�>�`j=�Ӌ��"[DQ�EL�����(�.�ĊlXD1�.��jb�(��t3u��7*[b�X�3���a�M=�c���T��"�Gb���4��Fiq�@"xFeK,��Xb�� ��9~i�h�G�4 �~b��1�E���������>�����G{��ėR��h)S��/P=�$�� ��-�@K�z����!�v	�h)Z�Tp�T��	�c�/�@K)�R��T\�z�wH��C|)ZJ��22�գ}D�2 )ZJ��2���c%S�[�A`)Z�T �T��	��D �h)Z�TL�.`="S��k �XJ��2^�գ�>���K)�R
���H_��C[F���w���"�����@q6~����|y�1����Ę��h��D{��R
��-�.2!W�h��D{��R
��-e**$?e��`<���D��@���D�$�h'_J��R��L�N�@�h'�D;��R
��-e*�-?	��0���ߧ�_`i�)��`��o����fR�'��R_c��ҟ�C����a't'�����1�L����n_�,�!�D��<�����}����� �Й�;8	��������rX;�At��7c��q;zƈZc�1>��i\m���6>����g���#��i���r|(9�Ho��H�����%���|���cn�1=�j�)��,�cb=�롆j衆j���j����j���j���jء�jء�jء��4԰C;԰C7�pC7�pC7�pC7�v��n��~��~������?!�Wޘ?;SkJ���v�C ���� !:A,H�Hy���HyD�Zq`��}R���|R���{Z�� {R��Fz�aҙTpF�N���!hI���:m
�j��J1��0X�0�G���~���9+��t5�T�4��֗�l�i����ꚦ��r:����-:�Y���j?�#��v �6�8����$��Y�hsň�0�� B��cfd�Zr �5�Nq�c��?^����w�Pt,���E���qkh�cn,�^lȘ��)��g���I'��X��D;317";pӈ\΍Mp���I4.��%�aݚg�'����о�Ę��PM�=h��ˍ�Ġ��]21V�k���f"���a�՚�9�7V�M�"8����jb�i�	Rĝ̍��к�+�,g�馆#eTf-�rA�hnN�z(�X��i��a>�Y�yqN9�uV��\�M����pb���5�v�b�ȴ(�h��$��5����pH$K�]y�BI2�cb�,�+-Z$JF/KY9��"�dp��=��1&���^K�VZ�@��a��3���EȌ%ɭҨ!�/�$wG�I��+:Z�fޓ�s/�]6Ђ-��;��T�����Ŝ?���lC���bΝ�\��J�}��X��@n!Ƽ���oߜvl��o�{����}w��ns3����}�'��$�Oj�Iş�?��'��O6��v�\���>��S��TE��^"V�8�#և��C�
{��X#b��D�U"b���ND��W���"�Z�Z�^-"֋��E�z�{��X/�X/r��E��"c�Ƚ^d��׋��"�z��^�^/2֋��E�zQ{��X/j��E���b��C����zQ�^�^/���׏�o�m-������y3I��V1o��~�������0�]��a|{��zSr��?}�^}�֛e7^����i��a@�>o�˧�������׻۟�Ǘᯯ��WG^��������_���M�{�������[�u��l��o��?_�뮽}�	�U~��^�z�yYw�S�-���u��|Z8	��)y�Y��~��ޙW���L��u������6P��t�[%mvg*��(}]�]K+D�+݈���%�ڭ�ǖ�����yS?-��H���nW�e�Ro��f����c����w��-�ŝ��w?���9�Q�?h9���r��ʸ�!3_��rOL��W�G\���V�wG������}�e����jZC�YfZc�Y᧿K��P��)���kI�|�������#���$��|��.OI}_M~Jr�.	�.+"Y.��t���r�H/2y�X��t���r1���⾐,w�d��'&�)���'�vZ�g PHA,���8(3�+��̉�	f�U�VN�)A�Qu���О)�ŌY�i�#RYM�%K�jJ�J�r��%��$Z�DK�h���	�)����e��&ђ;A���@G{1K2�V�b)�F��h�K���J�5.�Bk\*�ָT
�q�Z�RI�ƥRh�K���J�5.�Bk\*�֨T�q�Z�R)�ƥb��;�v������cۭ�~}?�|�߾{���n��������imk�pAuѫ�Kh¿�آt�p�l�˱|��O���e�����o�u˦��J��-|5\IX���ϲ��J���'U( LWXׇ-h�芪n�fG4��ƙ��z�>}zټ��e��-�V�n8���8�����څ�[��}�s7��C����n�U�o>,�7��T�^�Da{��,��jS��i�N�F6b��o��z��ӧ��-awgt�RW�[jj�������mmT�y\=wo���]آ�'���ˠam�Z-��}/���S��vC�a~���������g�4R�����y��c�S=�~[�{�����j���m������owa!�]�|����SJj݅���]��v*��۶q��!�+�j]U,�`qݛ*�D�B�F6�΋´��I]}cB=������mU�����+[���Ά�Nx��+��e��_t�>�������?����s�y��?��ͯ��?���˿܄�n��zYo���o>t���f��Y�<ݬ��](������W�4����)Af�}��M�>��-�-��w��b3bf������v;|����]փ1,J�� ��[n�߼����)q+�ս
�I8��~#�}���~�o¬gt��ݢ���$�	vl��n4EU���bQ�M�hٓ�$�wE7�6fwF�������~��^�ݟ~��7��|��=�	R��k�:��ņ�zJ�o�B[u_�0/��4t���N��s��zk�FԲ׍)D%�(ۺv8�/�.�ε�ْGz�E�o�2�(�uW%�T&2p���@��Z�-���R[�����	}�R�ۯ��Z�:L��Ą9Dy[4��a�����E[鎤k�38���\:Ai�@}��8no�X9|�Ã�R�_��P�rv��ΑaM�t�|��M���{�|X�
�-W���kg�.T�a���XJz�}I����'V%KYq_�R�)�R���2t�W\M�k��Of���1�rw?T.���>Z��B�
��54�)̽��U��~,g���}����[刻"���B�Wn� lY��|-�J�(���z=d l��a�v^ʽ�ֻє>`_�U��+"�~�UaL��fks{J�C�d�R�0xaw�ϕn���alE��\�u�;��2�����rU�b)�Գ�H3��+�e��
���ہ���u�<j,l��Nz3Z�
���q�$h�B\���A
5H�5;rV�raf�*f��V�70#��
 �R����_���{k���)����{�K3&��n�L���َ~Y��C��s�2J��+P�Y�	L��]�4J�[��^�@qK�Q�
��w�i��ЕB������3��1� q{h7��a���p���f���J���R^4]�:z���)�p2>��҇o��������M�D���*̝ڝN��R��1}�t�[4E�ȶpu���ʅ�a��e��E[�fL�{kʲr8"Vp���ە��O�;�&t����.���Lܛ}�@��@C -�4&@S�&�%m_�)�f����/LY��K��*,��*�!��<��3c^q�����͋�S��\�)���H;�m����Q��M3qOsTU/l]�q�jMX��U�ac`����}�<�0)�i�+��.!L$��D9.*�%}y\��j�;�ﵺ��U�J��@Q�8>�՚<�J�t�N`�V����uY{���WP*)"A��h��F�n�d�a����c�@�Lx����t&�Q3�������i�h�T.���j���Ʃv�9�?�1�yuBU&��a�"��!hʩ���Yc����p̹�9ߩ*ttj���/��5ou�Y?\&�E�ƆoX!M��Ţ���]eڦ���(q(���B�֕��nSh�_.Z�������������SȿN֜Ѻvc���O�o~��\�N����������?����ޝ�6��o?�W/O�7���ۅ�+3�e^����;-�k�?}�S�S��K�'����~}���/��_=m�_�W��z��ʣ=K-K�k߬^��7�~9�^�k�T�²�i}�ª<�@�W^��m&ӂ6�ndQ��*Z1l'�0�[��a#�,i'*�U�;����jJ��w�_�u�~Ynn�}j_�:A�洐�x¸s��Luu�Z�bQ�ɩ��U��.l�H'{e�xFؐR��Q�o9�`ܲ�[�������~�ۭ�՝+��KQ]e�#�X#MpGw<�]�n����Mv���6�U����9�}ީN;u/�7Z���a|��{%t�~�(��W��H��4�]�5����1,�?{�?{���2l�\i��B|����ߗ�˰���g�W韤����9���1���*��6���a1��Ǯ����F��e��0���r��n�Ӈ͸_T�~��0����u�1m �{Q/>t�����[w��?���~��`����߯�Ŵ���f�W�ލ����֡>��]Su{��=I�bu$����Z��o8�>��aܪ7FZ����vxc��������P�<��������͒|(q�,&3�&Ϗ�żJS�]P̹t����\L������O�[ua�!�+p��`�
(p�E���&��=.�A����Z̉\�)"�bi	_}�;M�)l�	��(� ��,�0��E�83�%J��[�P�V��G�4t~���;:�j�	k00t�5��gw.t�f�tHs�ugJ@A%Ey!&f�
�D�ۙ��^�}x�;1�q��	Z)��ǜ4pʰ�r4Q���������:3|\��LhLG}m�sô�*��^��z��;��$0��3����en,>40�,I.bo&0�8��B�U��_j�������B�a�4����95!͍�Fϙ�"���8�L��F��rŐ^�T�B��s(�j�ڕ���e�@�U�^���]�Z,(3�tB�IP3r��;&�Z(7Uʑ�.��"8��b��1� �RP1u��
�IԮC��7C.D��p'\C�-��c��qP��K��)���WZ��d����^_F�^�T�-tƒ8�8�%��q�X�2e�R6=��ߺr��cXnPqmc��P8`x40��,AƴTv�J[	O=/�Г��t��cG�w�u�]v3xE�q�Ν�&+�1-�V�8��M/��R��#Z22,t䅇G3xEB'�.:C��[M�z�R�I˞+����}�
r֒4w/-�x֒dw��fBC�Z����Q�
?]2�J�{�G��Tn�Sw�}����i��� "��g�7@��9*���gu�_'�b@%Ʃc E�� ZH��z躙6��3����h{�]��մT�ywi*Q,7l����;�澣��D[�쾛��\�W$��ʜY=.����b���=�^��������*�]їsUr>��R2��=��J#��u���b.Y��CJvJG��(����n�I෇C�7w�Ivr1��ᕵ�U�x�ꋡ������h�_��AP�*��2h?;���c1�Dj&018��H꼭fY�M��9�O;�� �i��� �w���}���fY~��Zj��pM���x�J��N���r�e��s��a�C���D?��!���r�E��X�@㢛2�,E��4�-��5��[�G�3����Eg�gM5����:D(���ǁC�wȯh��ؽh�|�T3�~�N-[�K��H��#Gߗ�j��ڤBrO������=��g��~g�m�{�~<.&��3l;��R�#_ 4Z�U!s���٧8�g r\���{"8D���^}��C\vc�~���\���@�+	��cW �2'�9Sͱ�6q�>��i!��I�A�5���L�a�q�á3��[|�؅\l���+�
� �_�3.�����?k�9v���!�b;	|���[�}��.ڻ�5����H:���b�<J�
x����
{��.:�=k�9v�FR�����̴�>/�I��ܩ��U�'b��!muBI����'3؛����
��k��	��yTh{�"b9��5���*��I�\8_I3��\H�ɫ���.���!�(D!I}�t��H�-�I���&��g�7��r�%zI�ńJ#D�#�-���]�>��7���H���!i{WC���!�b¨{g�R�p���	xY�ࢡ������P�Ѷl��e�I��c����O�����O�x2"�́�4S�<1F�%+���㌶�m�H���y�w3؛?��IC���x̚��1�V'0�3NCceJ��[J�?� #ɗog�7���9�P��%�R�V���2����\��R���Wj�o�(���.�7ot��z')�s���R��%2;u��8���v9��?�����`o�GQ����W{�'/`��
�x�L+�;tu��1D����3mNx/K�v�u����Yj��Г�~\,�""&�<��]؞�Ԟ��'^ۣtu�������͎#�Ӧ�߯L��ƥ҇�cq�evR�^�x�h��ޕP�En>;�u�EńNO-G("#ޫ��P�ץ��*J�|�����\T��B��ye*}r��^\�Q��+��~�ݹc�d�'�G�t���+�� �Iѧ6��|iҚ�1��Y��r��J��$��t&��Q^�k$�\/�zvnH�����a��vr�xo����/&f�
�D�۹o�e�0��dǣDT
0J��%܅��V��Hp;�2J���$Fǣ1e^��꒔b��&�����O�5)���W�)៦�d��u��<ҔB�(�v�Uu�h�`Ѯ���3<�������(��Q���_����`���B+�NSd�>�R��p�����Po���~|�}7��y�c�_]����~���㷛���l~Z��o���k��X/?��������f��f�=���f��i���_6��c����o77�O���͢n�O��]���7�S���/��7����f�y��=�7?������y�v�7��Z\~���i�C��,7n^��Ao�:4�ؼԁ�����9p�q��n���z�xwӼl6����[NV��ˠ�0���,77?/�_}�n���,ƛ]c�?����f����o�PK   �i;Y��(� � /   images/0add2520-d67e-4490-80cf-da78ad043e6f.png\�eP@�5�C��$���{p�����n�=��-x ��y�{��}�GwWuU��s����Vu����G��000hr���00p�00��(H�f
v���eu�``X���`��D<�MR�ɪ+���������<���``<�������g���;%K���H�I�iz���z���xܽi-@��Wi�b����d�iL�%?s�"�����>�>z�:�n/���=h��?��Uo�����&̳����������|�E����쁭���񚡡��۔OB%S��v��$'b��l^���=0w|<���	M[8;��x�
��s4noXY_U�Wpq�'��}	E�]/B.���H���;z.[�h����:�=ް9������k����*��L@��ז�g��g�pFX oi"Ǔ�\?��q�;x}��$C!������S��0��N�!��l��%q�EG��g|g��:N�?-������IN�P5[
������M��Y�C����jZ��K4��y�r���<iCҩ�E�g�N���͏B�&�[��F��H:ފqGQMoO�E��.�/qz�x庼ֵ����Q(9���Zu�K�?��cމ|��OR�Z��榛�}<6��}���r9N�F�8���Y�azZd%�.�qF�L��W)j���N������������Q�㸋��s�{ħ�Y�����zh� ���q����p)��T$X/f=))5ߢ5ܮ4��|r$�����!8��sA��f��
�ZW*�i��A�ɖp�)���q�~��ida3w%3�$��o�q������;��;Fz�WQu%�B��S�&{��W�)����������:��Ĥ:]G"[��!������8�����c}�y��3��{�A.y.;�֓�=���E.����6�)0�:w�lt�.��T�g�s׿^������ƶ}\����ɫ��:�$Y�	��WGO�z�?���B���C��(.{�x�S�(¿Rgx��Cumא��������^Hd�b�?p���^�&�z���:3�X1��	6���U���\ꄨ� �5���ս��<]�soxle��m�vS>5�c��Ԣ�Ds��0rm�]�^�����ʲ��%������49#A�RJK�a��J�A���Ď}�='Э�<�1W��j=r��YxIdq�2��y4����fA����-�������&�)�&b��2�j(�Â��C��:�K:lk[$��1w�	����˝ZQO��9���[�S�p��Ƞ�c{�}���$��FFe��$l~F��d<_F���'Z8*�o�硭A��[���Q�m�A�V��7��Vu����P���Vmk�u	.)����0pf�e�V.ť�����a�O�Tx1��B[������D_s���u��FȊ+d�q�"W<����WЭ��ۆ����h���>Ibm��J�+ߎ���N��&ۯr_OS��)��~���)�T��U��{������/Z�L�C���	��[T�	,����O��P������Z�[���E��^k"�I���8U5䘓N���v�o���xC�0��%z�w-O�F����\k-+�@�'KI�x��B�/8�/9��޳�eN��|n�5oI0u�%&�t?��5[?�dն��YU��+����[T�q"|<�]8���>�%�Gp���KF��������W�WS���U����2��y�N�'[���E�K�.��:��*�[%��1X5@�yҘ$A
���@��؜�P�x+z ��j��+�nyyzk�O�����f�~j҉��M���c���۠Gt���U�_��"P\�g�K>�0(N�j z)@�N��XL��#@l^��(����3G��Ȧ}G��bC��Ij3Z��0K��pLw �4l��K*Q(h�����Ɉc����??���.�M��fzV���t���<�٩Q���>���Dʼ�%�Uy
yu���lVYЕ�k$����#kv'�8䇜��ε���Q��P��}e�����?�i���M�}]h%�wEOgQ:�e�F���J��|�-L�#�a��yqq�fx%�z$閵f֕	�1����x瑍�����k�
/���1b��QAg�u.�Q���$��������������_�l�]�5�7`�������/�֪�_�%�?�FP0�i���P2qְƸ�Hׇ�)�]�x�7y�g�gp�w����,t��F��=ݠw��{dm�U	��D�d���h֌�肖N����"��I a���Ri��{J����(d�
x<�7+�>s�d�W����@U4R�e�_��GBbêD�Zy6G,Dzb�ϻ���	�Fqa�RI7�`�a]�%7����>�\�=��D����)-v���Y�d,����8��=������t�<���%�_� U]#����JY�p:�6qu�!��Mw�5>�W�2y�;P��l`O̢6Qܔtb�	��^'�~M��Z|9���l�*AAF�u��QN��oC���h���,��p�2����aw>ȩ�1HdQ���)m�d�g��h��ɤ�ſFZ3�F��%�.sz���v:��!�Q)v��}͂�q�����b��r�ߑ�'�`(8Nzb]�=�K�U�ܞ�"�����ѻ@���	���S[',/�4F�D�.o���97%��JW�)�3��}]��hz� �8�& ��YLK�L2�n9,��p9N�>�I�)�?m��[�~R���
_�Z4�Q��������{b*�`�A�G�ձ"�.�I�2�,���n5� ����*��E��(�����s�� � ��{Jc��)�a5��
[/�k��h��:e��Evl�*̇o��u\��]��)T����+���d_�r�|�+u���%��+�~���&W	�������X�^�l�-�(g%Œ�o�&�I�\���Ԃ�,��21K�ک��r����Z3@�F?�����l��c�����k��O_�����5L�q���g��zN%�mJ��M泲)�>��/+o!az
7!�(���E7��u�
��#�ٽ�d��97 ��x$���4_��S��D�'�k��y����ɤ��x{�9�?����yD�O[�s��b��kE��	�$gdQ1���_����{��N�����O��c��1w��J�'*v���%Q(�w�`�c������u��<�s�/FZ�'0��⤟�Y��UT�{�`�����0�u䇸Qx���'��V�/��V��b\ɓ2n�Z��$z"���,tp�"(빑�?%g4�w`J7��a���PF��8�;�[�L�ک��=(�.��L�������Bz�t���DC2��f�D�|��^��}�]Òf��|ɎOI-"O�{����/������9��s<�\��ů&?~���ɤ��qk_o�����s��u�rɵ�j�]��"�(|ϟ�/M�(����-_�������t�̀��N�� �.n0�ᎼG�`��V6�ݼǬ߆j��wwj�|w���=]�e�i6�P�r��<G#A�˾�l�H�Ѯ�^L!���䈧��@��`{=�f�{�I�KP���!�JM�f�Ք�f�p����Q�JtN֕[W�[�:R)���=p���d��;	����0�\D{���+פ��
��/�X|ƞ��i�zgTY�Qqzݝ,I�Gr4Aʛ�
���C�o|�~��׿�T��`���pK����d�~o�_'�S�R���]���5�C�N�[�_��f[���c��J��ة�������l�v?�j&Ǟ,rc���N��c{Ap��o��]�e~b`��W(���MN���^��Ay��)A���cc�eQK�0!CL�v���S��X����W��&�`�"��r��zu���]2��Mf�&��&yj�T��8����(�W�A�'�ħo#r'o�pGXM`
২�U�ǭ��l����5^{:�8�Y��W��i�Oe�9F���O[��A�е���	������[����8ԗʳÍ5%�_�v��\��>��~�v��E�&�F*Cl<�e�{ �{���3��5O�aMN	f�5j���������;ve�&����+���h��2ŗ��ԛ�t�
5A�ly�H����M��R�pc��W�[��`r�/��$Pd2�?k9�"{���p����Td���� p"H"f芇��MuZ���["(+!Br9j��x�3t�Mu���jd7��	g=�-f�D"�� $�<�
�q�o��l�� P:"���� �zkYPT�7�_
�}�1r��{V1m�Ǹ�,��/*�x���Yo%�P����9�'̚�)Դ��-I�!o���Ț����k��ߛ�v�N�)5;	�
�ޱ#6��I^���p�I�aJS�9x]�@E�����%�ԧn���~�����X�ӓ��!���񡺫8�����*HC)��-]K�E�����UF�?���vH9)j�X�s%�����lDM��2����$%�t�v.lxadQ��܅BMW+���YŠ席��@��i�'ҫ�E�{m���+�Z�P3�H�2'�<ϳ5��:x"�nj�G�(�h.�_P��~��O̆L&Sa�����6� *�f��;2�����\�,�y�Hp^�V�u:cd�,��AB>%��X���I��U��ǎ�#�*!%`u��G������>���_Sd�H㇞���{�V1.�f(��Z+�V<�(���UKv�����%��)A��Z�i"Z��5�T �7� �g��zf�yZ ��IT�-�H?�����zjD���:�^�_��n�cc�]?�軶�S���տ��9� y�c����b��Xz��0��_�mm�Jk��&�4�ź!�ʜ����6ߨ���%@&Z��Cgzdk���b?%o����_�S����9/?�^�=���HqM��n�G��V�êt��$2M���+g�������ē��9���_�Y{�Ն<s0�sw8�S�ݏ�=��D�H���,���y/�R�b8����M5��b�h�[6���a9����0�e�+�Sݞ�B�9��8��&6��˦O��7W(�N=Vӫ��^u��y!+���DhM���H����nD�X�
`�=b�u~H+���Gܝ��\�+R��H��~�ެ�j�ϛ�?q���p�ښb�"���1�h������R烖��;�`w&�8A�O�wY*��X����Zw�[����
_=���h� 8'$�A�f ��稜J��2!,eI�����  ��u�x�
��8��s̷%�3�m��p�h�oJA���d�5��Ԕ;@��<H[�\��6B����д�X���	"4�A@N|p��'M��J�P}g$���bt�z��&$�JI���8��bC@�z���/��rUAZ.!s�y5:7��1S�����	s$q��YF
>ߏ�F�37���-�f��rv���k:��,�0r�!muȶ��<����"�{8��il*�)��#�����>�I���+���ʬ�(�m�S�Z6<�*v��?w�/;-���*�	¢�*9u��6U�h���L�Qt�����{T!�����&��tNp�5��\�4#J�t x�#QK��Ju���2H����_6��e� ����C�C�����pT�x>���5�H�.��?��#[�0~�JW|-6üozɘM_�:cw��d(�<IK�+�1n%-����AE�є@��Ӗ�)Y���$��<t��)�����A������?�v�g�gg���ʿff��85�j��/���2��υ���KB��j�\��.&�uLM�v�%���r�l�wO:��V��mk#ׂi��-��� +ꛆg�}�M֍儃�ݭ��Lޭ�9F����@�s?��Խ�[��:�tx��ƶ�d>���\���\�[���O��P����$�m�o�a�Ͽ���ߙ�u�b��.\������%�>V��� ��H���ʕ~s@8p�u����#�%! mI�Jz�;������9�nV�D�� HW�Kl������=�]�oT�b��?@*tq�BV�O�U�c�\w�}��UJq��I
"c���*��Ҝ`�d�;���^r��V�����2��
���L��#Cda�H��2�I�m�ʏ��P�/�l�:�EA�޺v�=ހ:��bkK��
3�K���D2�dP�=�m��H��|�cH�N�����:qw}Ȥ$Un�[�_��V���|��6`�ŷ��9Rz��_\ٝ�XV�=�%R��ߠ3�|o&>��/]+˻�D_�ٸz]J-���`=�B3�I�_�ZI��VS	츨��T]�N@{�pED�Y�GeI�$�.ߣrP�z��Y- "ǵ-�;������2Q/�S�*�b܊���6���釴���H]�.�U��0\&A���o+3%�Z˞�x��q�~��Y'ʃ�,q�ާf�
�5Q�V���j �)��&|�/�`��R��]H���b��6�8^-�}��IBf�����#�@)d�|��X75�^�
,P���Δ�ȃ�<�y����uk\{C��+��"�浰��>t��lY�wt�t=#�]ƙ���y;��
_=���ױz]A�"ci�������-m/���)�Þ�#r_�P��6^�U$"��uٗ�����q�k+�cӌAm�\_�C�t�_�t�;�x�0T c�MGf��4O@L^��@3�6�l>�L[��ʄ�p�A�J����܆�٠C�7K������M��˒��{�����}@�R�x������=��/���JF��5�R���#���A��.��Q���\���C��x�y`�ӴmziW�:� D�!�2 �
Ƨ���P:\��R�jp)t�����w2��ꥬ Na��8�����eg:��x��`L�`��U&4+KpSKc�S����Z�z\Oqaͻ��)��*#�4�eQ�d���k��.ˌ�%FM�ۈd&&q����v?�*��T���#c��Ʀ�,|d�f��{b_}���)��"�rH�1-�����*���[ր)$�xX��FMV�IvL|M���^UL��通R�[,�^��}PԴ�� �!�N͛rY���$;�R��I���嶁tbgA�X{i������\� �*"��+��D��#<w���okM<����ŚKJ�ޓ��Y^&���N;1�E�����V�6&b(��Rhƚ�⁮QZk����[�<��"A�����/�����J�����0dJH�R�����(k�8eov����q��6��y�4����\��A2�m�Z�,jH4�09���O�S�ѫ�"��`b�� V���W�4G:+�p�����={�3�� y$�� a`S�����JB�+ �8�Nټ���lm(�`����-d�\;�F� +�#�x�W�B�l5	i�#���{��^b%+q���Xm�՜���a����L½!�%�����Ҍ̕���;他~ـ�VM�A�DN�Z���C}��	��u�f';1Q5���N�U��[��_N����Y�>�$h'�,p*1�g�FKG���x:DW��]�wd%�~Oiͪ��rb�:�L!��:ĐٰG?����$Y$�� Ou���yCj�6����C)�E�b�H��P�89�V�hy4��b~M���ILDv�\j�7}�N߂�@=�SA��JX��@%)os�����`�/B��u&��oXv���z�sA"���0e�}�P�I�v�=p�D�$g:��·˃�ֵSk� ����_�9�^�.�VF����./sR��EW��$�>k�²:���V��>��l�{�lެ�+�lM�jD�G��^n���M�r�ͦ�6�o/-LG�Xg�`��?���),GF-�����2��X�	��ƴsr�7��|���P�̰��0��,I�3�>Mq'x"6Pg�|������3�y�j�b�Z��&Iے j����D�&����Nj��Q2m�m%^���/�?dIX<��*�a�c�����ih��o�Dq���JRQŤ���*aG[K�G�q��j�OG���#�oPk�ku����+�,
�q��0+k� ��lQ���Pi{�;%׃U$m8<J�]�Mb�xkf��2
zF�R'm�����(�@�[��+$ev_QN�2X�j^��O@��ak����pY�[�?�:V�X>�9��!��ŷ�M��OJZz��@��7>�Z���|��ui'����	��:V��(n�t��L#�j������$�9���1���,�JHL��.Ye��."��ɹPGp%hu�3,CZn�I����)��׮������"s؝u�[�G�x�qT�(��'�o���G���C�ZJ&�R;a"e����I��H��;�)>��y��xdM�L1��G�^�'�o�s�	�!s'bGo��[`�lq�ɺ���#-j*q�$m�\�p��5����q#�`k�`�$	YE�Z���Ti�5���H���b{�^ld�j�����k�p����Z8u��oa��*��:��<,g��ݼ�@m~4�A%D��C3L�]-.WH�}hH�O]��<��p�>��hr����ĺ,�e�ކ�fk�4ew2+�\�㔫��6v]���;t�e����6=6<����b5��͓#��m��c���z!��D*)�2��p!�1�f}h|�m�I��!yԮ�m"Q�o��g3LH}ȅx�'���r19S%ͺ�EdKM�GP�J�C�����3
�30׮c����L�i����E�"r�<Y�w{�y�.
܁�M��\.�8%��Zj,�<�P�5)}ZL��b��!X�l�G���
w8�*�ʘŚ��kB[���q����#Q" x�Q�B��2\�������oZ�rI,�,V2c��J�9	��v��a͙)���W `VK�P���w�F����o|(
Ӄ��ېA���ިt���:�f�p���	�J<��"/aȘ8�_�$w�ϔ��*tx��D��q"�w0���h���j��ɳ鼅n��ל��bs���`�U3~�ZR�1��kA�E���2{k2����/��h5MVJE������\�v�9�\-�Vw����t3,���J��L�o��N��+�g&�lw��+SHL�0^���jln�;� ����!Y�!Ӽl��]��(���d�U�����J��6���g�W�
����o�￙I����F��d�3j��U�#��9�Aϯjrs���`oM@1i�n��5wNe&Sߺ���3Va.��˂�)�t�eS<u(�� ��u?ˊ�7���+�O�V�s�=��ͬ�0aT���s�*fE``���	�V9kL^[qor��F'ә��>s�~�:<?n	� g�.�z�i�A��A�i�B-)#:���o��ZX�0Rj�DG-���C��Ǿ&ѩ�0�Ϻ�͘Ia�Џ�z�g9�kDn�v�ˢ7����[Ku���&9�e��z���S��d����=G�7 OkP痐~��w]��Q@a�G��ī���L�m���<`����47X�a&(0�����h%_Pe�)�EX��jE�a{���й:��w.:v>�s���+ͤ6.�<=3���m��?a=�%ǖ r�ۘo���ػ8�s�I��4��MMZMa��`0���E�1���l:�X��T���8s�V!�������������0qt3�M��Zlȥ1��aLfj&5�_���!^"�5�)v��o�
2|a��v�I�ʌgػ��<&[ ������,�eJ�T5�?���f���JK�(�'�l뢕�3�xs���o���,���n�
`C?%�Z�N���O7�3hؾ�Ą�!1�A����w��j�9-ܰd߳����X���#F�H�\M���>��}��K	l��g���u���j"���;�P<4"�l��ɲ�,�����]�v�������s����Q���J���g�d�FJ�i�Mv+�@~��ME���~DT1�Ԩ�Z�ޙ�q2G�R���a���|Re����ԉ��I��x�"5y�4V�Juo�g+.ڢ�JeH�;�t#XS+�q���ʫ�u��vx��Y��Ǳ'���v%�:�Ml<A�v
�C>��qR�R24Ԓ�?�БaQ}��qJ��uTe�1I�N5!�E���}\03���Z�\V�T�,vL{��M�q>X.��xZ{ˉ� ��C�
�V������"#
�j���4��*������s�ym���:����Q/e�������>1�t 
�=�����WD�ȗ1r�t�tXc��8Y�>��xS�R��?�[<��:Oa��Y�|�x�s�\��D~�!��`���r�`��V]�}���Q��=�[��g��^�h��fH��o�k���)֎[HTB�]��((4O[5�8���`��K=��6���Q�/fh�-�.�K�5#d/a�%�	:�D9�^�D�·%���Y5�|�Oa�K���ƾ���`&�;C2�/��\S1���������k�E�j|;�>��G�3g�Z�%A��������"�4q3k�e�,/ª<U��:����29�l2��u�����Y�����>NcT�k��_ح1�~;Ŭ>�?��zZj�i6��R��n[������&�(;��V+�0V��~rs��>
ޝr0�qk��w���
3K=��?eǽ�
�d�ZAeK�w����6L�aA�&�b��~۾�yL�z���FnbWZJ?E����Y�{��=2M����)� Bq�y�˹ooDD���UZ�v��׀e�u�B���� � �Qr��z��A]�/����1�p��m�|f��p�8FF��Y�1��2����m�]-�Qi&C\rC�K�s˔�s4K�l�T�BX����
'�F�>�شB�Uw%¥��(f�Mǆ��0��<��7k,�Ӟ�gf��; ����캶�dg0�䨅h���N��Kyߔ��%ѤtF����h�@x���O��Dk��i��* +��1m2�E�����.{\��C4\�}�G�8;�_1�.��C3a��ԣ{#�;_����k�'�%P�$N7;��b�����?O�q�ğm���xi!�9+:�M���Z�vt�Rf?��2�V��7�����v0bj��dv��U��W��n�Ν$�.8g��h�/��8����+�]��E�+�K'S��q��A���i�~�3��������s��9+	>��`�?�hϞ�+jE�S̘Tj*��ѽe7���z�6�>n�O�Kmu��W������ӂ�n�<P+��>A��Y�o�T3Fa!kw1ɯ(g�C�$��V���������'�fq���M8Z��t��I�j|W*�9q�+���}�Ĩ��,W�S��]��~Ћ3�^�Q�zB��7����l�}U�`������!|����n�w*�8�)�q7ĥ����R��f#)"���Ϸ�-*��F�?��(u�����$��N͆;������'\�d�w���/j�Z1L Z���`�S![4 ����G��'W��/=�Z�����/�9�".��Y���G.���?)�Bo��5L�#g��>��ѐ����N�DT>`4j�%�$�3�"����3�Ă��OqY2�Sq@�$�W��I\�3_bsa	Ԟ�&���;@���v�C C�1��r��m!����HpĽ*e���L���W����<Bث��J:�▴ډy�YJ[R��N�˘]g�=���G����	+�DA���z7�bQ��nGss��ʘ�B0�����}E�h P�޽O��ַ�@2�������x���A�$��A�ܾe���q'�c�Y}i�o��{$��B}�{<�����-뺙B7fE�;ܝ 2��"AS=xl2\��Wi4�,�s�?�N�Ù��[Tk�9��B�����b��y���b�oc�|�Ő�ڵ�	H��\�Eӓ>� �p�Q�I�>-{��/	
��Z�2���7ÎS���FC �[p���b��1�4�/R!���x��*��%�:}����Zƥ񺜄k��:A�G>c:m;��,��fL�q6�f�d�o#feT��r
�1��7�FTr\D�jM�F�wޭ�Y��mB`%pY*\�F��x��)����S�=*��t�Z L��z��e���J���}�3�ĩ���x�M�N���$D�"�;��c��Vgļ���9���K�PtE���`�A�M�B�a=�����{�3��|
�����U��[^�5�A�XH%�^:O�e�&�o2�<�a[��.o֚�wu
JHJQF<��>���!�z����'��ϰ��0Ţ�F>�kMݼ����8��*/�pCܛG�O1�!,�Sǳ��YL�.0���§���rB�+%����Ȏk�&��P�n�tZ��#Y�R��/v.Y��k�������ͳ��"-����������繳�?�ɾ6]��-x�ꃒ<�'/f0��}Éާ��W�e����m	��a� o\��@�£m>�VG��B�C[3���_�o<�$���aU�Jk������̫KR@�AƏ[IB�$6�ݵ�󌠤rD�����ܰ�����q��h	�sD�߿������r��.L`!�`2��E+Կ �=Ԇ�jC2�%��ki�[ˡ�1�äM�|w<YbI=����� �W2>5]�%���jto����r�-g���j��+�����gM�@��W��vb!DNp�X�����P�*~��&�S �����b����U����\7��D�j�|�Upw�_&WL��ԃf<�TR��R��-�AX!�fTh@�ML_6��"�ΐ��ĄZ�9�lAx	cp���)'c\(n���"��a
���%#|-�	��G�e�m�7=�w�MdI��~9��7St������n�*5�_���X��� r�D1"��>&��rG���b���h��2�k
�E	��ݳٹ;���;/*�x��>i�L'��`�cF�������!�~}r�e!Jh�C���.���\Yj���|�y�xCgd�S����ΪԊ�^����OJ�"�������ŋ�8I��>	�K�i��_	б��d��֮Q��*8�ظ��A�Hh8��_D��P��ֶ�n��B���k��g�=�k��:�-jw���/,��=)�~���xc�,�W�
"��7R�#_-� sR���>�ǝ�n�t��7�鑿ސ=/�؂���|+-I���tBm���n�Ӗ��Y	i¤R�B�Ǝ�n5���U���pX�7���1Ζ��۱�0"#"yAi���1o�}F��+"5��W�	_�&6��S�p �<�� �,��Ʀ���mj��fA5{��㨢�� ��ŧ���D;.E��덾���̲_�`���{��{v�,0�d��\�e��(f��CqWw31�7+�&M̺G�ȋ��s�2�!{$�7:�)��[���AEݞ�]�ᏘO�g�����GF��6�/�n��"�0�*�����E��wmY��ٌ�%�,9�I�ț�]�}�wyǹZ�/�������������/��I�q�)MP��_+���T��+ۀ�Oz�vzka?a�j�`���ĲP.���8�w�%C�H�u��^�������'-�}�ނ������0��	ƭ��C�
n��w~��E*�NT&-��;�%��$@�qR"�T�p����̜��O�eN�&�O�|gh���޹�](���n+
�6�G�����q�Ɲ�Pm,ꚢ!�#�d�0�Ȯpl~�u\B°p��§�7�O[�a�LU9;Ƽ��M[������GR����-���O��.c/_{'RtH8WT�v�N�D۫j߸�����O
4+wT��\�Y��vK���6�I�ݜ�8�Ȕ���B8�4wgj��?�'�p�tb	�$Lf���n�.��;����4��ȉ����5���-��Kޘ=��I/��E�LP��Ϸ?Cl=J��������S�:.YV��N
Ik,-;��ҙ?ʉv1�n��b{�kxN˘��5��Īە{��]Sߗ~ ��K�p�i��@t��wO��k�,����S�fJl���D�b��+h���w�/<����	O�Ε��:�Av���{H�K��עJ�"�^��LDrA �NLׁ��Y4���=YD�L��/��B+��-��������i����c�8JuQ����<�5k�>�ft��Q�w������ʊM�Ҧ��Ǜo���~��i����}d���aXY�U��m�B�M(N{U�ҪF��(�]1͜0� |�&���-Y|MF�/0��6�K1� ���Dp͘�P|6i�8�K�&ڤ�t�Zup��8�2�2�'�A�� s���4�hļ���T�c��s�v)�x�S*���x�K�nf���At��y���j?&�	����R�2Rt�K�Q����R^V��<O�l4�Y�T����,�D��3����>5�ii��z�m�"���w)�4hCE���g)��J7
�@���juy���d�O������n��eǺ�K��. �� ?B�Ƨ�Jf��b��J���2"�>m�����F�i��S�D�� I1Rj=}�������;�����i�3EC�t6ƚ�� ';Q<���X�*���ʟ��o��� ���j�l��?��c�B~O<}b�\��D?����h⪷#WZ�D���GSu��x`DвȊ�Vlt_�p.j~2������{�\�ӖNa�����ie���N}1�׶�g9���|g���<2�0g�,fZ5�@��$b��_��%G��	��m�=*w�������i��lI)�$�����F�-�u�y��
?�m?���`h:њ|S�WE��g&k���Kp�
�H�L�ғj=��}�֎=B}�u
�t/�S���;�|�ɝ�A�;�e�V�j�q�	P���t8q�c���P�ǰ�H��a->� �+�IRH��9p��a�<`��`�`11k��*�^dMm��Na���*�X��?Nu.�1I!p`�/t.�o�T���F�3��+����q}J7~R6��������ax3�9pm�6��A������ƍoZ�1#���&5y,G�i�1:v�;������F�,P�����=������nH�!i��q8}?����-}!6�7u�u��xh%�/��$lʂ����"�*e#��Ԗ�h���s���}n��?��Pn�r�.Jֺġ���<q�&6ޒ.��x!Z�ӇdsA�r�dӔ����6}����cw��v�K�g����s��9���U��C=Ogd�)��TzG��?!�[R�U�Q9�ZL4B�c&W��GW��|y�}& �m�OwJ����&D`�B���(Ղ�	b(2��x���y3QYq�]�������X��=	���:�k���@��}���'RPC2КS��d�5ܭ���K�'bo�����F�o�G%5��.�2K
n���V7��\a8���=�N� ��K�����JN��u8��� ꈸ[�YK¬!�#����GO�e�}=�N�����C�x���m��#��y˞y��4ݘsC�i��V���⥯����ZK�6i��Z�� U�RѴ�kn���{Lb,���aRJ�j��YnTU�tE\��ͭ�N��M���U	J�R��)0$�����t��I��������*_8�K7%Ri:[���s��|v�����Rݪ2Z뺓��c��8@e�0��0�p;2��}�����fcD���ˊ>���-��h�ŘG�X2�.�l���n@,��*9@Mh���13�ƿՋJ���5�f��u��ɱ3Sz��K�vy��cj�s��%�!���d}}���D�#(�V��I�Q�6w:��T���dK$_2k~���{]�BBIaJ�_i�mK$f��xY�J��MI�B��.�儤�S]�5B�f��%��DI3��B^M�{^���PB3�eO�΂H�O�u�3�gafe��뼶Y~���Ҳ�c�[@���B�$��Q��g+Ŵ��XB�]S��c���Ҿ��o|�{�=p)���%-�P��`*��x�y�}��5Z�P�\ĉ��`�c�ˠ��Kk�
����r�t�:�Vq�/m<��^�u�Ɖ��jN���¬���]�> n�1
�7�F"H��Ҫ��Ŏ�n>�7=��w�R���f�����,�	���l�1�f�JIv�'��C����~&䫛*�٨�
i��2�U�пd�%�q���q�y�y�����k��{B�o�L�����j>��^1�(Y�'�k9A>�������-���$�b���e0���b�6�a�:�b���,X"��F�I��呻��������!i���� we�kO׳��l!R2@�x�M� Q�i�]����8z���݁v�M$�ʝE3.���U��
�(Rƥٗ�� �@]���CY��8���;���k��!Wߴo3��hP�$��9��1D���t�M���(O��'�%��Fn0�r�y�-@r���}�Y�|	e��:�5�]�=[�b\�9�ǉ���0�kPU?��T��r|_z>��11�\��fU��QNY�TeCd�H�h�o�.$x0��'�r�����+A�@�T�T0I��V�eSCL_T��'rۮ{�c�5�ظ������+�|�M�ne�~�A��G7`�R�=�YO:C�a��꿾�i�T�*tuJ���1C|����Ɨ~rC
E�&��O�ag�J�}�Ob���ʻ�	?hƪ|m���n���97��ϗ�ܖ���;}$G��j�?!U{lۻ��l�nR�G� �c��!�c��MdxH�(�?6���B�s�t��3W�P��-�U��%y�jU�X��p��A��*.J�X��\������y�y��.d�ĄĎV7Q��c��A ���b3
�Dۤ�kn��w.����lE��MU5�4�9���ܔIHj	��55�j.����:����l溛n扏9�g?��,_<����! !e �-æ�k�1Յ7"5�jQ��k�^��o�ߌ7��`3Bǔ�����ex_��lڴ����q���v1A.��1��sǦM�޵�{��e����s|��x����Yc1��m۷�k�N��Y�D�)��Xc���b�R��mK�E��Ae����@,t݉��?7�/'3��W=��P@`ʱ$NM�]�l�8��uU#����<MSF����c;�����NRb1�:�DgbL;�Nͬ���{�l8D�J,|U	�O�8;oM���H�׎]�S�)t�G��i��f�8�?ߩn�Q���$T��P���
e�f���F�Sx���1�v� s��Y9�k�B#���W�g]���A�VrA!�N�l�u��&��o]~?��J֟|"�s�O9��,&�N���o����X��s�8[�6��57������L>�YO�ݩ�{�n�̓�Cc@�/P�+��6���V���eR��w�F��y3�:��;�,��Trgq�謤=�SIK-K4���3�p�&��y#W_>�����.ڈ�L�ҙ�E�h��1�	ch6���/�Ƥ�7Qb����7��Yg���woa׎��!ŕeY������Q�Ji �I���䥴!��t�)<����߾�P	+!Pu�#��B$�bD1�,�UǱ�-4(�X:=f��}������#N��L=�Ɍ���L�[M�����OZ�c+��݄�i��NW�*V��d;���Ƌ2#S����>3��㜬���w����)<������nR��}F�'�~�
�N:��>�;3p-�d5Sg���"���*n�o�%4	���x�mw�e��u�3·�F�m���>�"pm�9F$es�C���LX=���h��\ͱeWo��+o���V-b��E�Z��%K�0<4���K�޳}�v�o+���Ǹ�V;�'f��W������B@���M>�~�=�U��ۻֶP(��K��"D�T	.��F~t�M,np�	k8i�q�j9kV�`dt��((���G��z��;w���-ܻ};{�G�b02ۡ�$�M�<XDʪ�%p���#��?Ǌ�+۳�F�A�m��EA���_C���ɝ%�s|���N��O}�_=#�s���ƒb�]9�;	5:0�;j���O�)��y���	�I�g^��A������-L#�������K�۶m%�b�킘ٯ�L���􃊙��3�W�ⴰq sz@~,V�����'_��0�����q'�̶��\O'�!��t�f@;t��W�&$3��W�B�s���n�K^��w����������9�2Ġ�'�<��&E����*�!j
Q����v@�B@�Lc�@����q5y�'"�����2�H�+YE���di�6�l���8����|�}��2R�wb��F�XLl��?>�b���1�2N$�I���Ynڛm,�����Nr��йD��ꤹ&��%}Y��2�+DTSŞ�ϸ�I�$�����<�Q��ux��c��z��zG����������5U�sw괜Vo�ZH��`�CJ�5�>0<��37<�VYP
���'��'Xى��8���Xu�#���	O��z(�rcd���{e{�ݻ����7u� ;L_$ 6��H̄�=�9�ͻ>X��y)���'���s�U��&��̱lŊǬJ�~�.h�vc��� �<�δhl��N�� �A��X��Bc-����8E(h@�b*-���{�R��ZA���qj��q|lz�������7
V�PXII:���Q�q����'Ϸ`���m��($#����OYczڕ^�^hG�b4`%�gIM� �t@C MmE�n%l�|_�r���f�TRD���&H�o�1ɾe.×%�������;~�(5&!j�@�	�P��;�����5�ip0J�+�����G�fy�k�s�����2�S�G�z� �!_t��]��v��:��ю�vuC;OQ�7�1r���8a�)ؑE��m��:4��f��؜�9¢�g�o'�C�g�Yd�����|�FM��o��Ҥk4��h'��������Px�@x���4?*Z��Ӊ�w�z��Ď��tar8�A��D�(���+_�4��P��\8'���b�ʃ`;��,���w���_��9P�hk�|틟b�qv� ��ގI��Q[�����~i�=c��]�}����K?��� <V��ف�&����0¯������yEʒ�'�<�e�X������^ ������R��x�>�WF�vfl��^0<�g����U_�z�AN�H��~��5�cG�S�h���M�h��Y�h˗/cdd���� �ݽ��(��ORm
C�j��'	�w^�săd4��h������lN�;+=r3�$�'��ų,K�el'piv7=v�k��TTC��1�I��x�0]P�	���P2b=ǉ�=�-H�q{��4cR��N�g����^끜��Hg�X�}h��SUhXȁ���G���f��^vetK����x黁�&�I.�=���4��}��O�E�{���i�����y۷o�,=��؞]�۳���ps���E�}`W��k�Cm��vT����»,4 X�{>��kp<�j?_m�U"�=��Om�����x[:�z˲�!�v�=��]<���t�n��t�Z���Q���b'vT�?yM�	EL�/KO��̺�c�b�"�$��\���
�r��{�&Cg��y��>p�NO^*V�`l����u�#�(&%nʮ�hFk;|�*[��*���T�[r"�"�;�<sE������v��YMN��DRbCԀF('�����|Gg�*ǫ�J���c(8
P����C�t��U�b�vD�θv�����S�=p���očIq�Q g�W�+^��\q��������Ν��K�KjT�R��]�M��t�{;�j�r�����������
�J	oۼ�y��������Ku �U�F���ҙ�d��������M���0�°�1ۛ=���%�@�_ğ��oU�a�l�8����עqh��U��&�{��e�&ڔ��ɰƀ�tQ5*�#�v�w��݅��Hu2���C�}�6K�P1�ū�c)��!�s&����8�V[mG����������>i��Ҥ0M
��a�d���}�$+V3+�N�0X86��Wp�8+�zp���~A1XM��^\W�{I��b��t@��n���Mu����B�L7�l�μ�O6R����A�`\%ń�6�:;P���*�P[m�z�(����K����H �����}�,�,�3/
�����.X����0%bPc����]�D�"��l�k�7k��v��<�\pqq�+!��{�Y��� ���8��M��W�b&o�@Y�~]�I�g2������J�uTj��1�zտ:�QMP5 ����t���!�.�`\6{��t��>�g�����i�%�z� @�H�rR���0(8V�QE���?���|��o��w�ݔEk
��I5�"خ�X� ��g$*Q�<ϧynLw�!b\�)���5G+�G�n�j��.�[m�:�����xa3- ��`�B]�2����t���}�����L�)�\C�g���h��*�s:p��gD;��JF��T���x�s��2�F�MB���7�՞,SWv�t:�z�:k��%QS}�A��yɬ����l������ml�c�2tŹ|d�,���{����o���D̹���6���R��X����Y��W�5N��<z�h�Hw���l�vٔ�kac4��ϺQ�������0�.$���&{v�6�L�OP��Ā3��:D5B���o�$4���YQ����焲��Ѥ����<�τ��!�b�+Ro@lw�SB��vd6�&�s�p� ��)�-��W1D`��u�U��3tH���.�r<��v��X�;f%���Ym�q��Sc��W{�y/�,��I���M���V[m�Νa��������ci8�I'��!��5����k411�ƍ�|� 8"��N?c^S��5İ�ý��,�{`kHEj�>vp�}X0��u���4��`lg�E�1|�|����RsP �����H�LG�����������R��(�V[m�j��s�p��K$"&z^�Ӥ�h���B��ﾛ����D������U+x��_O�2z��İu�����4�x��>�0��EA�ib�t��+��s�!~�*�q}n�Ć�2;��J_�qm�V;�,.�����k��G����j������tB�F��4$��Z��!N�B�[����Ԧ
4��r��p��1�k&���D�Ez��^�c��­�yF�ݦ�����-�3�5%&�)�W�����bMN��&E����H@������u
�wqd��K+��D�5c��������d!�>�1��n�v{�䥃cMRQc�m�rEm���tH�n���ڥ1�<z��\UI#h�D�h���mL�:4��!e(J�&����N%��K�����K��5EA#����)X>j9c����v˖,���F�f�ر�;︛�v��]���I4>Wջ����T�}�h��!vKr�]lL�1%�\��Ti��|��F����΃;�(}SmU�ZD���j���#�i�)���B��tC<$򍱪��Uy���>2���.��du'��H*Qt�A�E��%�Y��+Fx�9g��eP��ldL��}@TY��|ќ�[��W���w�Uc�p��1��,h����-p�9��ڵ؞VU�@3!ELS�E��f#��HīO�IO�tN�s��i��qY��J�q0�� &��o�� +�]Q�G���V�сM���@׳��
D*/�O��5��zR��x,8�h��xS��L����q�ƅ�<���x�g��}4�n&�����W��n%�O&X�"��~7n��o��F
5��:�=�{^�N�y�y��@��4F�"}��=�ё��|gT��)ɇդ�
�Y5Ɵx�y����A���3A�<�U�^��;)e�	��P�lڠ�hp���x�K_��w��|��lG�WM$��?����T<b�5�y��j;J�ׇ�rहH8� �t���n��r�KC�S��t�������)����n�dQW��Q5ݘ1
��C��m�i�lh�g?�|N\9ʈ�A|��*>t�ÀD��CT�,K�!���H'�`�N}��|���qk��������Z-��aD�b�AD��YK���1�����F���٤����F#1�ud���k�b���Q��l���	B4e,�(�HM�>��i$�x"������/���+%i��'Fr���opD#=/��;p���/Z��f�y�ӱr�;vg�^�9Ͷ�oe����=��s��Sى�5��a<�H�L~�t����b�Eq&B��Ynfޘw�R"�����1;��y�8�ښn^8�9@��o�Ńj�����Mz���>���0Ⓘ缷��M������$��J6���f�$��l����+��g<��	M'��D�$"�%;@�KB,A"y�$D%Ĉ3АH�<v~�i�������ei��qP�l6��6]SJ2k�2b	��"�1<<D�#���R�o#`L$z��k3�X�1D)
O4�۴�A!�d�`)4bLNģ�����z�{��A?����T NV��@��V�7� ��<̌а�|��uL��0f���h͙L�2�D?Aڧ�@�C�PO���v0��d��yGFH�*K��'>�<f״��!F���>���~�=�� ��A�C�N��������!�eO,kgIq�����F��YZL�M���-Q ���m�8��]ǉ+�qa/�B$n�n+�ю_�f�Lɬ�{�N�5d֢VV-CxN\�q�����nA�h��؎J�"(�@�>e�!�2�,ɴ�Y����a�4ɜ!h岴��PbF�`��3!Cj-6[� �<O`C�\��	�؃����6�C��f��UU�T���c������8#��սR��q�w��¡d}�C�c�5c��M��o��nbU���8oVe��or۠�s����3{2�ֻ��j{0,
�.ŋ#�g4L�V�k3>�xk-_��h������U]ˉ�k�!��y������C���N[��G�y"y����e��ī�aGx�Ͻ�O<�:FY�R<쾟�}����^�6BHt��iƂ�NZ�O���ƻwh���m��P9�8�g�_{?�,F*���m�����o������6��Ió��T^��/��㸡t����}��7>���PР-�H�8�����̖�n�󵌵�E+(ZBf�����|�X��~���֏�!��
DZ"�;�����*II�����Λô��*�>��P�-/�Q�h����ע�Lq֕sJ���}@6�BYl�c�%�<4�bw��z<�V��e1��.�bhƀ�L��H�J.�RF�Y�JQ{�j;�@Tbr�����M1���N���g#Mx��hֆP$QQA�y�O=�'\�S���\ќ��l�:~��M7]�׿��50�Db`�D'��G�Νw�q�q}n���)��-�����8c)4H.��:���_�<sډ����g���u�����u��H�oW�իGyӟ���=�?��7�@����e��E���q�e�OD��b�L�c�x3�3��?�~x�uĘaM����>�'�ΐ�*�`�YF�(�.;<���9^�dX��h�I�t�9_*���Si�*6ˉU��|ܧc�m�B���A���M}�4�b�˒�e�Pփ�����6|Fx`������[V�����&�f�2�<�d��e�h4ط��L�&g��=���B��t��Ot7�T��yo-���m@���fkk!��X��iY��\�1�RR	�;�8n�%���-�BP���<�i�����A��� n�\�d�}��p����|���h�J�P��!�~�rn�s��RK�ᵆF�vl�\����[��2[��������,o�kx̣��i�ϥ?���(b�;���|�c|�_`�XA����~�׽�ټ��O����kv��DB����ɢǚ�h�|�S�ƪ��G�����a�b\V��z��`�T@Jˀ���%C����p.���lj�+�vQ`�KS �A�bLp��
�<��t�e7G�����U¡���B�����Z��hm�6K��e��{�ct����al�4M�fni�bt�b��ݻw�]�vaCA�i�ۿ�}c���-�f�XM ���5���0 Ѡ`E	
J�ƤM#!�^\����"Mms�i�2���ɳ&e$�ˏ[���\@Í��4��@(K��fl�p׭��]�nF5�2C��!W���Vsӝ?9�CQĠ�ү�<� Ӏڜv����q�y4���Gs��'a�؄���~r�~����%�R`�����~��$�qZΙ�Nẝ�A"�bh�аF�3|����e���g��ߗӖQ��Q�xx�ejK1�
F#V!�JްdN!�`��a��
�*Q!%�H�9ʎ�{py�2g>NO��X������U��!�I��q:�ګ���mƾ��R�z��V��Ӫ��P�H�X<V=�-Ln<Vڈ7)!�U��O�kD
ψb<�I��j�4Tm��D�& ��I��n�v;=�]����0κ�V�q�*�xi�n{~�տ�1�7�''�	���M+3 9���W�wo�?������ԇ�'�Z:�(!F���m���P�u���8����v�)�6�}/K�:Z����{|�!�%�-A*�C��J��TwĊ�����\�a����O�c�k�����Z���:`������e/�)rR�����w�U��y�ǡ�~�f^���s֩��rV�M���&w��~��=�j�3���G����~٨P�����|��O�:N����䔢J�65tf�aɬ�I@4�EF�rkE���:�����n#!J%)�WPc�֏���
������������y}�j�vJ�R՛�y�CD��))�6��E Ċ���E��Y��I���Z�{����ƢjX��5ä2N�!T���G�K�.Ǘ�Sf�	42G09'<�����P$
")�J*��~�);G���6/�!���~�a3Λ����G���W^ͥߺ�0��2(b,N�X!��=�����#ܽ�~~x�Fbh`�K:��)�o����I��_��1�탟g\��7(�$鬎jy��<��AUM <���%,��+��J:�<A^��l�z�T�=:G��~����))����x�(��B"$��GX��u�o0�ݘPܜ�nm��v�`T:�:�Z�h�՜}�idS�j��N���И�{4&7��e,�nh���Q�2WF����C���6�`惞�qg�L����2�C1�Ӟ\���|& 9{HS�ͻ�x��'�����u����žΨ���BZvY�V�v�u������"8c9���Sv0���3��b�,c�ڵ�y��Āƀ�4c�p����i��[?#�vx��^=�B����Ѩ:�=�|�|���YNY5�Ѡ@Q�t�Ȭ��X��?v)��+	2
$���i3�����g���|��W�o�~�4Ȳ!
�o���="LB�J��"��������TҚ���|��E�U�A��!F!��q�vǝ�Z-��ȂA5("�+��	�/��bq�&B�>G1&��W���EC�	�>�����'֠fj��[���8`2�9*d������8>��XU7���ь�+��tq�����t�@t�.�c�ru��1���Z�d�%��-[F���{����u��0M��0��}$z�)�T�N#!�q���n<g�Z��q�M7��o�
����P��YJ�z��!O=s�/�|�#�D��c#����g��y*��'�ԣy�O]���s9�f)�z�K��J]\�0��I�!��f�_��\y�-x�)�pf�l���I�;'����R�����x(�H��B�����(#����0(h=ɥD�I����{Vz�}Y�2�˞�l.��7`��2":S[m���2ܦ'�6 �`�hrŋƞTb�<G1�uԖ�4��!��t��6Q:�B�_̤�̤4��a��&JH�ΒJ8�v�@�v�bS®Hrk#��麻M������f�4p��Z�%Q2�oW����/�X��@7D�&�xcLUr�b�O�a�"1�s4�%Ź����s��F�(�:�l����?�������m>y�F��T�Yf�y˛���<c���Wyӛ�D��o�����8�_���lo,���+�����_xዸᮽ�,f���&Uhu�Ƀ7�U�$0�
!B�C��Z�s���c��=AP4�c����v��Te~�ɠV����l��΃Q�'�4��
��� 8H��_M��9���j{P���2G�~:��qx\����1���pxq�
���8�����N���t��K��/i��bC�
������U�����Aؔ���Wv�g��X�P��}�gw�ޏ�M�sh6G�2�}[��;��%�T�{�F�Z��RUv��]-t�F�1��Y'/�"J.`b�9����j�}�����>�i�q���'bգ
��H�){����gl�C��^���`�]D4�MNި
�~x�Ox��?�?�����WB�x����ɫ�b&�����k6��Od2UsV;�Nܔ�^N�����'2�WCP!%��2��s�kQ����S��P��bU�L��S_�lC�d�`���?�{I�y�4����W���2y����� ���Ŧ��V޲/f��b�^oӌ	Ӡe��cN[��3攒S�1Q%ݎ��o�L帻R����#i*=�P�ŭ�?�@����R������*�`�W���W@{syP�q�΀5��j�׆�*#. x���ԥ����A���4�:"��`��F:���W@���BR'c4p�m��xD��}��g3��@�Q���b�1���4B)��2
c�V	��qbpyzX����-�y���?��|����OF!e
�c�"PZhQ����O<�����g��?�~^������& �Eiq���>�;�A�1�2?6tr��Lf��6�|FEĠ(�rk�r���r���+�4[:SE�Q��%��v[�SVJ:�]{ʰM�ԓZ���V�Q1�v�C}
�iG���%-I��#u�h<c�=c-����?w�g_	������q0O�!b�֏U��l�=��8�!y��u��ٲg]6m?�v�������]�P.�-/��hQ���3����@������4
{���1�E�S�v�غ}KV	�BT��/斍����N s�(��v��ծ,1�;w��*Q���gd k~.�x�������z�c��;������B#�˯|>��ڟJn�mE)�%��g>��^��,����{��⺛(d(e&N�e�B�e	�u�J] �
LG�����͇���x�9����^�Ú���h֤�;�G� BӬ3�ױo��aJ4��L .M�K��U!���/m1�M�3� ��Fe�MlI!�{F�,���� ���XN��K�����
���:7��ڎ���������0�JJ@t���|1�ޜk�,|Μ7���$GMο�+H,�2��!����#+�|�43�Y����������!3�>��6/�ľ" �- �v�Y��ֽ)@4�ݶ�kV`�EQ(.K�����'�����-�� &>��KjXL�����&-ip�=[h����䘬��]�	����.�`O{���
#��}�k��^J�Cl�I���"k�5y�{��^z����-|��w����I����9�(��i�ʯ�����g�˙g�Ο��?�o�+�,�[Vz0&�Ǣ��R_г0i"��ʐs,�i82��ݘ�0��{��O�l�l6����'�ߍˀ��������6�m�;�t�#B��_;	U�UKa0Y��S���	��o�%�k�P����㪰:�����+���=�')�N2�J����x(C��8�z�����d'�Uȓ��hW�C�d)_t�)N3��>'g�GhyN�P�"�4���c���r�`&E��UM���4 �� ��A�8��ynX�q#�Ԡ���\�Ƿ�_~�w� c�*�G��P�)S��	��/��ܖؐ\�FrƢc�4��-׬>*A{�o��� ʖ������v�?^��~Z��v�|���ӟ�4�l	-�Xh{Ъ ��m|��7�B˷�#�xl���Dib��BK~�����ox���ͷ��{>r)�Zj{0؂�IurVy_���sc�?�u���3v�N��%�y>�'��l���\��K@�1�s��9f���F�_�_��}:�69������0Iv��<�Q�V�Nf�>`*3�n�CQݰ�Nrd?�1�'�H��EA����w�hcL���ʲ��lR�e/͘)�)��4&1@�?������L�׉��k-���q'���N�����<�ې$ ��m��M6k-!���7鳓���N��P ���c���Ƞ�{�U�xL�1��b�X��D�
�@R~��$�p5X|z��:qā�k.+5�����X���Z1�*؎B�v�ĩ���ν��&��	6b"!���e��0z�kx'�F��*雏��y7�.x�չ!��d+�+��6o�qg='HKrch����߿�����X���� `��н0�߹����ɍ�i��W�"�����cB���r�V�������g�P_�[A��%Mb���&�>�������r��xbHڦ֤�-U%��İ���\�ė2�c�Fq.��UO�b�]�q�S_�P�7��ۜC��V�<�Y�A<@6�3��'�,I'6�6�dRPi�-�ت*�E� 5��L[�ej߆����z�t5Nc�R���+�#��u��L��9�s��!t�[Q8�eg�n�1F�*��M}!b��gYFaZf�4���2�E�=�d�����s���9߲,�������|�sn���7�� ��팩�F�v��=��@r!�2����l"��ؕ^B��q�goJ2��%���1�@UÅ���&U�Z��̜d@����	���5ڷ\L��⤱ġ�_���Fri!q�Ɉ��>������+%�����՛9餵?�ab;I9�ق�W>���bl�G�w>�|�#Y�b5�vo�[n���@�K��,UR�rr�wMv�������!�NR�1Pm���ˆ)|I�=A�9�K��lO��ȝ�C�f�iBĊPĈ�sZ��A�X��j�>E��c�C���mr��&�TV�LɜPj;�j�3�\�_���b1F֯_Ϻu� Q�T9.���ܳg�v�⾭�0�Ƙ 5����]p�<���夓Nbtt�����o�>��6n����_? ���v ���#�V���<��v�V�bɒ%�ٳg?��O������εc�_�bb�A���^x!�>+W�d����پ};W_}5W]u;v�[��w��=�\�=�\�?�x�/_���0{���{�c�-���+ٹs��x!�7�H����O��SO��jq�e�k#�N��(��H��'��ŮH�t�r�.���+G�U��
OQ��O������ p>aEq��@p�}$l'1U;e=��J��}P$��#��6 ��JRա�-:B�k�?� [����#_��u����3b�/AK����#����q�WPV�p1F���&���mi�2���w�`�-���AՑ�]�5� Kb�T%6ۅg�9���$(U����h٦�C�bE�`�a��&� jRs�X�X��ȢEC���f��v�QiS�BĈO��5:��X�u��>;���٬(
��&�zֳxի^5�v۶m�ꫯ�K_�?���f3ϧeg������կf�ʕ�2����Y��c����o��/~�M�6M{�'?�ɼ���� �� �Y�z ��v���7�0ಞ�>w�������g���,Z���C7f�c���Ѩ|�3��]�z���ﶟ.|�{�ڵky�_�K^�FGG��������j����>�{�����h�]t�gF��k��[�	 *"H'�&V�c�h�ƺ�i�e:%1;U�&V܏����ܹOH=Y�1S�6u.p9I�~��w$�t����U�S�c��!V�D+�y
:ú@P���j�J�M�+\>�D���vC
����tw��r��q����x��dE��~F3K�7h�-�1Q�����ECN�rE�k`�0�}�׾w+w�%�O1-�ݛ!�?B�LuN�C6�$�1Θ$ .��.<b5����w��XxU�!�t��d�	�f8�h��jpZ�e�@����Ҳr	�(�A�dfr�fCba�/���y�w�Ǔc2'���֥��իW��g?�g?��lڴ�����|�;ߙ�9e�U��7��M��O�� 3�?�u�%˒$ފ+x��^ʖ{��y�f�<�2�'�t�\r	6l����0�� oݺu������~7���g<_U��|&�����p��N_L��(/����=�7��l߾} �v��9ǫ_�j^�����˲Lq�> &�N�X���E/⢋.��~���뮻��T-�t��}��������/�@�[k��? �T�t5hb>}굫yl�5U�Qc�0B��X ]�qb�Q!�M�7RE��<�	ՐȖ��M�y� .�n��wN�ݰ(�G|	.o��B9Ƽ/t 
Aq)4��̪#fF�v!T��Q�(�IF3J*C�����<D���@�I�⚟��'�H�Jʨ���1�e7��f��qx<�5�%�-!��7\�24<D).SL���a��W��]��;����K����B��8N�!�*	�ss5��R��I��PvGB�nd �x��M��J�Â���fD��MK��ݻ��,�יe���]��Zׯ_�[��>��������ub�F�����E]��"�޽{ټy3��s�v��˗�v�ZN:�$�����~��կħ�o~�9��Ӻ�/"�}��\y��{ｌ��1::ʺu��⋻L�1����������_��w���׾����5� �|�{����og�Νw�q�s�9��O�TL�p��'�����u��t��Z���~�7s �(
���*n��fv�؁��u���G��9�Ӎ�<�x����/��/�n�gL\��+W���o~3���~�<wP��Q��da��(,�&#6#k��hX��a,ylш�<�X0j"%�2���,�@;��5x#��hs�+k!x�Í&h��׿�G�|N7T������n��/���ĩ%�S��Z����ڿ��ϰf��p�9��|�X����f*��'3�C��rI��ݜl#'���:Zn�>��>�C�z�8s�r�<cH
4��R�"�v�mF�|�n�y��l��B�ޤ:�	� �=�ӟ����h�X�B&ӣ�������]�n��k v�k���s�ɸ#�2Զ�>{(������\s�5x��̲e�8묳�袋xֳ����0�J�e��/�"�<�\r	@7�g2�=��y�_<��~��?��?�aZ�V�y���<�y�S��3��L6o����8�v�,˺��o}�[y�;߉Da��ͼ����+���j��y�	UUV�\�����'>�{�y�k�ַ��Md��C�����?N�"�,���'y���������#^x!oy�[EU9�sx�3��W��)1�W]u_��Wx�s�K��|�3��}�c׮]}g�!�2.��"���7a��:�ڵky�^���^Ja�����w�y���of�ʕ�y|ǎ�^����$u*!6$��X���ǈD��F�cC3(MF�Tqq�\'�d��-v�]�,cWlc���p��F�0786����N�S��)%�q��'Q�p6 �L��az	��c��( �"�#t}Ǉ�Ng��i�S/���?dQ�O��e�cf�.�G��{
��sW/��s���q�j�8\���� ��gM��㞭���M7p׎q����)�K�w�V�3Ϳ����d�U�v������l��ܨ�C�e�L�v�3M�"��H3��գ�y�1v���Y��;wr�e��������}��o���|f�}{�ӟ΍7����t3�'�������w���|���.�e�&&&���?ϗ��eD����n��&����B����@f}'��c;w��o|#�x�;8�SPUN8�.��~��N�믿������w�wy���UW]5 {��@�����������k�O����׾�M�� ≉	������~��?���o���ڮ�T��eY��o���ۿ�O��O� ���>�^zi7�lr򖵖�����w~�w�
U���8��sy��wL�ˎn/����*�K�1�˛4����;N�����S�MOH j�*MzQ�
6D�W�+��]� "6A��ФIH�(�'�����{��ǹ�N���n
$0��3�dwg��r�s~�)���Y�8S��R��l�R|R�g�rz�Wгb	�ޥ�`;8��gXaM�j�ך7�)A��.��ǞG��"Lj�r0�7�O�~�ưN8��G{"���V�ecZ��g-<��c,݅��\�7��:��5������6A�;Y�xI6�C�
�#pD>i:�u�.ϋ�\��yĮ�Q'����P/���T���\kC����3S���8�g�p�X6?�cx$M��6�X۶���M&�7���mol�ycۘض�o���_S��t�9繟��nr>i�y:�&�B��z�m�2h@�}j���F\����	p��<j�q�����䉎M�B��;�3�^��A@�S&���kc��U�5�0�&n[g'�~Ax�{����gJ��#J��
�C��N.|�$��S1#��ǎޣc������`���-�r��sfD�Y<O�>A�|�RLj��m�11��Z���W\�\p��kƮ���G��sF��m�/������!|׻V�C<N�)�1�t<�ۯ;Y?��}���'4�;���\iZƓQ�";Lwz=;L�ݎ�ܬ��߾L��`�i�'E���B
���la��-a����-��:^;���T��AӼ���~޴�&�Q�(l�̦���dL�[K���OT�50F1/�'L�X�;��O�}��Py�ĩ0B�R��u&Q�$&�v�`����3�>����s���Vn}1�����C�sض��ّ���� ~[����,�Ⱥ�b�V84�^���Pa���f��RlY��Y�����6;��B�qF�6�R°"2w~���8Mm���2	�R�k�u�����v��>*�C$V�.�N��� �DD�׫+~�2��ð�W�j����G��~�����u:D�_��eA���@�b~��D6LrHE�������㛅͵���^�4O����]?���BM�$M&U��&��y�ݴ���1C8��|�����1�"�ޓ������=���ꗩ��G �;l�Hd~�*��G,��<�| �1[�Lh&�C�<�hU���Z�m�n|aސ+�m�#����aÙS��4,#^���o�D�?��Ǌ�g�]t�L�	!C�����C|6�&i1WHD��'Q���
�|�� �R�`Y�i��@7�7c\��Jk�of������_7.����)�I��~}}�/�N�l��= '�������f���v[�+	��QG�.P�x�PN.��h�Ǉö^jׄ�<�~b^{xDl��9�����4�4�x~Wz�c(G�E|؃��$*R20^9�T�(�dil9�h���CRI%�_n1���t��x��0k�MM�Scjܦ�x6��.@K�Xb9����1,����F:��đJ�@���e�������mi��8֬�Z��LU_�ZO�MMM��Ȩq4�qꏋ20�z����B)�z[��8�(��;Z�gE3l���.Y�_�	#�
I�.�1z�34S]�K��>�`�~h>p���=�#q���
��@�߉.}�r{p�s���|uq��.��q��Pi���	�C�B�2�K �Ѽ���n�6@�>gǵf�]dF��+m^�7wfJb]���B8����f.gU���vo�\�C��L���AȎ�o�{e�n�tad1E����p�k��W���#��j{9)�0��X��X�hۊjl��׈ ��4Y��[Sۣ,'�+1��LRt������!�7���&\���8M�0x���:Wl��X9�mm����ԥ�h���r\4��u%�	�<:�������l�K�p�T᡻-��\�kk�UGdSz��� N5^o��2{�F��-�Q{�5�a�N���-��	G�!���H(*;M&K��ݦ/]]�xw��N�?�� �Wzg�C㖻B.�VA��w{{*FX��YE�:1��]ʥI�,Y_���f�(��jj��˾�#"�˛UP�!���_�M�g{?hxxz�{�	s
�� =	|�l>'���|Ue����[݂�����n"�D9�K}�=��G��-���:Vi;6տص����qF��c�:ɻ��scc��a0G��������W���qg�e '?ߦ��a8N�X
#��`��(�5L,Oog�a�W��'�Ǻn2�}��vQ=�:���s����o<����������aШ�����J�}��p��_�uB8j�� ��/U�#�[YXP1�[�`�.D���Q5��:�����y�#�qIw����K��h�9O��0uA4�l�\V�r���`4�X������.dw�#�F] �$W �M��/���Uy��~��3������>�vKґ�f&���r-��Y��b��PN[5.�e�6���t���b��lF˾)3�Ts����dE]�親bK�|-<�Ew93�J�m;�&����@N�B�w��@q�����߾���k��QY���~���y��Q�\Mn$��y��-�=Ym�����1z����Z��5�7��3[.
��Qq��\�_�濲��y��ID���:f �a=<<�@���e�{� ѩ��a9��q=A���u��{tyuW[�ua�j���|��r�%�I���k���'�V�>�Uv�ek<C�����у!I�(m��1=��ZՊ-[�O-B����h���5�CD�&�?��5j�f�s _;�+����k�[�M�څ۽j|�{X:f/-�x,!�G0������Eb*a����l&�L�Ȏ�k�T�	�ɦO�[E��%�r�y��i�o�����ْNqP���W	$"��	K� �1���{�V�8�t�a`�&�7Tq��A��������a�&P�$IbH��$_ZU��g�C/}�s�W���(Z�ͺ���}�@���oZ�+�� Ǳ��$�@�Fd����Aҥ;�)҅>�EQ=t�;�|�]�J����!;m�U�Mk6��ͮIy7���ۅj�$��`ɛ��i��.s��+�Vң�B�0��OC�[![�=[��eRA}_y2���IN��d�(;y7ŚW���bjJ#����5���V��,�G��Rʚ��ut��ň[f#X��h����h��g��7M�W�Co�z�M���>��o݅���񣋌+0����,���
{ވ�M:��	�39��$1�Ԙ#P�&e�pw��SQ�*�l���:��/V�i?����a���%C����~7�|��9�b��S�~���@k�VD���Í�w�nkk�����x���u���ӵl*�_ "O�W!�I��ڧ��g_��D��8�,�A��ك_s�G�V��������
1'gg�_'��;�+FC�+�m�aݴ�}�Mx��K�U�A�OU�ʒ��7V����V�C�ڔ���g���4�Rm�m]Q�U�;��7)��/�Ģd������~5X[k����@Dj2��sWh�}�HY�y�̓��Ғ:�s�_~G��Gj2y~��8�N��c�C�_Ԅ4vl�b����L~���@D�\�˰�0����ژu�����\�_N����aœ��^�*���b��U+�*$���#�!��.j�:��mMA:%*=rw<��zV����i��cL���b[���z��p�u�@�!��sYeQ�Qw��y#4ݘ���1��������P��_� J�����?���VZk����(��K���m<� ������a��д�q�9|$��_�dkP23�YUW�\��q[���XS�����U�k(��!ߖ��o�5@�֥=�s���A�L�0E��#�����@K�n�0��icjLs�� $y; 7E����o��s��A�����m<����rN[��3�����~�h��q �U��^��8��{3Ds�JD�~g����B���r [!�L��^�ޞ�Ъ�����eC|+����$5��_�,��aŪe;X���F�������u�����ώ/�+�e���	�ErG���p���X�q��-n�L5x%�¤��$� ہV4�8��͕�տ�<��k�+��]^��Y�T�ʯ�7+��r&�s�=���rͷ�:�	i]g�8C�Bil�/w�,s�S�1|��豉K/뾟�_���Q��N���܄�X1���+�.D�Ҷ��PgA���X�ЯA	<h������1,_�3���3S�6'j�Sb�7$>����o[0r��ä1g�g�� l�.��F2YY�����wm���7���G"���5��h����m_��ϊ�$*ꨙ���إI�tM�xʿ�+��7f������R�]���B+
����=^B���X2=�r�˲/�����%�m���3h,@�"�^$I�
�&M��%�� ���l������L�v�sl����<���&�
s����T��Oɖy�L�Kb���E'��\b���F�%Q���#��b�� F��?����x'��י�٩�I �H}�+j����q� ��Q��2�^�'�ی�h;��Þ��]��������Ֆ���m���/m]Z����x��N�a"6A�|��"�������>@�V�BqY2����d����E:b�B�Q� �"��A��L�B ��헪������'}w�j�B*�����D�Nl	���@����!���S�#���#퀄%AD#Ĺ�9t��UJy-cD����Ιʤ�������X�G	L�.��_G��y�D�%>f�,jA/oH�V')&��	�E!uA��8|�#�����7���"�����<�]7U�=<�&�3�h�E�� |�@���,���~a��mς���u�����*�_��ߞ3�-�|Ch�g8�R�kET�$�ˏ�ü�W5k��AᰅP�<Cr2��ь�O�Q���������%ѝ�4F��ah�
<�@>P�<v_��M���#�t�E�Ȭ�`r�P���}bq�@q᭳P�G�>����[��9�d������z��4���Y�pAd�Iܸq
��?mo�N���3�S�s�k\w�9K0Z��L���n����4�o�����De�%Q8o}��'�Ժfx��$e�hY������~a��,9{���c7�=-��n��rT��L��(�1w��6�$��W���8�T�MZP�Nִ(R��w��ʂ���'�B��-�ya���_�A�r����?��Os+Ѝxh�� ��t�7�g����&���DN�JTP0G��쭕���mݪX2d���L�C.7��3��=�*�Ĭ\��ZFS߹���*jE.e	�/1���C2�E/d����`�,�r��|#�w4�o`@�3�x@z�bh����}�i�|��n$Ϋ!.�^����pG0%@�j�OT�u�]��tG0�*��=�53�B*�;;;#s���2gˤT̘�V�������l7����HW�z����W���v �+��H�%R�?}��(N`�"��x�_ u7̈́�0,�.����R�4f�W^��E���<���dV\˻�����!s}�9��
��[29�e�Ec߻�9E�-�*!=)%�|�����,.��x�3��*�j��
��l�����i�v�H���.XH�?*:�W��e�	8��cg��mD����t���f�B�K��!qCv��dE�\����EЕH���$J�i���6y�LC�I��Bi^7�i�[+���
3F|pe|���RX�פ��p�5�/6Vg.�4&T\��!^�))�#y<:oL�����evZ"�3�'�?-֠��nɘ�u��|�8i�%���t�-�C��Ȋ%���ZGGG����lE�a�ҿ����C����x�d�b����G�KP���e`�
���� d�$�::9�1�q�m�e�i�� ��6XO.+��Dx?���:ʖ�K�?P�6�o��_�����H��u��Nס7�j WT��C�����t�+ e�P��W��̓�G�+/p���8M<�^"���s
2����Oeq��6A�5��9Q츖�4H�z�j�~��WA�4������3Ìh��%1y�*�=��;��tZE?�#��A�(X�2ٟ��l8ٸoQx�@��'�O�=�r��vZk���dJu���q�m�����K��I�F�8��!a��v=����A�Q�gǑ+�+�!�y��Qh��w"A���,��z���G8-�"�?F]�	�K�E�eˬ=���P<�}˅qv�}c��8{��d�J<_<�DNɢQ��t���n��=5�|���J-��$@�h<,q*�2�(���|�������|	���U$�fC���X��4ސש֦!��<��׏ݟ�`�-�?�ػlO�K���-�}A����t�PL+"`7����靟�L��w�@��x|ϴ����<�Uύ(8R���A%?���(l����>�;ڄs�y����aUp[YP��Dp�8(����p�)�u�A2��@Fv��Q�m��*d3G��n�b�i�B�ԕ�0�E��˔+c����R%��0:���/��n���hd9LQ&H�ExsEV������n>��k�瑾K�F6Yc�v��9��������}	7{��s4�͇Jm�Е
����A�u��	.*����៥�ĉ��f}2ĎpEa.E�CvuCz@�N�l��=��M�u�2���)%(�Hɪ�����C6����yÜ���+�0lӆ�֗w�;�lv���?�r��Za�e+T�a/%��z>�Ziݽ�������&��x��F�������*�ڮ�_�=AyJ>��U�kW�d��Q޴-uV���'��Z/?gS���=/42���җ-�Jg'�n�8��Q��o��Qj���dw��y/��>n�.Zv�w��{�`��[�6,�k��$�@��:���l�BP����� ���׾��*.?���8��m<��o�ɽQK۝G�WJJ������^\��0��]�c�.&�������S��C��hl$�	5�Dq��)����ۏǫu�8L��ƹ����^��?ZVC-#s���P���"5�IbX�v��VN�yo�*$����k�ƿ�%xJ�%���8����]�L�S�uT+N��%�J�JR�	4ݐ
�~���Ej�����>Z^�q�����Qǫ���6���p�����aWuٳ)���F������$�P#��>;f�fF�$%�z[�IE��e�)�_���k#�]m�S�y�~i><��q�_���
+���Rt{��! ��DE��FJib�嬚s��y1-��e<�*/�lL����_�o�������jH���t[�*] rc��L�d �׷7��	�{��4%�������.<�ng�C�얘����(C�F��!�.�����F������f^U� H�SE��=�x��Aާ㖪2�����#��`�j��~���j_�!AG�}���sdb<
�8��*[��yS	���N2wAw�V�Y:���PB���J&�^}�z+�yE�j��\'W����	�����:���➒��Oں�+��s\�#��&�J�j��'���C�90��{��8�E��-8�Ӕ�廉��3�yNK�$���8�"�A�����mg�>��*�֨1ل�� d� ����\��*�F�ґ�:/(�&�*�q�͚�I���K�.�9=�/Y��-J�Hэ6Vte �`���^�@x�T����c���q �?������K-E�uo���/�`wE�bnIp7E���3�����x�89%.d!v֊ê�ɿo�t�H)I���=�1�q� ��c9e6T��Z�(ǎ`ï=���.d�
#��:�7��x����h���@�F풤�6P<u��2۬�L�L�B����]����Vw�R�����#�;�LV6����`�*�yv�*�����%��`�Ҳ�n�w3���(���"wHe�h"Q.]�L�ȟ�y���F#ș� g�x�X���x�,�rǎ�U1p��<5�
�8`�%�������w�cl�]����8������v����xF�|�K�-�s���w���ۿ�7�ts�}̞��牫�rd��sl�#y�ԉnV�|�&,��n�+�F��2b!����w����H-����fG|9��B�DᑻU+�b�{����dq9b&	}�Я�B6׮�p0r�\����"�VSdq�[d6�����O�|@�ݝS���͕��׋�ͪ��t�Ѕ�,���E(Eú��~;���SV���_��UԀĹ��g���ϛ��(,�WtṐGjd��f���h���*�	\��*�v3�n�0��J�ѽP�PA��$��>���y�8��s���Yg^�=5dgG_v���Z�x㔬��(ti�(|0���:���,B��d-�Lf�^�����ŵ�+�I�#����|�A3���qF�~87��f��
AN!0R1{2 ���vy6�2s'���j��3��������a�1|�_{���؉��%����0�~>��
��L5���6m�j�K�p`���v�ئL�%��g�}?9m~��w��f��}��I�|~�����|m�K/e����_�j�N�jp�~ ��#��?%�r�i�A�C�r,�|�6�]4�$D�* ��Rp����N��~�\�'p���y��f藀���b}�����B
��vs��Җ!��Q��()cB�m@3��ᅅ�(F�H|2E��>�^��
)ZW�$��M�a�FM U �>��K}�'#�)��	4������48U#�[!��S����1�:F[�Rf$O ,����J��O�~\��x +��Y�<��P]��nj;��f2�74e���S�'�bs!��H������?��ip%�O��.��{ ��Al�t�"WI"�5j�я��5�@\�ka@8��!J�,���[��
����;�4�p<�&URѰy����D�;:��iJ]qQ�md2Di�4�EA�n���Q�U�B�'{Bu��R9�&$�ݿ��^..�?��ʄv�0��E8uzb_bQ���R��_P��s�X���V6Q��ɡ�d�N�8o?T��!���B��ٔx}�޸�ܕ���>h¯mn����_��5�@DU�@���Q`�۹䧔�����]�,�i�3�S�\��؉by����ȬpR�<Z���C̌P��_/O!��1XgV�Zq~~�u�F�w4���okky'��p��L�!B���l�2~����h�\�S��&�0���M�K8�"�w#��0�������P�_S�����}QƷ��>on4���NQ�fs��S06h�v���$\��� G��=g�F�	|��P�{���A�P@����IT�V�VdC�v"ю��OO#dK���aqB
��md����A��Qk!bn�z�����S̚��E��Ϛ���a�׺�m6��`�xJL|>a8m�t����8j#�g#]�֫����=���6Ӱ����Lcԏ�Ǥ�z7�8s{�z�M��#�A�Wy�}˳��%:&�&���M�\o$�򇉉���_{��O)�Ah\��K3�V7L��]��rr�i� "�%���X׫�7ӻS��ܪ��pC遮]
тfM@+t{Ly�����B�dl�x�(5��&TKD^cAy�3�e+tɿ�����#��oh�2��G��-�IX������&+7��e�ED���[�.�Y-�+��+஠Ą$�Է���)����=�K�p	�3?�w��^އ5K5�u�����⎎#xQ-�Ӭ���mVtp�i�Kvh��
���(ͮ]��NbeD��]B��#Xtq��߱����5@�׍���)�*�=͘`��W��ji2��� :�.�b��u�nT��m�F����Ӌ�z�_8P�H&|Ұ��b�u�S���!_Kx����6s�����'�`�j����<o���OQZ��h����O����R���+�۝��� _~��}���#��|���s-�,�-��2~���b�zIf�n��8s}�́�xP�Y0I�B��=����}�)�q����q�x�~��v�3!/�0�^M5�e�n�Ӑ�Qݙ.:xW� Қb����<�6Z5-%+�Y�c�~����8�0n,O.�����c�ᰎ@I�$��/�<�!�*)�4X��k���͓V��m8�C���0�yXBp`�ǋ��6��E�\�|�n���s���YAJ���~��˃�P�f��&�K}(54k�j��z#>��fM�!�bz�^"���:Ċ7z8W}b��7�8Bys��9����2_B-��?�M��r9lS���kәP(�6@Z�9v��(�?w�/{�8����6�ҥl�O�E�S�/�:3��Q�B��jf�����8���خw��x�0^�l��Rp|�ϼɲ�墸���$��ǄE�l��Ui���|���8g�vA`���Ӭ+*�ϝ����(Yo�K{�8�F�	\!�lT�#�gOܑ#��X���ꇐ���^`&sIf����1,� ���9����ղP�̀�'[�P�7��W�t����HxC�b_Y&"O0��[O�Hfk�� 鱔�`��w��0j��9����/����3H1�̴�ݾꅚ�����G����m� �?(okį�Fv�]=h����r����< ��^C���O�L[�מ�Ű��Jswk�M�xZшQ����iq���n�����+�G�P����n��d�Ȼ�5�B ���(&6�~�R{}Qe.�C�m���IK�'������{���84LG��3d���@�"[���ăW=ڿ}�h�����-�lm���+tb��x0��J�s�ɺ��S�+ Q�|bw�&�C�u��q;�<����|���j����yw|��:����?k�|�T����j�1��ٰE��An����=���jM���ca�H���c�ҊŞ�Ӫ#%8��~삗����&�^wQ5P3�hTHS�G�:O���{uSї�&����!�'���Ф�-(z~}���RЍ�.$�X���!5})-�}�^��r9)���:�d����P��Sau��I��s�>�<�G&}ѯ�����v���zʘIâYeD�����E��>�������[�>��$7��n{ǣ�2�^E�&{�e��~���G*'�S���˜ԉpY\�o�v�l���R���LEaӐ�q,Ǖ�?s{Mf��p�'X�p>��xF5�?`8�LS|ݩQ���_�>|4�jyciC�8A����U��[ůѨ1��u.�B��$���b��O�Hѣ$`���k��wT��\��Q7R������.@H�ƻ]�Ɠ�Mo�N$�m8������#U�R����s�[��O7���E]�O���v���7��o�S�n��3"�͖�	���0s"��\\Q�[v*�c�������I4��9�BIĻ�f�.������*��沝�7���1Yc�LU���9���]}6k��Q
\aʿ�����ߏj��E�߂|<D��p_��Y68\�^�:|{px��(�k9NnW�d�2O�Z	N���q�)�]��������<������$��I�0�B������f��&�����Q��U2/��ce��т=6��5$�,�^R�;�@�]Tti��VG��g�Ϛ֊�����޼��#Q#�mH��S��$����uG�E�!7KM9�d2��A��D?��U)�����wj�#�Ԟr�Օ��ıD��F�{�l�T"0b�����Q��� TϢ4J�4x(��ߕ0�lD�¤�����-����6xؓ�E��1�ڎQ���$&ee�b�ۤ$��cpGp®
��x	pQ*(�Ts��RQ�G�.�Ka��p��%j|����?����,�s���3=|���C!(Eײn��{�t�� }zI�?H���m�6�]��d�]{�g���2�$A�'ڨ|\�,	r�Z@$? �ZT��V�����Rάwn��6�r��SŌ/���1�6�~��~��p�	���[y!E*�^XB�B�v��!(���~ӹI�к��c���ĝ��k$��#��e�����ҝ%�RA��#���Z[�n)�� ���yp����e��W�0���I)�Ik�]1exQB�R�L��+ǈ�kw���O�@ȇͬ�O'�Y��q��x�Ts�(ܡ�Bj��	J���>����˶9�\�jX��ֿ<�-S�(=����W�sM�[s�/e���]/m����ŵ}T�G�����<۝����J�s%��ݹ��&��|����Zm��^�@��k��Y�q����J�'Ҝ����E�`�B��X�H�t�I*Q'A�$��];���[D�AF�FH�y\��mNa�[�@�iYoV=☻B�-�l	eh��OqH���}�>FP������`�fhq�~h?I���'r�� u�|�R<����H�RJ1߆�E/D���~�(_�z��`�<hz����S��eQ(&�+��t۔�z���9��/1���|�^3;����ϣ?���p:��_���2��>z�'��}t�%�m�,�}���3�9��B��bȋ�
�d�X�G�/s��zT'��Lm$M������-e�CB�O��  ��:�<rO��(f�j�u��)-&�ʯ��z�`,@W��whi(�����"����ё�Jb��D9��cr�J,~�D���bY����v��F�c�хvd�����vc�]Ε�0R	EiԲ΍u��|Y�t������5��4JB�D�ɽ2Ϗ>
%N��ef�<��e�|�?�v��'��
�������@ti� �/�B����I7�H-�\��oDw�V1��C
=%�����#G1�:2 ����ibֆ�����=V��k�ܲ�R��AiT5�9���I"���hs.0ij9<	�a���4��s��c=ǔ*Oj2Rddң��[��l��2�h���;;+���^2�����U�\�T5­ZF�n�BcEʹ�+����/�X�y"����2l�ި����ز	Q�\d����~�����iG���^�\�ߨ�����Ҫ�߭TԺ�ahG2��K�y�A�V�D&��&e��C]�5����71�B�ʍ�gH�}�[�A���3`鲝��U2e'���:�4e���P��8.iE��h���.�}�;�N8a�3��#1-mMV��Va�],-���6��迋[Z�怭n⳶_�^��8��������-��Ñ��]��h�!-G-��'[��$
4�:V^����b=$5��K������]�Mͼ���>t}�8��H�̼e���l?FV�U��4�S�8����Ff����XR]�w@�(X �Z��jY-v�*ǹ	QmH���T�H��.�#��ת|�_w�k�t�������L�h����T�W���t���c,Krk��_�-��G&��$3|�|`eW)�}�#1�}���6/]6�y7�J�؉^>�� ��\D���y���~��`���0O��ښ �]�_3����E��=���<[�\�Ϯ^�?��W��,Gc(EIU��냓"S��>�T �`���[��e7]����Ǎ^�Zq���՜���l�j�pA�9��R�$4�cwy7u�5���%U(0/�}��J�����Hw�� `,�6�O��Um��#TDJ��kb���p��t�%C���������ţ��3A�0`��O~-��:XS��l���1�׺�q$������<ɶ�S���p=�v~�(f�|�e���ỉ^���7�i����ݡ7R�����;g� _��V�i� ��.gx	����0�%�������Õ�'q� ��cȯ����W�Q(�f��{���a��\�?k:+��?��4�3�:#?�LMn��،������(q��_�U�w����j�}og�c�[ry'Y��\
���7P
�AL����xkMC�<�����S�j
!����/�B�Q�n$Y�>V�(�F90'��k�3Dϩ��)o �+0C�Ҷ?1,^j���R�y�	�##��.��Ǒ5h�δq�,%�[KE��wB��ɭ��R�L��6&���z�ICE�m�j���K�nݱ�,Җ�t�c���)��"�.���X��U�̽_�a�hC�\�l�F1�*�����KN��B1J��&x4nY���{�o�n;�Dz/!,�O�]aխ������ќ�h�x���'���p
���B���ѝ��]�Ҫ��vR�����x�fT� sa{���,�T�-��ڇd'�յ�(��P��0!/�
�?��{�+0�����1����)DY H��L��N�m�SaP������a�H��D����Т�� y����>Bn;�z\!\7y����T����񟞏)��]���~h��­���"*��"94f�)8�dC*�}C���h�������pr�lwj��<
�����0Q^y�2a��:���������Ϫ0v�D5*������%-�<�H�������P�fs����Y���К��0|��(MI�G��Y����=�Y�Em�ςm�,2���.S�܇D``3�i�4�jO���-$.��7�,�n�D���7[���2K6^+ŃB�v}�c8��zL��!�b5e*��Eի�b2�/}�=����=Ir>� ���o�	5�W�!t�C՘��יv�Q5R&�6����vC�=H<�!r�^�q��n�J�`w�Ez�CT����t�/�#/B[�[FeV�n���W2�w�j�<�c^`;�"�fT\�<���*.9i��݉ �tg�7?�J�՛:���ڊ�� �[o�%��~�V����f{Ӝ�8bsS��v�=��o��Ǐ�b [�p���C�?Y뱮o�ރn}�MI�Â�B���,��ym�m�n����(�A���)��m��^��?��V�Z��4A�٨�߂Fa���L'�&�rL�]�o�V�jiXs��e��;��.7x����r_�KYDe�K�V��ˮ��Y"Gx�r��T*��ׂ�#U C%
fٛ�e��0/p՜���A��;tU�2E�"�'�"��r��@��nP^:�1�R��
��;fu �+q�"����C�BY����z��t���}���!�'�n����A�M
d�B��T��s��8�|�ђ =.����FG�|a���e��҃I2���5�J����fɵ��@b���{�&*S� Pc��U�Q]���TY���Ԅ啈�M�2c2���Q�8`v����挋~yy�,P]�KC�="���sa�ɖ�J~#!�6��Gͱ��KçABJTz�+��&��T�� ��kѱw$#�*О�����G� �ËB�E3��mZ,���H�7c�� Sݦ�=�6�=��Mb�Y	hl�g���ve?�x�
��J�����T��4;k$�������I��Y��&z����>�s���?p���"���z�N����f��[6�%0�vd	��q��
O9�,0�`�_	Mq�h���_�����1b�����<��'wm,K|t)�X7�Lhmb̄j��h�`X���>���N���;:��ԥ:�'ɹ{%;��r��D'�_�
:$�(�n�-������|�
����ї�����(#�"���u�P^�Xf��L�{>e�m���i0�?���w���ײ�y�:�������2�6]a���S�a��9r:�8�;�Y3��YYl*f��n����Dܪ}���u9��z�J��{'����Y�)�����!���w����$9)[e�r�0.� .%�4#F�zX3�,����X�_b�t�|����s������[��
y�I�&ӎV���I&z�2�MTz�7N�a�m��L�l� �������\a��kT8pʢ��2[d��S� R�_�V~��<���y�ieQ���Ii�;(�����>"��)TB��-�)�2)��#�;37O�DC>~��X̸hC�ȯ���EG�j%ik��������rDW�p�&B%� ��%�g��.Ԧ��9����j6�k��L��w#�� �L^`n�`Q����J�>ߟf�B�G"��AJ&�`�Oꍱk��_�>9�T���bX�o�X��*,s�ٶ�X����'�ʅ���͗/��?�;^03:�{B��sǺZ���g�
D�/��YA]ͫ`3�nA!�b(�O���_�z~���W�e�Q�/�%�I�wr޾̵B#I���=a�BA%4"��"�@�۴�)�Ć,�<��t�ϰ���hPۄ%�@�.���(P6U��1A���i��Rye��ߏM��}�U�Z��;&�x��B��bǨ��e�O��s�h�O����}��� *bf���� ���d��BI�+�O�ѐ�r+�#����{i�K��I#��I3z�Z.�Xb~aͪ�y�V<�~^�A�փA���8��Oy-�~J����� �!�te.6�J���D��b��V�m1}�����ZlR}v���!B<��H������Q�k=�^��W�X�"�y1�T� ��-=�y3��o�����!cs}��������ş;\5ޮ���qS�9	��c�ڎ�Q����e�M�y�ˡ�s�&�ޖ�4KT�)�2
n� �����}���5�~�M5�xꁉ�>v�En�m5��oZC%�9��a؃�<�`']6��~���_�c���؝����t݌R*�e��
��e�%�[B��\2''7j�y�_s����{N6BV���%&����|,F��M��ʹ���s�,��D��<�����ӿ���R�P�?n�'5m��1V-���n�H�&H	�l�ƿ�I�.YŠ�8^o~�j�z#�����O�M	r�c��3A��nZ�� t@�����	�N�P�rN���9��3�h��h��$��v:?��79��8[�O}���|�KS�l�����8�Lk�'g|��.��x�Ɓ�b"!y�{��;����w���c}��E�r֌ZR#��l[2^��w*!PJbC�!�ɽ�<��ʤL͠�£0.BE�Z���R��5��]�$I�8.�UC(I�u8Q
���R��yL
��(�8�U����Pi��$��C�'�>���I]+.k�x������	�s))*$s���|8~��)����u_�l���
~r&[N�F�K`-8������{�7�t�����\ �s<�C�È0�%+j�G��S�d�Yɺa�v�Ģ)ǚ���>������e�<�ĳ�F�`��洯���.����%��x�އ������#��'��������o�bao��+��>|�kc��;��Kf�K�4'��u�uǽ,^
{�=#uʵ��	\��T*#�a�|�#o�G������_�M�%l_�և���>�骇F[�s�`"1��(��-Ze�e��d��ai���I��%i���Y'��xUl �;��m4U��iۇ{և�jǿ짳�	�u �2.���[[�{�Ԋ����厜������ws��vc�Wl��t~~���Z𝯟N�����s����|WX�V���������/3��/�k~Ќ��m�C��ӢH��[9�����i'sڧ>�w�D�����x,5����"]DxYf��η�{��n5��~��|�s���8���p*���_&n�:~w����C���˙�v���m��9���#�e����W�������?�$����M7#3�d��Ba�YQ�8d���ɷ>�y?�.��ǥT���c��!*ݍVERM���y��|��/s���O�C��>{��~�C���Y���!�b��������.��R�e>��mK���{������񱏞�y?���B�(c\��[/��>? d�1�!2�+�P$D1ڲ)�����^mZ�x�9��./Q�d8�.2N�΅r@��x�BX�Af������>�-΅f�P���w&+�h̊�&�X�+o~Ʃ�h���8��c,�H��k�U���:o���Z<�U�y.W�
��Lj\��Дh��u}2��*<3{>��0�+FR�@��ߟ�Q��O�r~Ƽ���d s�;�Y.��lƌ*�lAJ51��̒������
�dݒ�\x��R��bv�~2��s�@M�7myBe֬y���9�Q�J�,�j_��L��g�U'���'9�S��
��yt
/Κŧ��eV�R�띳@��0����v�{	�>�=.
[-a��X���<���g_ !�]�6�\�q� RY�������f-�:iq��râ8�9E�f))���I�ڊ\�9��)[�����ߏ�
E��q�
G{4+�-����_�wĺ̓�<�o��g>�����a���~ƍ̸�6"�&�Rـ{｟��w�ݹ����Q���@6�AY+jIH��Z ��_�q%�1+dPב|��YIR�y^�?��~���� Y�ʫ���oŹ?���}'R��������qءs�_/�ʈw�~ϛ�W��9"Q������W��3�~�����?㉥� t}�P�4�t�����T��Z.�� G��23n���f�O¨9�%"]�Y�*�8������G?�1��q)�r�=\yՍ�����E���W��	��m\v�߰N����o➛���%ˡTBh��{7>v��������+b���Ѹ�%5ߴ����ܳx�ϫ7o�}�R�:��,�uD�h^_�S���x���YlvC�T�o�F8|��4�)�Y>J�;�p�0���̒������E#d�{@���?7n܃�l���%z�'�1N-���& �m������н�!"Ez������\t�l�o}���Ug�b_��x����Ky��G;J!�
�M�ޡKR]���cy�5�cJX�|�#���c����ԍF�Q
 ��9����".���D�W%�p���l��G��7�'�s4;M߸�|�����������T��b ���KK��7���m���O?��R�;��aL/&Q�t�CL?b[��1~~������jL��i���~5\=�曵��3�ht�}w��/B����f�]���[����G�sλ�vj�.�ى�8|/Q*c��#�5���.��1(��^�n�-7^��ݔ�
�a�<���O���_ ��#+.����=#�� ���Z���U�Ț��'������N[�]/HK�V���}��g�a
����R�M�Q�r$IJ-uH��%�,�7�=%q���11%�d�A�k{�77_�;�vW�^��\�3?ѾL�6�'�"DBsnegpR3qÍ���Kn�Qv�.DY*��r'����xH�2#F�aʸ7�t�DL%�Ԭ��`��������9O3�R�k�NjR��L�
c5^i��'�u���WN��|�^�R݉S�g�� lѠ~�h޸�$ǻf������"�/}�C�֌Z�g�e}'�C�2�m��E�!4�5�"�����+`����(������M��Y��1^q7�r��u�ޤ٪Z&֘���4���͕��9��;���*���D��#	(3������@F����6uC��(F8�&tgIi�*k�,x���M�/1mڴ@u���9�Y�b#GU�2t}:k(��,�IIm����سsѕ1�5�Z��w�(*ћ~��?��_��V)).�S�Z�V�G���Hx��H�b��o���3��o}�+��}y��'����vt���C�`���y\��316e���D��H��7��Y�X�0��(�Ƌ;��6�����Qq�P�#����Z5`��CxQ(\��܆��fz)QZ�LB�2RgQ"u�m�	���]o9�w���� ��I�E�RCo"�����v>���÷󶷿�7��,���tD�0x�sQ($BzLR��?�=_�+�pecT\j�GdCGf������)4R�(t�{'��-$�d���N�Z���o<^H6��):�w��(�y�[@�$���@��Eݕ��֣F���qo�MI��Raв��%!550%5Q�q�YV�8�i���uH��B`d��*����8&uilأH��X�����_��Vc��OQ���֤6E����_۳}����ȸ6� �>�rf�/� �0����Y��V�|S���V��F���m
��k����8��#�5�.�� @�#����sZ��$q� ��9N`51�d���@��Ȁ�\yDT��E�	�|r���`�"�#������[wg\E"�B�4�O�RF��ט7��z�F(Fu i7�*&��@�Ǳx��ko#���P���ջP�/B��D�J"p�	���A���w��TD�!��K��"|�B��˱6��Q��%������	<x�T{jx!Ѯ�i𾆌$K��� ���]K��)Rzz}��"<�]H���)���Y7#��!Ne%h�2�`�hŤoH}��]/���VD�ZM�[Rt!��.�E���L�M���5ߔb�u�-D��.�K)-Nu)�"���~���\{ŵ�y�/H�@���%zzR��5b�;��xɯ8�̟gZkD�I�H��A)�����*A�l##"�?y�5�QRg>�a�ø��PT�Bg)ǒ(�@�*Z��2Ӽ�X:;�H-:|�f��ಿ�����t�
.�
E(���V�16*�<b�lL:�*���*Ӄ�IA�Y�&Aw��Rh�TX���g�%L��9QtL���R����M<�=)^B��MHSI$�RY]O@���g���w��o}������|�r�q�J%�{{Z��>���S4��em�*N�~�Wa)O�hYn�9wY�֕D�}~������:A��T�W^�Wd<]s�;WwoY���<�Og�B��Q�����AB����٩�����yL�]�o>�k6;�H�L�I�h��T��1nX�90�E$T��5�3�[S��ӝY��Ǒ�D��)Jt�����"Aa0�#�jr/.S\v�=,31��E��52��&}�C�(�,qx	ݔBm���'�q�Z"����ƳK`��ᆛ��{n�?w\�~��e4�D1S��8Hg9Q�"���И�shۚF�k�F4���-�mh��Qr-�/rMي�Ǹ\�������3�?�C�*R$̙����^CbJj�L�;l>�b҆S)wT�5�9��a�BQ�1Ԫ��;Aoo��c6P�e�?���:X���j���8���@R�l���gR�I��k-�K�YRg0&�k3������s��ŖԜGG[���DQ�j�j���gR/z��^þBo�0�IE)��"�1�Ѐ&Jx�L�3s^7�n�c𛦆P��Uyほ3��y��2w�b����V�VtV"�⥀�������]�U�����n���wt]e"ۋ��PV��0f��k�ĦY�hpl9�.�����h�Z^�����뚎�,���W�ݠ��5�#DȽ苇|ón��ጟ�z���J7IbM�R��
���y;�<��^Q!U%�n�ܮ�p��L%��;R��(�U�����T�fEO�˪쐃�V��H*t����r��'r�=�0�Pk� BT�0W�v�-��Wo$t�-6�'�Rn �{����u��B,���o�\���?��h<2u�j7]���/��&u��������x�Nb��	H��J\u�e�3�H)�u��.2;�+��6�f�G�z����:����R��z1I5��H�Q�ȁ��+�5E�5��eB
���j��淿��v�̟����ԉ�!��ϋ�̆c*hG��p�l=��s��e�n���w�(*ӡ�_>��P�dX�0�V`��G���ͷ݅�~�� {�%�?�.޺�\ѹԖ�byR姿��mv|�x�piVK�>`/N;�3T�Rbz�*��E,�YƱ�=���s晧Sf92�$�z�����볁��M�^>�qX���� �esʾ������Cy��M�L���\J4��$�I�����XzL�]/�n���9cG�B���nT]¡�X�C���=w<�}O-�ţ�	C�Jq�ۗU~��!06��8�={.�}�3�c��	"M�� �qYqM+���mm[�˻)f,�[�C���O���׿����t�-���^v��>�Q%>�/��?��^y5��q�0?�٩$�$�1�+J8b��R�ċ�4V+�ru9�{���͹���x����}�c?�A�^�yɢ�:ө��$	�e�*����Ay��e��T"x��p�o����M��·�R��o�t����?Y]�s.P"�����|�}�>���7���Na�'|�S�C�����;pQ)Cc�w�����.:�{���o���,_��q�{�]�G�(q�_.�Y���w���|�3�j$
�7?�ᰌ�4��)�W�'�z�/����;��7�=>���,�R�=�۶~�ϳf+A�\��c[3iM���9�����l�h�@��>qYop"d�!�V�U����� :Ie����摙��ɤQL�l#&O���JQ�e� T/�aO?��<��;pjD�q�K�� |�ΗlI���
D\C=����X�k]Ї����BIc� ̯��u�l�:�G�0�4G�^��f�3��75p��a�(��H	ހ_�I%'�xbQ���C��B��%��#P�e��P7�ƷIhc�Ըƿ8dϫ)�T��E�����Xt�̓����+~��tJ�w��>�_����P��}+4-8�ң�R�}��=�H'��c�K��G>@�2PHz!5>u�GiL߆�L��e,
�l +�!+�@�����[�k�3���cMI��v�u��?�8RU�ۄ.Qc�3�8����R�[�U��#C�.�W��gR��#r	NT��7����EI�_�=3�d��.)��".��m}7l4n=�(�R'��Tئ�}(MT�ɾ@��a<�n�\c�c��O�^Ţ�B�t�@4����N$8�e�t$6���=<���(o=f$JJP
%5+zzY�S�fR"݉�A�g+ 3�B7֠7�% �+�9gdN>�h�[M^��ֶu+��Zv�� �9(P�����(�e��<��C���|�����@�e5����[F�(��\~�H��tph� �ZsKИ��eu�9UXho�����u�2�N+���yװG��Z�lsm�{��s�R�4P
�L=�y�����f�%�� 039\/�,����)\V��о�4��M���0���'���M��KR��\��,�m}�Kg�Ic;���?ܬ���ʃ��� ��&�� ���{��,Z0)������6����x�T@@��l��r�F��h�z�Nz����%ms�nF�i\����Q�%���mkۺe��0��e栳����:0��^g:�Iqx����'�cm��Y��$ox��g߼ھ�t�f�/���\����1���	�� ���5rU���Ӳȭh`�Ȼ���Y�Y�'�,�l�.�6^�P��3�꛺��1��rnE	Y�~~L#��.��K��`�m�i2w#��	��4E?�[] ����}~o��%I��l10��Ce�����\���=Q\��k�JI�7P"	!�J�8��-!��e��)�����:��@�����*�l��ub���/8�ʣy�CC4���r����7;'Zǝo��/'�[_�{��^��|]��J����o�,u/s Տ��@5�Ck���������̷Ƀ��"2,� ��1(3	H���>1���O�̧���YM���X�;]��wٗ
��kѸ.h��i����b�dj���"���'+�"��xQ�l��S�i��V�f
70����(E��I{�)l�i, ��ʖ�Q����,��׉�㕹c1�<��:*t��G e�\�4�_���ep�>�Z6��m������8j����5tE?���~E!�Š��3�����[Q�x=�x�h�|I��p�i)^dܘkT&J��Z��d/�|���/��*,yT2�^?�<�� ʦ}c�q 4Ʀf'9��F�}���l�<5��>�����ڥ��8�}k%�n�{���fq�Fy܌�0oȐN�1
��^���m��Xǰ��Wo��2��{R���RT(W}.+�3����J���1Z���S��c�F�eT&��,�-��n%;����Vv�W��ȭ��8m����^���7v+f��I�? ;�1$[��BMw���x\;S7Ŀ�U\����^�k]��t�ccw���>�~�K�5 �ֶu	uX[FJj��r��y�uM��f *���s^
�?�:s� ��ۏ�mm{	qK���͜��E�`��VȢv�1��&�6m[��ֶW�:#���mU�j�v�۲��(��-m ڶ���Ԧ��
�9��9��B�����~mk[���J��I��T��)�����G4rD����h[̤ۚ6�#q6��ixUSJ9B�z��.���+��6�)^q���3������/H��"��Զgh��ֶ��RM4)V�6j�;���i� ���0iר�c;"ڶ��E���$�uI��b:(]�܆Q�ZbPZc �t�#	T6���@���,u�X�.Wp΁�I�挼��{I�-^�%u�ֶ���h½�M�m[ͯ�φ�¡��c�X�&�R�o ���M�޶��^G�6БYYôsxdS���#K}v��DK�s^�ť�T���J�:�@��yQy�鶵�mm2rim�l��ub/3�h�o!�_�u�-�cJ�����x|��N ]�uU����@��}�ֶ���඘�9wa�f:$�]y#b���d��R������ݯ#B4 ���WJ�5�Kj��U�߰@T�`Y�0�ZE?�Tmk[�֤'ɚC���'D^�[���pk�� P��%��k(oVr��%K�Clr��MPV�� a��1��ň��DZc�b��.^������fY>��xJ�C�wGD[�p��KO��5�ok&@%��_��D�'ڠ�mk�Z]����Fi�w�R`����i �:��[|�;j^����6�2�ĕ\��f8��/�韛5��B���l3��Oi;"Ӷ�ۄ��`�f3r�"�*7eX T��_+�7��I���6 �x/�B`M��|L�^�PH˚h�w�
��e{�t嗳�;o�[n��4(�	q���XSHe�#O��G�a��nR"��H�@!���P����fg�W~9n�/��rHi�"�G��<}ޕ/�r-���m̀��X,tļ[���ŗ�Efz����<�� Ǔ��h�n���ܥdgݢ�!p� X�
 �mm{��֊��"uD���w�4n��r��E���ƁM�.fs
h�B`�J%��퇸��с�&�u/�ߧTb��u3���w�ײ���)�*�,"V%|&U\��Y��V�ô1L�l2�͜��w��e�	��Ij�%��~�\N�_��5�qj�{W̜�r� ���g��]!���m[�[�X�A��e����3V
�
��F.�&��aFE�m�vl�	}��T���͕l\�O��6��m�T��E%�r�9�t �w������^#mlM���E��$%-^]�σI~�S 5'�K���{Dm9S�)�ggƎP(���1�3Fjz3h��Z:���6)3m��\s�yzN75	*�����:2��2�/�q��T���l H���b�o��ֶ���Ő������E�[��zlߢ��:�L�JM���@@��Y�C`����#�_����ֶ��dV~���Vk8,JJ��`-J˦��o�X�����{�t'�̝� kRʁ�ڶ.���%1(�����M����F,jشZ/ߒQ��c���GህG��(���ĵ�~���[R�Zi�c� Q�]�άވ���-%�9,!�{���Ρ %I��kNڶFw�N�-���J��xa��6�w����]����E�KI���=A�B��8Cmև�p�<:�8k���u�5��
��7/;}W���phoޡ�����~ϼ@�ֶ!�g�깿�=�Y3c^�&}=�����5��h�/�52|�v�!�
��u�Ƣ�0��@�N���b޼�v�PUb.IQBae�u-^DԪ)�J��P�"t�7ք5�{�H0�x-=W���U�]X/A��f�5D�P�o<n�ЇC+�ԝAC9R��>I�:�8�P�/�x��h��(զ9m���:늱{��îO>�'�K��,]����X��h�7h'B�d�cϽ�W_�f����R�Dbjw��t���5-(�om�@�/V:߃ΰ�&,�R�7�η��hEl[�ڶ� P�f �
4�2��%�)|�q��?���N���x�klBy�Z���N��xg��2�Cpؾ;�!z�}�3)��$B����x�N����1,]��ￗ��soೖ
��VXcP*�,o<pw�t��,IS�T�hxm[�H/�ʂ�X�Y��1���e�Q#�JJR�Y�k��t3�,dq�
R5��1�y훫�*hװ���>�Sv!�����/�? ����a��>{Q���(l���kn}�+��YLڡ�Қ�������Q9t��N��`[f�/M^"s$������yj[ۆB���A�_o��7y���*nH��� ^b�z�W�9�C$X
��P+� X3FI�w	%Wcǭ6a�%t��<�9DTQM���	L�h
"18�2j�T�=xS�:��,Z8����|*�Śn��xaQ��q%�>�l͕w>��*O��UI��o�k��7ա� @}B��n�1[o�6�p$U:���x��RaP�hR1{A7w��9�����4�
�ҕ���x��(hVλ�Z�,Wr�>���铗n��m��RbTD� �r	� �m��S1���<P*�PJ�����+������ܠ�ch�5�ؚL�����i���mh�i%�� Q�4����dkc�+qEM9�W��W��\�����&)J�уl�	O�d��	��<'��H�v��WC�PQ� �BɇH��F����]��nq��'����ů1A ��Ȍ��#�N3nܦ��ɓ�ُO'�1�a=%)����n�M�����$�h�-z��Q��Š� W)��V��H�%2�
)���9p��2qL���sKP£��g�qz����l6*f��f�n��1����
S��
Q�q�g��]�R �:�!��k�>��� a��@yP.LB#]��k�g�� �c5}I�x�^�Y����_�u��8���v��X1XzF�9Y�;!c��;'K8kݰx&[�"*k��g����+o�l����O�Db�E�q<�Գ8�Y���l�3T�u�Jl�mm[wM�歞�g^�F�˲�s�� ��5�I�����?;NE9�6K����SOq��k��_����p��s#��::��;�x�����{��ٿb^��ۀ��U��ʣNHU�_�����h�R�<�h�.��1���WH(x�iv�)�e�v[N�S�+�3��� b��I��?�U �M�Yg҅���u,R�8餓9��o1v�(|��#�`]��m¼{�)��u�X�Y����ïZ��Hg�6�C'L�x4�n[F�)�-C��TH�$W,�
�w�PT�4	SF�x�!�s�ݏp��/ⴣfS�����M��(pY1��ك��E����]d��<m"��� ��q��\N>/���O>ãO<S L�q���"�vP �2@&q����XX�k\Yt�B������]�΂lPlr6�B?Pݶ���m�D$�Ҟ�rE�S?�{�؃�ْ� 7���c�g��m��T���.	M�"H3we<=^�h)�t�d�n2����-�����W��eF��"�B�}�ٍ���z���(����s�o��a�R83�R��J�ZCb��|�-(�����%����-Y�A��#@x�.�淾�뮹�R��)�'�B�xM����P#�v_�H�x�	���V�����T5	�B�q.�}CtI����[�H�s�n[P*�����AƉ����̭�ET4���Ժ)*$�;��Q�F��E�	PE��Rf�Z���F���¼nFCm�w�nO	��o��4X�]��"�.��
\�-B"�/���F���%W�e��`�o����f��p��пȚ�s���q��ֶ�&�Xl��w3R�:ǰ����?G�A��+�=��_~-�^��KL�x2�n=����]$6&% N������>|�;y|n�޸�5��<��~�8v�R�?{�,������[��J"�$�7�#e�?�=������>���_�z��*j��q��(E���F��bRk���$+��l�ͶXc�}�9Mi����k��o�ԩ�!�Ə��,Ij�Cp�UlVr�w�"]J�N��A��#2Y��gl���q>萦��RY �8��H�đ�5ʱ@�Q���k7�Z�r��Ϣ+c1�����-�N߈�eWV�I�E��+}�N@6Ԁ6$'��5|�m�N�PBfT>K�{�r�l���_y���-�F�0��Fi�sC;�V�049��1 ��-ْ�,A��Ԛ@W���m[��ֶuܲz��z]x~��o���\J��Q]$>����x|�,n���ش���gʴWs�Q�������o�⫮�cx����8���3k>��x�d	eo�s{����W����Ȟ[nδ�ǳt�����$�C�%�ǎ�[C�����1��ҁN3�<7\&�"pO��O�B��� S:F�(�4���`���4D=�#b��׽E-�t�#U'K�%��oy�l0~D���x�b���ZfΜI�$�K!R����x���vߚ�s�����:W��C��$q���\	�� .;oRe1g�Q�95IB�\�Y�5>�D��P*EX<��6�AH�*�{QԎ���3�C	��P���S��c]���p�����>�6�6 `Ɲk��b%s��(R�؋�g�o��g��~Jw��2D��އ��-�z,mk[�ڶk�[n��2����9�@����D	�>0�8�wA�Ԓ"U��-���El��V���]9���կ�M�p����؅�Ftp���0{�
.��v����x��q��%�i���ʘOWG�R9��B*�����ɛ���~h��Ф�%�x6�d]:!�L�ħ��*������r-���2bn�����n����&	���84֗�ħ?�y�*#L
:�M�]�S���~���}� #��%�P�e��~K���!jޑ��fH�X9���H�"A����n��­w!�j�!IRjTT�&%<��Z��q�HM/^*R�|��tҋ#bRT{ƿ������m��S6!�
g!Y].8��� |�M��Vj��yq�f�rB��g#)�R���M�Og)�g�������W��>��:�
�w��Q��;SK��"u��mmk���p��rտ��G�ȁoy���ˮ�Gf!lh�����x�fi�5�
R ������"����;x�Ỳ��)�CW��UNK|���z{�ᚫ�q�m,����u�a�?_M٧�B`W�A3�� ������=�r�~+-��5B��n
��&�I�u����1Va��ŗ��3ib�7��b)^�84�-eʕ�|��2F�!�Y�ăPH-�|��O�_~���ҽlZV�J�G	��i����Gy~�!Ѫa�!�"��p����ᣏd�m&Q�n�ܹ�����y����o���1^J��xak	ox�A|�c�vZ'`����%<�����_p�Cϑ���h$W_r>���s�����ޔT�@4�]}�� �:��z����P���I&����k�9*8U����;����o']i3[6���8Ԛ�����ݯ~���Fؤ�aZ%�g�}.�\v%�Pvcک����Uk��v������䔳/��7G��|��� `��^�z�?\s���_�"U�ʈTz,XR6D�� W�W�ʘYs�P6���F���5TT��b�}������[���������l�~�.l6qO?�"t�Ʈ"��P�_����F�̕���ϲubP\���I�ʂ�.n�Y#���[��B��9E����6O�I���6[l�p=��;������|�#'�e�B�xG-M�Y�E�����k��GOo��dD-5AC����V��GW}G��z��_8��u�I��$TD��Iǰ�.��SN�G���g�V��?��|��Ή�0�3{�%�ƍe��v�_���%$N�<�iߋZǵg�h�q�w�;�&����M?���+O�m@⼉h5_��,�Q��^��8�*�F�L��5�U�=�P��\�ke.f(�>�+��S��y����4Ҷ���6�?\W^�elG٧�Z~��p�{?Ù���o���_Ą1��sw��S��c�ơ|���C�kP�l���N=o�RCȔ��QZ��ә�	��pBi�TJl�q�����>�(eP6�h!���5=�
��I�:�9GI�Q�����	�e�u�!�>���?���a�p�!���'%�Q�h��k�ډzl[��ۥ�p�U��S7�"kH�P��1��;�|E�-�����%�!�B߯(q�����?�O�<Nx$	�{��2��x'Cb3�"�4񈆌{���74�g�=��o����O炿^��:��2q��n�y�{��&5R+jY��K�~��^3�����������[#��&Md��^�q8�Tt����d���m���w��U��D�M����(� �mV2XlF����U�2��J��a�T�+����y��tk#P�A2�m�6#n�O�=�����s�QMm�*,�����tF��Jw��%�g��勂�}7�}���� \Vk�y����6S�f��B�D�d����L�R$��]�toݶ��RL���gQR"D���R�AӶk��Z�b��Mm`����us~͖=UʥcR��|��~�$�S�45tv�d�ͷ��_�_��|���O�Ώ}��O3�p�"<J��XGTRl8a,%`��y,�����)�g?�^F�|��|�3��u�f߱Ϯ[�ᘘ��j�"� TX�\�� � @-I<�.���FG�q�	����Jl���L�І�M��E������݌am5DI��7�,^^��28���b-�9�%��ݐAE%�β�$K�P�Ef��O�\x�#�z|?����p��)Q)��Bz	]�.F�K��P�j��ww�:ѽw��}�AZH�����q��?�1��B�܀W"u�es����[��ڛ���X/AV�o�=x��!|���q���"O5�xj�r�z�V.��&� /�A� ��r}��&����%�l�͖l<q<¸A\�Z����A��	��Dp�}�#[ɖ�A�k&7�����X����	^/_h�^����7��.ƪq�H5Lv�X9����y�p�ߛ:� ��;ԅ����e�
�$I���O@e�ϝ�o�"��h��ֶU�އ�����t���L:ѻ�D�֎�R2w�"}�)���%D���ׅ5uoC�R�LJY��5 c�JMO>1�O��n���l��(F��d�
��)R�I�<����HGo6��C�`4����F��8Ŵ�7f��F�IP�3��������4���m���=UZ�L釢��|�^������Pޓ�x������E���l���3~�a�󅿣ҡH�R�E��s�I|	kAˁKW�� 4u��E@-D"A+w��ѭOd�\�j$�2e�����S#G�d�|S������^"��]�f�M�9���H>ѴfQ��8���"������������%7�J�G��2%�QV�J"uD��XX6t���r�7D��ݔ5�����öDB�zY��(�F�<����wߍ�!#� ��:\����RJ�Ը~��j������he�x1�Ғɤ/�1(�I���?�z6xB�l��l�@5�b��K��U�?��e�=�"�)�?;�p�d�e�#�o[��6Ȫ+$�Hq�޻2y����Jgޯ"�wCK>1�=1�Ǟz:�v� g�>�_
���XD���8"��M�T��^���)giPV�A�)V#}�:c��y'����16��naiR�7.s��18���s�/�*;�N�|L";��u;���އ��w=�߽�yCV��Gխ<���L�d�[���U�.��S���۾�"�X[�{��!S��ӏ��O��RH��Tmʳ���)��R�U�u���N�sD:»�<R�&S6��)���2ְ�F1wγ}�Z.��~9B� �8̾��'\}�����8��o����/�����E)S!�EE����W��lK\R��ŗ:Ie'��*�R%tF	$0iH�TH!���>%�}b�b��eQ�iAEzFH�tv��l��\����Q ����!5�ݰ鱌�M;ߏ�JZ�l_���^����=��rI�Qc�b�����&w} �B�Mh��h<����EL[�w����7�I/2�4**�7�]��^���Ubi���AyCI$r��q(N����R��:�T�f=*�����/~N�Y��?�)sUyz�llZE��.���w��y�R��� �ucE��'C�|�-%jT��������u����g?�ə��<W8h�pՄ��'#]�Z�������c<�x9[��:��9�Mp^c������nv �R�xn�r�.qL#�n��5���oT�a۝vY�b� ax�����ҿR� lBI���%��U�S���QHh�ĚSV�Ҏt�O<�{�VTk	Z��-S0�7(�H�"��w����>��aF\��)���;9�����y�8�(�:�(�l�Rf>�4�͸�?\t)�w�]�H�d��#��<�ؓ�Z�+d$I]�����T6pB�R~��j�Y!��pH�-�*֎���o��'H�%B:D"�U�ظK��c	;ƕAk�2O�8�\�R
���J:��()�:����	�*-��{k�C+�T��d�q�F	$��RV��Om�{%���@��\���\*�jf@T"
�*��K1o[�^��U�P�d�����(h�U�؅�3Wg���`�u.��b��*t�g|��v؂=�>�@**K�����fr�/~����<ܲ����?cι�ާ����*�V@Q�F@AT�6��F�hLr�޼y�_�{�{soroZ�.156J#�K#=�TPT{��ךs��s����TAU�<��T��{�f�1��;��r065^�z�R.��rJ%��k�����|���I# F@��bďsԱs��;n��u럀���/�� /����xë^̙'�ĵW_��Ō6=n`1QS�1��JŪLk��6�
�s�uw�׽�D� Qq����/�ʫ����ujCK�f(	v�ΰc��~�W�8���6�-KNJ�f�l9W]}3Mu����I�Z+l�:-�Vs���͒E��96l`!s�R��������F�n�vYkiƀ��W��U�����k_ɉ��q���p��'r�KN�=�?���Q�Z�3�l�
��~�Ո�l;�V�O7s���Ԡ��=�L�۵��gss�tS�{R���(�o�4j���|�i�֤1�~�C0��J�կx9k�/&�J4�$F6�9ǝw����H0Ӯ3mݟ��S�S^|2�f�.�R��(�e�x�{?��z"���4�;uZ��C��J���؟�ٷ��v?��6�b���Y��J?��B�|�����x�=�%{́���pߺ��W���΅�v���Q�70�$)�v�R���7�ko�>�i�)���f���%/f�·���1�� ���{U���^�[^�b������n����EKh,@�'��PÆ�c�|�z^x�
�F�!�XXIZ�_��?2��X7��E�)�����`�&��R�A��%�r�Z��{7���mlj�j��n�	��:���hl�AYv0gbD�oz|._��
<��c]�s�v��َ3��	�kޤnje���Jf-F�G6>��O~�_/���9������/8|�0����w��Q+FX�~�}̡\��)\]L%u�I4�T����F��#'�-C(M��t�`�r��4�S���'V23��9c��z�F�N=�������Ţ���!�U�F7�}{^����uѣt6U%�@T�M/?�z}8=SR(�ؼ��e����0L���Cg_#{.Y` ���8���=&�Av
��>r����j�vi<Gum�@� t&�ef~^w���'����V��������\��������|%͘:�EA�m�⬷Pg�\�9F,bJB�d�#�Qf^�&��׾�y���_��1$_N)�`4��(Xg����y�oML\�zXB%��)S�ԇ���6	�c($��`x�2YQ��FZy�ԍoİx@���M���"J���]LƆ'����ةC ]]�:��0�_����F�Rd��Xk0��Z22���`H�O��TV�l�22����+�sD#�&jd�,pev�D�����H,�7�A,�6��!
7�w?�������-aQ-"Zr��]�K�9��\�M,��TZ���U��X�(3=�f/r�1�B��qD{��V��*�^�k&���u3�{ܭi������E�){^�g��ԵI�)�SP�Fz�1ja�Gۯ���q���%2J�1���E�\K�F��Nwz^Sn(�j
�gv���8'k�q�z^��f�|�#;��=�wQ*e�х>w�U���^�ѽ>b��>AA�����Z, ��O�9�_���C5�Iv�(%o�2@)uJ�S� �2Ęf�;l>LP�F����\�����5�|1e6�9�K�-�dd�`z!�l�3��W�$�����Z�J0�R��`�d��|`�s8kK�$9=/����]~�(a�B,igᬄ��B�z�XS2P�	��&Fy�i�A�}t�/��F��R3a-M^�m���9���=H�ТF�������pN����ʗ��)@-�ԁ�A��A�bzUR���/0<�W�5;��0��w=��SH�3(�#����.��ޅf��Ff3D
r["q� �P�J`h��F�_z���k���=�8�GeH|(�4�5�<C5��(u��(푢-QŤ���TC#�;M�8�J�M5F�ˑ���� ��_���1��{j.O�p�%����D&���U��ޗv�Bv;�Ą�WH����o�ÖG�3Uj�RU�*e,)c��)�wk��Djj"��ʉ��b�bĒYCn� CC�������Z�.)�ׄ`�6M�Z�]�����7U栛�NkϨ!F��O���誒k�e'�Q�e��!N�D[+��������h	���3r�Y fu,Ri�v��n�:�D��`lj009��=����t���d�R����u�W7m��G�>�^�?�:t��^P9�|Z��9&3����&�>)�h���1Y���FqYƶ���]�}�f>���TSq�*&���O���Bx�1��eR�02�f|u?'�A��zMxb@��z�Z���!�YC(�XI�ն�OH:�H��f��ǈ�`\�14�f��.��l��zi �f�	����˴���*�:�Ԏc%�9�4�U�b�Mm�퍜��m\w�v�,��+�s����6:j&C��FJ,�`���m|��;�V.&�㌩F�O|�:L��kc���bP;��l� K���jc(0\�����[�ǑVwo���j�E��8W_y	�A�8�@(=;Gx3�==N�l���T���<��O�O~��yډ<���CA^��$��£��������[y�c��曹����A>��O���?ȊEu;O=�q��E��e'���<�:�J�P��
_�BI���8Y9B-n�v��cd���RLfh��o�,���Z��}iĈi7����b�	��e��`^L��Q���Y{eW����Dz��i��ne�:@,���{�:�<�CR�h�c�d���E�-S�қ)2S���0.�M:N�b������ݕ��>�ֆ3Ӫ��y��AQ�uQ1����|~�5�S>[��߶���g���c�,�6 ��@rn~V��o�S�#�M̓AD*�%ƈs��Z�<��v���ǘ��fG��;'ة��g^�����l~>a��5
>��N�E\��u|�q�#;g	c:��K(�"ƵN#�(�QJ�&�4d1ޭ���;�����o�aS2H��+35��X���Uh6?�����p�ʌ�,�𩖁�ｉ�7v�7��\��h��
��%�\Ƚ��D�5Ѣ�6Pc<D\}�u�v���������L%4k����x�?�O0D�<m�BX��(���_���H4tT���?�+���������8��?�#��f6�\�_�@��`�+��ʟR�&��+o��_�Ƕ�3
M��osY�����4��XG���ؤ��/�%gH=�;�9f�?��ũ�'�`�T�X�U��ٲ�	�x�I|k��f$�<��H�N�.	(t63)%:ss����L���t��.�=�#��u@�l�wNGŪw�{b5{k�g[[�ۈ���a*�ǨMN������)�I��zi�P�3�7���D�,J,r �b�l�3�?T�f�I�e�	�3M�1k{��=;-s�����S�\z7�-_����V�l�0CuG�h��h�MOmc�����<�}��-K��t�����h[���!E����b��� ���L�cMd��;����_���s9��z6U�����G?bxQN͖�N���#D7D�\���n�=�e�fQb,�Ї~����n^���9��U�4��<��z�����o|�Q�)9�P4F���W?��;���Яr�a+Ȁ��-;ǹ����|�;�y�`����EZ ]�G(��l6SI����"�Hv��D��r�J/]LQ<���4�,[��Y|�w�4Nj���^f���Q�XZӵiv�\(˂��Y�Q�e��t��|�մ�m"�I�a[ t��;zg)�3]5�j�ɬu|�r�
H�v�������N!�d͜�y�SR9Njp���N�S\��?�GFڌ�V�V'��8��{�tS_�8����R�8|��n�4�M���4W���7�ޣ�l߾�իWs��S��ٱc�<��v�`�ҥԲM����s�b���ޓ��M�ѭ?~��`b�z.Բ����f� ��l1>�+�]X$�0T��jOO���-�o-��;9��#0)$T
2Ùr�����|��F#I{pР:�1�җ8g	R�Qs��p��[�n��UOW�$	eB��N=�3�������E��N����跋�qCI�Q͜�$��9�K��K.�jBSk*Q�h�v�h�h����I8���Қߚ�m�����F�����QbS#}C�٤V����ܹ�ŋ󎷿c���e��;��w��e˗�'�H�H?*����y.&� �&�y��Ⱥ��4us�e��-��q����D9;��yO�X5�aR�l41U
Sc5	��36MCIH�.ژ���zCX���J_b�� ��I�_��B ��l��<Xg�!bHSOd��0%<2��ν3R2&�BIcf��=���ST��Ϥ�P�
<�<d�E0b06�o�FS��Ma}�ph�?�c��z��b�ߪw��!Gd�T�����2��N���0�1��Ո����1���o�Ŋ΃��3�b-!�kB`���y�v�a�ہ?��^�"|��r�-�q��\�"ibW��bd�R��%ke���Ը]�U2L��f 9��k��m5�ĥ*oSժ�����-!R�7��S����(���G��F�h="�Ify�����_U��Z���aL-M_��G���{6"��x��ä�iP�	@i|%>y���I2�h'�����J��w�a�U���I�����.f��3��x�ok����C�;G8���o����m�Z^��8��c��k�|�2�u}��!����Df�ݔ���Q�4If���6v6#��A�Lc1����+J�4��z]�2+�/�1bm^}��8���P�A�ш5��TѪ.�eDA����9LquĴ���H��S�H�bF��q���|wSgWj}*/a1X�(�'Ɛj���c�,ǫ�.L \��RE�� FE}h��zMFYpu�2��g��@���$�h��>+
�* h��b5�ŋe: j&1�F�9e#�f��㛀���L^�S�t����f� �r�U�
�	E�1.����T�X��D�Urs�������ieYbL�O=��|�;S@= �xN>�$�8�����jժ�#R�߾=�����U"��&�mV�ie�b�3"s�?����QЪkA3K���f�e?[�x#�Bf� 1�	0�=�.۩����x�dx��;z���6J�(��2�I]0i��+mU5M����'��8�Tn�:����d�(�Ş�7�$�,1j���n�B���
�ǟt�e���3Ng���GQ�eA�� ��4��Y�;��N.���X��g�ǳ��IU��7$=s�$�|ǱU@$�a��5q��kw��dNY1����%��4�U�����[�1�ĩ2��XCP�4�`ղE�t1F=V���p5�n�ɭ���TN�j+]=ݍPj���C��Y�|P$�c�4���x�R�N��1�V�t� z�r��k*v"e�ʢ�:ǎ�&���[�4pM�$/}:6kGz������@�����G�&�0##R5�A�����)�z ����=�b�q���n�c)�0c���g�� N���g٢�/[T5�6��|�h,��h�������)�'`�Cb���G��-TJ2��r�C���Kd��$������L�AZ��Oa�EUٲeo{��Ȳl�la�%VE��l����7p�E3<<��2|Y�S��V�9�y�7�k����I�X��ı�s$6�ot����Qˬ5��Tw"�a�����۷��S�a�Z��Zt<�*�0�t�Y�oۛ���xw��1
7L�F���2Qu7\����?Ǌ��.G�j��!b2��b�d`�/����c�kY4���k֢T����m��8��Ӹ��{p�M�j�b�	��m �(DzG�N��ֹ������!��}$F��д"S�0bu�	���ǒp��!��EW\�]�?LQz��)��39Jj�+}A-��ߚCy��Ϩ���4��)5㺛�d����V��n��)=�X�d�W��<2-pF�@�4�7�`�?���fY�� �)�y�|
����P�6m�|
�����J�d:�abd��G�p��/���b�>�B/9���#HN�3��Х����CK��t=Z�\*�R�����~LK���M˶&?`�e�<��v���E1�c��Yz$�G?��[� ^���1:��s�Y�%/=�UK�dm��HP���_|�+����%5���zQ$ib�ɜj���ݮ����O?�z�>	xN��U�����K�r��36>N�>�O��T�g�ikXJ���3����(�E�a���&gsJ�^��UߤZ�mFC�[�m�ǯ����q�B.K���	�� �3"����p��Opӝ�s�$�(�� P�N�j�Gh�H��T�]���I����o_�^����@�0����;�B��������U�Ve��'>ko`�&�"�v�r��m���o�Z�ĳ�m�}���tӍ,]�;���3 �}�Ev?��P�Q���'N1+����.�x�u��I�<����"՚���%�uV�T����j�n뢂']Jgw$�S"�Ҍu�Ӫ����;z�����%j��82� <CS�qA� -�ؤ%8]�{���6�
�s[áE� �B�ּF�ҥ��h5�A3dX7�����Tڕ�&�W�N�r7U�+�J��6���%	�7���'�o*g�Xk�����ݡA���҈��1K�q& ���Z�[��#J�'����$oKF�I��A�4C�[����۵��
^M%qSC]5�B:�M˗������!�6m�ī_��D83C�nVҗ�u_��WY�jդ��۳�D�k��U��8@aW�7�r�Y����j�mU�qDd[��uw<�������p���q���*�����6m��C�6����l�i�;k���r��۬�����̶���</���@?��I��s�e˗��Cw���=�v�z�1��i7���.O@�W��%��lA��|Q�@F""YNz�v7�$ɡ�2iR���᫺��k��ĥ1}Z}^�ٵ?�#FofpZ��0횬�
��Ҥ 3Hw��H����ɷw����ZK���0LŶ�d�.}��Xu���q�ubV �����`�j�S3R�:�j��֓�|�Fq�{�{Kó7�*F�5}�;��	��fFtٲem߼��j�0������ٟ&b�ۿER�h@@ꌔ�adC�7<����5|Ԥ�D3H�C>��;���R�Ւ�] 5����ƍ�@�/ᴻ�}�z3
�����u-�gv-�ȼ�gъ��JV�.�{_��5���^�zFt�cE"�X��[�vߞԪ��@T�j^ڳ6��ҒF	=s�5�X�H�Ba��(���m/���خ7��-[���7V��kڷ�6���)$Z��tҴ����h�y��s���5'e}��N�~|ݠn�׷�S���n�� Җgb��^�cd����j5F����}{zi��B���T3d�Ғ^&u,Fc�V&��y�m�g�9�m���t㻬BY&��GFF�g9׿�}��Mo�Z�)R�bR:W�, ��������>B�_bM��zb�f����Yg��HV�;ژT���cm}FK'0VY��}-�ʅ^cL��wmC띷�J�GUbLd���n���;�JU��k*I(ӖIr65��d�1�m۶-��>F��Ǳ�,8�߷�=�@tzOc0�3�-����7���W/�9̫�޷�B�C#�1�~MR�f�De�Qh6��FE�^���Ei��kL/�;ӿ�� f:޲���x5�s��2MKqI��eU�S�r����b����*�#�Ӹ��]�T��l6;��t�o�:��,1b���'�2��(E��^�]/�)}5ha/ �"�#�<���a�֭�y�/��r}����8	X���ac���]ߊTmL��FMt�o��ۮE�Z-�,]��a�M�6�)��Y����'O[�[1P-�+�@�Cg��7��F�͈:��l�B�w�t�ڍ|��ms7 X���Z�eA��EQ�_�2�T�J��V��U��]���j�3�1�z^RM+2"���s�(ʂ#Y����Es��-��[R a���˚]Z��ʲd||<��9�,���eIY������bn:8`4E��	�+����GaN�����i
���H8-Y��+���W������_p��R��>ר���m]��ЄVQv�� LN�v�+ 6ud�	��+MK�Qg
������3����g����Z�7������Z�V缰���q�葝j�#����X{k`��Ǩ�FX)M�v၍�P�e�Vd|+CyFP�J�� ��λ��Z�/�J�R�O>�$���XzF�#F��+�I�o�8�zH�j�aD�I�H���������
��Ӵ�	 W����N@����O�7ȴ0�h�!|����f�/^�M7���'�<��_|��,^���o���i��f�՛e��a<n��b&[SN�B���I�-��:IJ{��w�W'�c��6�5�=��>'��z�N�p�*;v�`�ƍ�]�v���Ƥyhl�YL����g7���e˨�j4����	��}l�`hw�%1:��q��/�s���A��&�o���ҧQ��l���BUz��%06����9�Q3g0�
JTz�q�F�N��z���I���4��э�R���uJ�S�:b@L Z-ܙ�AU{�I7>�(�6��;F� ��A��4��G��x}�e<��Qr?�~."�Rr���c���Lm�Z�G֯�i�X��Z|mт����F�<����[�����1�a�!������������49���͈��?of������b�F�Z��I��v�<������i[���'�d{s[fp�����C�{��<�h�.Z<�{+?�!"�^�!�Xk�ゔP��7�%m1��D�4���Pkkm�+�(o�|���K3�ٛ�\e�R��"��7�4�4vu.��=\:U'j�N�Y0w]�V�B�^�ꫯ��G�T+*�5M��-�h4����l�R���&�Й��^S�1�l4�S�
E����`48B6�X���ń�֦}5�N̗��0��)%��o��)�(� Y}qI����:��y����~�㌁�\@�\�b>�;�`gO�����} ����q�R����7 �uk����͛7w�yVuí�c>��<��!�����5�۳�p�U �fVk�O5�[/�U��ߖܷ�������\u�U,]��s�=�j��0�-�v�m�r�/�a�ʕ��9>�Y�z�g>%���������ϊ�:N;����b��Y�ρ� ��P����,Ҭ���>*M#>2m{J��X��2����Xcv�Ft�m�Z�}����B�b;c�t�2~򓟰r�J�9��:k���Q#]x�F�e˖��h�}���`6v2;-v4�b>}a!�D'���v�	nA՚1?q����$} ڷg��Ўl�e8�h6�|�k_�9Ǫ��Y�t	۷mg�m����k`��EXc���}�2P��V�]w߇3�g<�i7��� H[U�S[Qx��9��v1I���eHc��P��`���ԞBl�i[�b�ݝ)��Q�S�m��}k�'�t/ �]kB� ��<*b��l�o|��(X�xq�߷m���� �z�Z���ח�{֘�3T�El- i�F���I�Of�HO�L�K��:�&���M����_e}���JŇڀ�%��l6���& �u�u|�j$U�����@���-m\AE𓊸t����<�7 A#B^f4�΀D�.H��va#��߫�	���g������8#�����4*s�� bQMAD�*��ii��;�B��j�g��2��|3�:絻;l��C�jR�
�j4
aa
�9�oJv�5o^�m�5-��m�fVҽ������.���q�R�KrST�fa���*��)�%�=��5�� �_��ϖo^��S/+5�U�V�������TRUզ�$GWb(YT�Ĳ���V�v�0�����a �#<�c�ǟ������L���/#�׀H�Z)V��M�B�@�o��I���<�F��y��g�)��:t����If�]I㡻�A�s�c뎤go���_eUE�rء�`C35��J��p�Cm��0���Z�|p���kE�ƭ�M��Z�U2���s��S��Y�b(L��[Fw��r�!�|��.	%O��_p�(�Ē�044�~ˇ����ֳXƥ�?Xe1沆��T�y�!��koW)9�%����|�Z�Z��1�]���Z���� O����7rB�XQV,_�7L{���e n�g�d���,ߟMDb���ZK(�O.M2����#8�ȃY�('ӂLX-P�T����f^9���/�[�mw> YΨ��l e��4�g����o�a����sB��Z�g�z��v\3���l������+i& ���y�9���J|<�rTeժU��ц�
��C�sn���W�\�D����G�:�5Cć�>��5�H14M���P��IH�^+W��
(lVC��G���O�+�K�p�A�r�@�jRzh�zba%',��Z���I�MO�?ѮSl1�s�p���Y�r��9^�����ε�.Ę�#�r��t�4� Q�Ѿ�] T�.���N7�3T��0�ak���Ӟ��04�~;=����b5`���g�����Yť��νO�X���?��)$�b{_p�6�]���J����爲�;~�6���)G)>[A��_~҈����z�Fz���U�O;���{��� �Y��,Ͽ�JSW �Ng%vZ��޽kH+Ҩ!���,)��bU�4�y=�� Đ���.�?�s��i@���B523O�骔`�������(��@Y��g�3 �'�/�ְ��*y���z�Fe	$f4�ЩG3��eU<5�32U%C �]9B�,�F�.��}g���!]W���F�Cb���]�i�6� tt�P�}ģ�U������4��ќ�:��m_��q�\�~�Q�p��(.6�9���C%�,T��&�q�_T筯9���y�[��Φ�e�9cn�Zb��TTlonjƤsqL{�M�.bB�h�W��	1P��)�G5�e)�-�*��ۖ�h�1z::!��$�*D�،�46���>�$�6�=��|1�Μ�&&`�4�_�&1q�b��1#�YҖ|F�э��YN�hb��ԤT�Q�Zcp2:wH�jzR��J�։�X$�R��Q*����kZ}NS��T����t��� ���gfEM��3D�1��$-�X���Mߛ�Ԝ7 �H�_�a��0I^�TZ~
m?�-}7�Q��:>6�\�}��"�s�P[cNۨ��c�1CP�kJ�!3��8�Z�(�TՌ��N��-�	��~�t��P6ɬ#T#C�<���m�Iz�@-s�䟂BDz|d�N���m�:j;��|_��#���|��}��`Dw�?hj0��`���12@�}�w���ߡ�����ϐ��m4�Ơ`&��ގ�I���t,s���~�8�ۀ+Fy����c�'#��́D2k(�֤ZO��h����Z���H�I>��n�=�p�_2����554hך�����mUDn���DS̯���H�l*�Gq֠a�)ť�w1�f.�E�v'o'����g'�iH���cLѝ»�����q3 ����:�E�e�㛹��W�f����v�!��+����7Rwv�s:���遨��$FҴ������!�)��|�7�(�Xu�o�m�^S�"�*������N��|��L����}ܭ׼�IWVַ�	�'��j=Tl�̓6�MUp5��1JŮ���� �h���i?CS��>�S׫N��Ky��y���O����k���n�y��N��j����f�
m��m��֚�H���7��v�[��hI���)�?��YÀ��H�B�h���B��>P�e��3��dh�����
F<D%�q2�G����s�!�������]	�kʈ ��[beg\H��K��E%C�T�-槛���3e�H�Z�lc�5�#^��G��PA2��m�	�pcD����^�_�ʧ�ylL�Rhb�.��~���j�a'Ӻ���`�ɀ��?ʒ��w�u۞#���6Cy�Fg�Ԥ�$Q��8��DlUJ�x�!n�滘��j�ܖ�L ��O $��N}*��(_�yI:>4���*��sm���u��3'M���s��0�����Ge:F�N`<tN�X{�(���1�����ʥ��ٯq���+[�ցZ�jj&�,��^ָ�1�i�k;sQ�^��w�w����Eū98��|�B��g�N��@i*���w�o�=�#t~Iި�������mk���2��UG0���Z�$�{u��ߏ�$�4�}�b�X��s�~Ü���Λ�2FU�f,*u��2�+^�ZN=�%�X$�Rɓ�\s�O���0Xw��X�E�A���c���S�{�$HN[ �5���O��ǂ��o�d��K8���j	�g,V؜�"�Ԗ�<��a6l�̶��“@�gA�Q���T����+��9���:p�2�hJ����*e���F��H�������3��H�Ukc+��IOt���')��B�� �60�X6����p��Nj�00!j�P������)/���;���^���:G�&#hW���!ѵ���4.-�͊���[�� UZ�e��*�Hϱ�aEQ7w�X4�A�%�"�:��x�9�io��K}Uf�:�`L��je;��A�E��~����6����V�Y��&�j&�5]�0Z,���ҡk��b+�5x������*}H%9�n'к��}�q��^��4��*�Ƥ>�]�RelRu{*��.�d�JB.��)���5�Ï���KN?�$\:F%ePb6�����7�|�V9~!�
D����K�z_���l~��,eP\�Q4�ጓ�a��o!��UA:�;O��h�TFY��p��'p���H(�g՝��q�0h+V�^u0��y`�f���~6loblF���LOTl�G��.b�ň��R��H��#_�v�Q���aN���`l����q�-wL?�]>"r��7�sAR����M[G�h�ӋS�ҙ��zp�F�su��_}g�g~����`�z٤�٬NJ*V�Am�Q�p�ͷ�ۜ2B�s�:�@��|�<�J3Z�f�\t�������׶�ؙ�4��8L�6Q��Rh��|f�U�2��or���aς8��<sMz��8Ь&i)c,΀WO�T���]�^��HG��G(�:TťZa�!&�F���0k�|1.#��R��뾃J�v���-��[_��t���i�e������c�A��2��*�0��X�
� ����㲞c�)��
����(�*c+F4έFt6y~9�����&QQc�:u��8��Z�
m�F�6�PP���Rs������Qb(RB�E�E�a����Rj���c��&�V��H�yN��Z�k�Y�."7;�3��H�`튜�\�)�)1��(B�G<�׽�̈́`:rx(�&�\��y����?��{﹅��a�9�B��9d���Y���75Aj���N���u�0D2-�q��O:��N8�A��Z܁ƀ)���08Aأ����ӹ��G���qn��"6K��twP��i�z]T�F��x۝�{dC[�pOQ��Ű��D��sX�a.<Lz�~v��|���i��I;���UGo�ns+.iH�R��w��YRH�,���o_t��-��U;�fԊ�[5��L��I)��9ۖ�؝k3�6��4}d��-\r�M�I�ѵ
X�8}|DŊ��8��5V(���F��뱚����?��]Cں_sa֚>�c�����i�iG���QF���;��@��p�T;���o���t�1�i^8����T�k�b�r} ��������AIAT廃FJS��ՠ�Yd�:�f�u$�4�\~��Hh�6k?A�w6��f]�ùeL"�{�m��h�BQ"/u�M[vq�s��d�P�@�M����L�&����4|��{��� -J.���,��v�rK#�b3����Nm޾�#����"C����{�9|��>ÿ~�+4� �ֺ&u��pʋ_����r��_�5�Z0�/�x�+_�o}��p�2�j�n��y������?�M��Ŷ���J$���5/�������2`�V����⟿�/\{��)[�1���Z�q�P��@�Q�D-���m�:�ż񍿂�Q��~ܴ}Ν�E���7��m|�)�Ĥ���ㄣbæ��dW'�ͩ���i&�X-rc�{��8|�br݊i6�Inr�
�v�[n��U���*�Yǯ`���s�u�� O)F�~� ��/��F���yFp�=�K�=ƈk�"���5GhNlC�Qm������@��ٙ/8�$��fQm*�R����Ќ�ԭ,�k�P,�Y���S��O�̮�8KF=�U�ݹ���HR�W�R��J�u}���PǺMO�a�d�S��])]�:�E����N��c�(<�e;On}�]
P�[�3Rl6�Q�%e�^�����;�Ū��
�t�F�T�w�a<�5����S!�Y�hJ)Gq�fCO�� %F����Q]:6��bS9�쁌V�c���1�\w�=� �j2*�@!�%�4Ɣ�A��;�iԱ��ظ�)$xjYb�1R%]�P5&�3:=�RU\hEn��8	m600PUJ�u)�T3�w1-�ִ���;0!L�����~�&���y��T	:ϛb�!4�gu�.��*>�k���x+W}��+�!`+����o}��8��>�E2Sc��!.���9��Y^��;�&0��q�������?��?����6��_���s�q� �k˖	��z</9�/�/�C���fv��u�3��q���RJ2��v5�,c*��2��y�1U�Zf[CG������!>��_糟��cV'���.�n
)(J���M�>��0�-�h�s^�Q.A�-X
j���K��yԎ�xGn&�Z���L��,⼗��o��
�(=Fv��� *�Sک;B��)��<�O��nMWG[ojg&6hb:T�����C+m��y�r�J�d��;85픠V$>�vy�ڝ�*HO���rqkm%Adf��
�b��7U�����\6���I��=�M�j�^#�uD_�eY��:������d��9'��\�m'u��XF����aI����T��h{�\�wJյҚlg`}R�sHL`%��@������ҀuI�r���"�+���q�"XIE!T�.E��1� �82k�0���:����v���P�Xk�h��T�hhC��	��97h�t8�|�$�Y�٘��W|%$/�!�	��ZJcˈWl���F&1�f� ,��J��:"�	�qiO�4�0w��7�ݥ�)�Ρ���$n��,����g �V+�M5�F0��]���=�pK���7n��h��cVrډǱ�{���}$�(�##򺗞D��m�r�D������s�Q�SG����'�����HdXu�Ny����;�L3�x�`�ߟ����<�?���s�/����z���p�Q|����f9!�l�1&a�j����O�lX�Cu֨�"5�k��ձd�
��$ϳj����
�M��>��+���i3��B��\XT3<UD�N�ܴ �U|���jz����5z�)0�:�yy�0�r;�VI����#jF��n�HQ6���V�0x|c'���x�A8z�R^�����+�؜��K��k-E��䤍�m�+&�pg��A�fIY'B��Iz ���Ij ͢I�>H("khG�*	�JT2��h4�1��HѤ�=�$�j���W��u�m�TZ�ځX���MC��pLb�B�f5���F�M'%��4&隯k���Z3��̞
� MS1�Jf�j׈3e�f|�x�&�U����II�؝�1Oﰶ��ǊmH�S�+^'�P��9�a:R;�����ZSIl�A�q�91L����I�=bPR���5����.�/
Τ �Wȼ�i��W?k#J�L��,1��̈́s5�0��z2-�}E�k����m��m�͞��fcz�
R�ֵ4���̸�XfV�!�=H�A��`���`�$=l&^�˾�#�m*i�V������ܙ���L�]������@ѦOz���/�����>�,���;i6v"�4�Pd�8��s��������Wq����W�	%�ŏ���B�	n ��n�����^A���W��t��	D�/��'\z��ٌ�RFa�cO�a�&.���T+�;���P�AsV������B�Kj��Yx�f�Z}���J[r�%y+�� i b1�f�#ض���T==5�,_2Ė�">ƪ��ӎ���s����X��+��Q��^�q��S�[qՁ�����Moyr<��Z���>�~�?)�j�!"v�؂���{�½��`��U�`����4��H4�S|]��=�8i�6'�y��ض��m�9�m۶��m�ƶ�>����W�f�5�s���g�r֕�|1��-[9�␈W��K̟C�����mh�m�è�"I[ψ^�(��70꼧C�:�aD��>o0kn=(A1	�z6�i�P;]2Tz ���m|����:����:E��~Xl��|����)6|��cvsL\�!�!4��E�?0m}O�ɥ�����y�UrC�p�<��9(ѫŔicj�00rr �xGB���璟"�����I�O��2�����١A�w����m�\\+�P~N�7Ţ,M�f⹕M�������6q�c�C�C=!�XV�gh��I�q͞_��'��>����$%�O[�vC5*�E��ڼ��e;;��X毯��)��e�X��G�,2Z��?�x�����щ�rN̸@�r��R�ܩK�@�j76����~�l�s�nd�8�����7�����~�&H+�� �F���#�ebLQkM�f-dh�I��2��W�N��_��wI��F s֛���vb}�R{�E�5����+��ez�|�&�����VslMly�-�v�$)�TW�}QѦ,C�!�=}�,��Hͱ��C��ǳuAh�4d�Y��g�1�n�'�<{�t�*S3ic��]����Z��e��V�Z߈��mc�����A�v_����p�y���oO�p�+�Ԯ3�@���	\����=��J��D�\��b�2N��;RF��vQ�#Aݐ� v`0;W�S� �O6PE�����H!���l%�Ь!{���HFʧ]�~�b�ul	O��*�H��W��&���9�����wLZ�Z}��K���u9S��j3Ӄ$?��!5{4�$��.���:4�bC���3�1]�Lhtg����G�zO�����)��|.?�{`�=��� ��x�I6�*�Ē{�T�Hv��z[�U i�/i�wG�힪����2��<E��2��q��9$�a 	j�*妅�'P�ct�mҿދ��M�ȶW*�@��m�Z�KA�^v��Ⴧz�"�l}749ו�R�ٹp��9��r���a"q����ǌ1�&~��ͽ�G�7E9෹R��o�K�rSDa���?��p�����]�}ѩ\�J��tn�8E����JT�%�@�����=n��y+3\Sc�����ף+>�B�AY���s'0�&���EW��;G{�E�9��	�]�l]l�������K \��g3�����!����R�J2|�E����18l��J���c��w;�D���g}�~�^#����>�Q����CsM	
 �$�Lt�Nxuףn�8�Nf��W�ϽG�g���z|��QV�QԬ���u$���%i�b�U�J�΀����� ѻ���f��I����\SJ�387�n��?ߏKt��������=�[b�f�1E��/�k�OX�3
ć��_m^���XI���$�Rֈv��9�afͦoĬ�l�6okn�MО�?�5�b���IԖ�z�˕B�<
���~Y��L"9�;pM:	S�s�|�9{�u	������'1���n��bU���S�O��E��,n����nuiCI�l�$��G�,�e@�<%��Z�h6�rVRG����W�5=" |#����7�����R�#��oڟ�R;�7�/��<���C����ٴ����G�����WW �����>nu�����O��Խ�O����nu�+��p�̉ҾKؗ��ڣk�R�\o��B]zp�}�kܾ��jz�:���<f�n��$���0N$z���r�l��,P�<ʃr�/�V��?������~\�r:O�f�R�J������t��c�o穾}���3f��{��їW�eL%9��B2�='"�����6��׎h|�����of��խWO�:8sb6.�pD�*�4���n��P�`>���eZ�#o�B)��U���bwR�.�4������KTF�xN.oyK���4������47_����e0�>g[�����ā�l���z��T�s�����(�H�`lT��AFx��b���Dh�l�TjE������V�G-�d�u�D���[�Y)b�/&���m���>-�J�+-ߓ�x<=$�Y2��J�����t6�(s�CPX�o��
C�q8(]p�at	4��w�(�� �q��4{�z�
�TU�P��6N����m��p�������,U9Q�\���V�qg��c��S�J�ºw���^ ~�"��h����{7_�[{�F�B� ���ĜA���Ai�t�)���0 Aʕ������jB#kľ:�WٝZ��v�n�8u�k��EA�ˌ�"��(>��ޗ%e!��γ�� k��nE)�;�E]��Τ�x;s�Oߌ�ٲ���I�Ӏ��u����)a����$X:KYǞ�v�K$��,��b� 2ݣ"R@ʒ�研�K�W�0Or�M7EC��V�vu���*�F��妕zaR�L[�������.��+��_��F[(evx��?ʗ� ��22u����Nl>�/`�{�O�k��:��x	��=sj������p�m�=�Ɩ$�>���ck���f�ӵް�+�9��Ę	1FPOa~o� �iN	���+/�ң���Dy�0��0���YA��l�e���xS��5XN���#qe��!r�B��_��>2�Y�'��Gs|DI�e�N���|w=�-�G{��큅�hҢ�������/{KV�{	D�cb+�j�C�׆��%�ls��b=�[���]/�[��L�!t5��y88�yi"���r�E�7Ī8f��E\��m����s�1$/J��XbWH���#0��痞Dh	�̦�s�0b��b�����c��aD"
���w�>f�r��u8�֢���p��V�+�S���Dg�(Uw��E:�~���:�9Gk��0��rLx$&�`��EȐ�MA��{���F������뿭]!��:`��)B�+��R��5���)�'����V�a��O��6E��Qa�z�3,��Z=�k��:�sJ��/�m�˹Nsj�H����|���gR��mtT�E��@�Q��5̅v���Sī���Vb��'Sڸv#��C�r�@O�b�46	��/:�Z����~B, Mh��c��:�oy��DBKbU2Z��[�,ʄ,�d�D.�sׯ��eX���*[�(��?D�d،Ϫ����CV6�y�|h���ָ�����f�Z=���!
����G�jwJ�6�����.>�>^�>s�>��x�l�\ԉ�R�	��{?Z4nB�|B"m��:�:e.<R	Z��?w?�>��v�l��и�~���~�xl�l����׾�M��/[�u��x?pY������<}�k���#ټ~r������S17�;��?SܺE45F3�a�'x+1���Q��w�>0Ȑa�G��8�ܐ.��ƈ�6�� QnccP!ٹ�}D���-�ۆ�*}��ye�RY	,���;�ϵ�sUUsȎ|� �(�XTq�yi���[5�y�|-��L.o���^��\�;�͗�[��'lǻ~+N�si�U;
��}Y���8�;޷'�B�KX�%�����ȼ�'���ӓ"�x�R=#Y��2���э��k�����<�op%�3c�g��m��qﻀ�B*���!/M�]��<xd�-�8F_h�6��yĒV���1�о����kHW�O��ϏKk�'�*�3|Jh`��ǣ�U�;Q=etx��r�dM"S��j�;����5_�oK�,w6M�px3�p�B7���.r���?�������t�cEO=x۞�|>�ȝX�z����$(��Fx�I^�ɉ��#�^��a�x)�:P���2���\�r"حj�l(�?6�����<�u��xX�{��6r�I��z�G�g}�*<~�<I���:�w��.f �� �������C��Y����>�>��%f���qS���f!qG���.P�.7y �_DT7��у?>O���ԊF�����Ns;�d�M��N ���4�S�xWu4r�N�I4�d�d�5��L����[�%�(�q�.����q�#�o�D8�¥l�� g>��g�A�v�=�RL���~��V���������m��)��e�y %��
x�����n��bslƆ�FK�=��腙�iO�M������2~�0�.S��H��E>Y�/�Y�]�����������Id�a[J_��J�~�w洃��o��ЗìHXl� 0�!8�qOg띑�MeА�_�#J�6�MA���%�h�}��Uu�QZ�����m��F�ϙ��>��z��(F�a'��]t���`�=����usT)�Q�zUc�m���a�m�U�uȋӼ�-2^�{��y�lv�ؓ��������H�ܗ�~��vx=G-��W����&��*{���H�D�`s^��ػC��Zo<��C�y�>�i��$����F=���h{�bxG_Qj̀[Y����,9"��1^RE�����D�ȵZq �ĲS�����@���xARW�?����CDàVw��x��e��سeR�>w�ej*���� Uّ��f�t�/�����z�^*|��AL��jUZ��.��&���j��n��*����8�N���&_B�j����S��R#H�r�����,C}'A\��{mw��51�Ϋ��>:q.
��t�p9�����%���#0Gљq�d��o��=��ba��Q��g��-��X��+���JMzh���^���~=N�Q?7�Qs}����1�OÒ������)�s�Hw
�{a�c놪)�Ȉ"�!�X�Z
2�TJ5F�{��${J���d�U�g�@�7�)�7@/�m��ګ��UҰ���?��'�e�6���"k.!��6���V�#-;���Y�*DH*�8!i��l�r7>��x�8�q�=*�X1�x��-��>��6�ix{\����=����(���[������\s��#E�w� Ux����d�"�P֞�T������E%�A���<���$� �T�z��=c-ySK�n2'�  �k��WZ��n�֤h%�/�qc�������\��t)Uf�x�,��-�x��7C!�윽Yb��d��.�G߹K��}["r���VK�o#:�UA��Y����67��\����D����(S���;�U�-�u��H!'q�-���h���L��-�\-J��7��S������ն�^ݖ�5�E	�B��j&��1C!��R��� c�@�:P�R)e��Vc��-˞�}Zl���J��qB]@w�r	��%%�Z9��W�o��N8VW󘨣�S���aɰ##����&Hр`���kt�ͩ��P�u�X�*�I'o��!U�ʅK2��Mv6.Ya����2�U�p�N�>�N�9��i��GM�����2��0[˽U�e+N�	,��ƼMNb��hh#�D8O�f=�%�=w�
�N� ��N,a�`yo�73��� ���RWv��2��H�8� n���%�����i�ѳ��+��'^T����,�lO�c5,Wt�D�wd9�M6����Q��D8�a�0��hƓ�ݬ�yP�5�����=;���u�+'��-��$�2y�)�o;�p�e�"��W]��Ū�dK�e�X��h����N���ɧ2A{-^��`�	�w�8���D��Nl�j�DS;�8�\Tn�%v#���ߞ�����c���]�iQԔ�`N�U��!e0��(�gYF����ilMds�pj��]��	O�R@�i�n��97�Z3B��������!����q���_��}��ބv�Zt�|�Vz�^����Y�;�Lr���gk�����,�hc��G���)�%�����狙��g��t��p�_����i����4��%�H��OC�����'n>j.�h���~72�o2��2����7�����]m���0���TI��S���Qg���;�t<~\er�a�ogxQՒ��+h��$1?�Vi��L���GGOU��U���w���e�k�B7Z�g��PKYN��G��J�Xo��գ��?���KWg(�b�B�V��WA�@�'T2���W�g�C���I�8�����W���&d���E�Uu6`a�3&D~5�-��*��$�gѡ�VGfo6��d��9Zs���(#��ӄ�^9A��EOn�O�E���π�KBN}dfA6w��g �W��>�G��$���<�FM�Ǩ�kX�w���f�z����v 	�x��0�/�Ϥu16ѮX0�,�P�#�DP�SFE����C��C⩯sk����,�Ng�:,]��+�'���V��<s��J�l9� I�*���Y[���Ķ�Z��9|�fHR����O��l��{���;�2ԅ�(�m���(VfN�c>��#C��o�W-�~���TX�Nr�k��]Z.y�8;�9B*b����*��0����3hΟ�/B�[�xϬ^.A �3z�]�����3�Y�S�i�ȵ�����q�n����C�籡ds!w6��b�:��=X��hTψM4���c�ƶ׌ �Jk�.T��9��dJAE��1\f.�A8�ܲ@O�)4NA��%����$B~��*��#����WSq*p�客![�H��D@�� :��P�+��|����Bq4ݬ'
;�,���>�^��A�1L�� Y\���-N�-.3�Ы)���&��"�ڨ\�
�|`�d�'���}���.��0�s#y�yR2�r%	IQ��z�g��2�p�i��]���SYz�k�nS�F���$-���� �+��Y��~�-�Ữ����q�k���yY�k��gRg�kYګ$*AC����E�\r��Xྡ]��g����쭒kK �s�N�J%0Q.����6Vh�d"&z���Α��T���?�l�㹯ew�Q0ˋ�yDT�V�|�h�2=أ2t��$����lq/*�v�_��&͠X�t�́ͅ$<		*�0��-4l ��E:Z��Y�LӉ>
�I�S�-�ʓ*S����6Xoh�X*EKUFT�����Eٶ�vdw�dx��E�`��.�}m�l�7h�����]����v����Zx��� 偛N�1�9��
t��"�>��r�.b�`�Pg�t�����w����#��UX��GC�9���=�,��̿K��P`�bH��p3��j�0�7�mb��n7h�^3��$Nߌϓ��"��ҍ,7	����䜲F{/(�&cȞ
5|�W��<�>��F��oN+2e��I����:c���TФ��#|O�چM���� ���>�N�i�j�m�P�:Z�X)�\#���=d (���+DB���U+�ג��1\$?�XwbF��q*��_`��Ȧ�����+��͚u��O���B))��k\0ڳ5��d��I����(wE��c���S�CM���[E�[�t����&k޹z�E_+�p��=�������k����/�v�f�${�:��'qj�'h��!Ed�M�W �a�jYw�QcY�~\��G=�-_TW �T������m��yb�7gd�B�QUb���H ��b��(���_�8Wss��cyW�or7�1yyQ�N��+��ۇ�����Y7n�,��|a�#+`��l)Qv�Ql�^Ն����i]|�+���$�QΕڝ��[z�f#�ʹy*Μ�du�⯡�?̱vLO�v˚���@���l����'�3�*�'�2ݮn�.w�F ?Ӯ��T��T�yy���*oȡI����	)��r%�Ё��4�a�H	�7͸��%�$��o	|+n�]-��5�j���\Y���V7NÍ�o��_����^���*���}�kp%@ܫ�-�WЛ�Qb2�qS?O�
2��0�ٲ���Mq*��j�C]?y�^�M֙�[d=$���_�_J���o�0q�O�|e���Z_^È7fZ{N(�L�E��H[R����/�_��2؍�#��~'I`e�豲�����:��Y6�`s��j�xO,����y��d�0\#v���w�)���@� �4Ìk��Uǵ����0�un�m����g�iO���Ն���·U�W�9�G�L<2w�^�U<��':�h���f�n8nsj�����us�9;~|<�������T�Lӧ��H��ӘW⤖H�q�����-3�:�x���~��Y�P����p�C���3kqUW]������t�$��N~��붵��z�@U=�)�z�?"eS��0����i�2[�o?;<��	\e�C�i4�NUC�<�e�-=牌�Á�>C$]Ge��N��|2�?�`-S�IGZ`ŲЉ��/ (�Wh���#���@=o�������mS�a?;JdO%�P��Z��o��tW�t���߾����%����9��$��Ԝ���_F7"�d���#:��h1���R��Ԁ#h�0=��#%(�|y��:�ϟ/���C�`��o�����a[܈B�28�y�� ֙��*.O1	�]���w�N��ɕ��j2�l4��ސ��:�DD;7߼�������B<�CG�>`[�S��� �&WDs�1y��vnk�Xbiz����lF��/�/\]8�����yi��������zZ ;q�6�ʹ?��8d����@��-�\�HJR^�����Z!{�S���x��흆,)I��r�aѡ��vFq�9���[lc���? �<�Ѓ��6G�益Y��G��-̣l��]@C��S�l�� �I��|�*()eg��#4�w&U)Gt2d�zT�#������M����@��Z�[CNYy���)e�p���l"��)Z�������!��/U���oC��	\���V��Z�"��w��p��R7�ؿ��̯!������ڕ<��o�95'EX���0�n%�[�^�2�zyZП���zs��=!D�g�8��;x�`��jbp�p�^)�Q�P2R�e@�����lR��q]�(�����K���yJ��I���/E��&��Z����27<��v�e�~�j#��$e�`.(��6�B�1fI0<��	��^!�)��a��;W�gx������F�f�[��K^���d��%��[����i hu� �j��k	�A8�b[G<C4���ҖK�=̵�˝Q�^<\GizC냟�߬G���ϐ׭��l5j��
xD��hi��#��0���&�^¨���\�i��Oa��a]�.ht�9u�źF-4ڜS."Xg���F�n�ئ��ُ-8��m����U��3���n��/����u�*�2V�锚'0'��q[��~�(�L�K 	��N��G���^�� u�!��6�@��pN���cb*�gޜ���/��5.�4Vt��񿇣24��L&�^���8Q����ei�A������"[/-a�hW�+og�i�²���v9�λ�&ck�BI�p�P)���Ű�ʡ��0�O�M�������9��T!*l�>��s��K+�������أ�yr��Pܟ1��l����3	��7�*h�BPP��^���B��1�����ϑ�����:J���V�7��gZ��(O"���^Irqx���Qڸ崝Ti���{��g=x���7#G��+��h$�>HzOQ��ڿ:�w!#G��V�C_�b8��<޼�j��Z��~�&TDu�驉R��!�����*�i�BB*@�� Z�yJ����o�[&���}C�2��cU�C�䇚��J��6�D>A�W �`R}#Z5��\���"!�!}˺�wT�iS@�x��������ǐ�B#W�����K�,|�aW����A��=T��-w�W��}mu!�F��'���G)�yMf��T�d )F�4n�>�'�0]�^gS�=�Ö��V���έ�E
L��7bR�P�r%.�r>���GԸܹ�z�8�K�Z�/-�*�t�6�o#yF�%N�
�?2z�I�o�A|,:]C�*�����$!��/�an)�P��:���0v��u(�a8 d���`M��pH�i�v ��ov���Rǣ	^`�*�L�Vt�F�4�*�>&Ch∹FϧnT2臄&��U������C}:��a��ŀ)��\CG~թI�B�J���4��aX^����5V#ڥ��d�仐�/&�ME)xQj���ӷ��qWh��̤E���	�(fD�Tp��w���;�����ј��e�9r��Y 1�Vy�`!�p���W_�/�)]� i"+�`C�2d�w����#�]�U'D�Zǐ*5)�
H��-cU�|7��4��P�T�#M�fK2P�3W�:~-��z	�>��y�R�r�[�QǱ�O�e-q��U��B[�f1+��-��� k8 *W���ӽ��%��I<(2i��N��Ox��3��F��5�Eɭ�_KEN�⥨H��϶tUIS�ܘ���(n?w?��C5�yT*.���T�k+4�\e�e���i�E�Zȗ=�qO����}I�#��6��Gyr!`�lV��۬���c9��:9DG�,:H�( <(ch�+bM�[f2���Ŧ�Y���̸j|�s��������,��&�i���I��h]�8�h���_�C�{�����~��ì����q bZ1j���S+[�Q���4��!��ך�D�����4��=:loL"(Ҕm���]E�Y_M�z�a�%]��s㵳ř��L����~�y{L,}�C>%�������S9��++x�=�n.f�VحSZt�g�5���T+5�xߵ���13�Ʃ7�2�>X�z�h�}��U�����z����;�r+��9j�c6(*�zn8�JIjx�SD/t�u�5��f�%t�.�R�V�[�NV��?���2�v�!�[�6|f��Zv�$jc�Bm�F�ݏ�i�����U���M�K�cXvRU����]�ixͺ���??b���ĺ��j�\����p�Ǭ}����2Jؒ�1��>�p[��`��^iW�}S�ћ!���V��/���xފ��T��؄��類G��������a��`��?Y�g&g(i�,$��:Y\��'�&x��i�ՆeޙE�����s���1'�:S����"��5��2�8���JF�	��d��p7T����&MKM�X,U� ���QX��^+t�h�C��bCc�;�6^U|�̂W$�@b�M��	�nG�dj!J�Y`�P���_<H���5�/�cF~�pI�S������w�ΩT�����$���������.�q�y>��� p���c�Y��'ʭ��p����V�GܦO�1��z��<�����k��5\:/:��\�����\�W��Ui:MwG�N�,���,��~��;7'LXq��.�6�p�H�A��#�(��u�3��_ )vϩ
p��i����ǩ_Ǳ�T!Y����ng�Z��ʡP�Ш04"_���ʀ�/%��� ���#��9��N��ɖ"��	Jq嵸�H0:ﳺM��+݄�/�X�C�?�4��)-���P+�=Y�������%J�	�I,��sn�B�x�å�*H�;[��'+������46��}��k��zO|������Y��]ʹ��ll-��}�3i�.�gs|ެy���SF�������f�-%zu��}��^�}�y����4�s����b���w����%6z.N����� �>)~�'����ۤ;���i'�	x�
�y׳g�����eQ�����mԭgJ���,iKV���0���n� �������s�H�Z~�{<b���3����<3��>�F���"˓�l�w�����Kio�-q=�ᓹkw8�f%g�$�RX�o�����J0�ؒ�3�~���+��
GZ0e9�Tࠫ��P,�9�'S��A�Hf$�b{��h��6�|>Y��6a��Z8�Ѽ���#�]���+�!�˥��s �>���%��~-&���v_f���|��]5�7��YgC>��>��~���m���-LM:�\羻�e�G�z�H�E/j����E��8?�Rx�WqY����3����΋bE����f�`}a�gݢ�(Q�8�VM��y��Yu����F�#A�fFw[�PM˙B�"j��
�7��؋���dK�6��+R2}�V�~��%����=�eeP�Wᓤ��0�v@ӇX��M��Q ���y^���D$������a�.�,��&d��A���l�	�}PWw��v��Տ�j�vd��Q
��φ�cg��ށl�.���͌S%8�
����e<_�/�eqi�����/�b}��� V�����[�F��BS�i���#0s�������7Y���&Ya5D/:��[�'�k��r_�V<����3r��α�̅�-ς�IY����#p������R��X�Vz.�D/K�;I�)�<�������[��2'2؎3��f�'&��M��TA,�[�MX5�ۇ�"[6����ԭi����D���n�]������_��Z�Y���=5�G?a����.6�u�ٵ|���p,��誤'����7�@%��L�l7��L+׷ˬz���4V-o7�M6(Y���L�į�a����)̇�,�U�U7���Am�����\2����8��y�蘙C�Y����ͺ��rEH=�M#_<�%�po5C��{ ύ[�R��#��NәՇf$�|�/�H�	04	7���X�]و`�QFG��M�W�Cg�4�æ�(	�!|���O	9���XG�i�cO��?������}B���Q��4%�u�~uy{֢���5�?�h�o�ӎ�ƕ����M
�;D��@�*��tX��޷u7 栄�9�${�4��9�9�L;R䶵���]9�E
����Oo���B���K�;�]>�u6��g�]�� U�ImyA�Juz��$#�I�b�h�J*�`
R]N��E�}z�������R?��ٵ�XG���=Q{����=D��7���('���W6���\7��=���\G��]����Y)M��x��"V{Z���@�Z����ke�@�ř����,��~��u����?F8�"�
�\v\�:*0���������;�X��B$��o>����~����C2�Ay��S����J�Q�2?c^��X�%M��o�88@�ӌ`���E����,w8���q�kg#�ь��,ؿ�6�/�5���=�V�F��c�آ�_�Ɓ�h��x&��E�!!�q��Ub`E�J��4���:r���\��K���GOh�:�p���#/�ib^���Z�W!Luxx�k3��=ц��=x���+C%���mH��-j��M��1�k�Vd��?Җ��s�����	�B/mr��P90zD>�:��ꤨeA'p��xS��+��s^>Y?����p?5k���'������+S"8�oI�3���	(yR��%Y����t� �x΀��&Դ�3+R-����ݎy;�A�9K{���JS�臓�^Y:9���H��v�(@&'>C�|7*0e�h<;)�'�J�h@�*a��Vs�ڟE����[�]�$c�ͩ��A�R]�<�[��p{HCx�3}�]�g�ѐ,d7\cZL�V ����|k,��Y@-tm陀���{S1�E�}���rR)mL��<�[���	���|PJa��KF��Fr��#���Bg+��C�G9������9������
�#M����g��t,ՀjW.}7+�:b���d�w:L���Ǖ�w �7)Y���&�T2u�BC!���3�����y��4ֿ�2��j��KE޿'+O�\F�,�Ġ���nf��q��u
��?�xzi���������<��(��,`���=���7(C)%�#)��ϯ��6�����o��E�%`��!��U�r��~�͕T�!��l w���w!~\o���#���o�UD�Fk�?5���>��go�k}�
CY��n���A����=�
���~�L�O����F���]�7���_gl�A��[o#�.�r?I96��@�s�BՃ��]j93�|?;=>�+�1��&DP7g��]W�΢r�=��xe�����~��6 �*gT��6N�;��,7fiƐ�Vy���#c�Y�nLS3�%5P37��<E%B���x'T�nӖ.A�,��dmK����#t���.e�Y�G���H���9���9�&[������_�h\ �Wf�!��7xJ$d�Bݯ-,������L��ga%�d����OU'x����|��v 	ݽ�s3�w��m�ĥ�2 �BJ�#h��{��7G{����N@�@f���*�j��v�>\0���q���H�`I�q��.2�ٳ�T/ޒś6j!�����H#{ƫ����O���l�{<3����C��&�Ps鱊��f}CC5�ӵ�]���"7�]�Dܟ��QA�pJH�ЇP2���aۣ��ߍ(\���
1�%nu�C�4�<�� |���v��!`}�ī�~��۹c�c����l�C�}��D����՚�T\IGbt��q�~X𛮜�͆ E���~���g���JT�oD���n�jH����E����9���Y���ަ����3��(g�r+P��������p9��4���~[ӁF�0M8T>l��h��\�fG򹨔d��k�*Q�Յ �UU���@��z���5P�-?\�w�e�4������; E�����1���߼P��/p��C���5�`=�z�9>�Q`_��o�[1���{ru���/j˓u�U�Y�ڿ�8��#\Ln�\��;�B
�r��NvE���_��R�+`��#Lđ5Uw�"���]�JA.ֲ���u5���o/l���>0��ْ�Ҽ�К[�փ-���L��x�.���H��З�<=q�O+/3�;|0�*Lc�yz��=�j����ȋS�+&�?��JcQ"$�s˩�g��j���� {�P�E�0V���9<#�������k"�)�.���os¸��D8�����WXՓ�*�C����Q��O��[r=NY>^s�K	����^��Q���)�f�]�\T����7����"�q�H7f~/aY�S�
~7��{L�����c�pN��zw���;���q�6��[���{	��X��-��/�4���E�W@�A�K�&^ю�@���i��?XUe3�P�k�JEN�-��g�z��D���t�t�2a�J2)0y援޸p�� ��L��{���8Msa��;��b}���������
r	���2�����\!=R֊Wc��QL?a��f�j��!�SG��<h9��HǼH��Dh68�&�ӣ����f>���*���K�Ѳ��ͅivq&���(Vԙ������(}W��a�?�V��B����&ӯ)$b`]5�c�E�M��2����BvFf���נKb���ykp@?��|�ᠷ8nD���	��ur�ÄC��&���Z�n��$xD�R0�pQ%fo�}{��o�ņ�7�-)Q����4[Xr���Y���R�'��%�p���p~��*U?(ҎE�c��k��0����5���O��,	�)�GV�)�a�LI^RIn�V!��
��?��DZL���JA�	;+�|N6�4��"��P.��b} ���S_�d�,6ɤ�?v�1˜%�P۱�G}s�E���3��e���y�Z�����1[�r��s����-c����~>��W��V��T��%c��h?�G�/�{'�Q/d=�����]BA
�G�L`�������l8x��#�Tj�Wp���O��k��h���_j(s�^v�fZj>~���Y^���֦hY YZNp�S��e�\ھ��n"G�ḁaY�. ��@�ho�c�~X`{T�Yq�gvٽ)��u������kc}�PYW�u�op��}�N'?�S�?U�M���~��{�z�h.�M��s���Z���^�n�m�K�e	qDz�w�Faja���˒qaCxhU�H��_�L�H�X�:�Nf,���}�)��򌈸��W�٬��:�О���}���]�,��Cc�@AG\� ��R��8#��®7�Q�og����o��$���1�%!@�~:1���H�QH��m���3�c�Ldc�� �}���������I�bC��K@��!�2���x�{�^Ms%�{6�G���k�w��m��w��?��C6�G}u���"�xV ���,���ӝpR;��L�a2_$��xQě�V>���`Y�h�a���[�6�Smwxj�����Bps��"�wg�c���Ј$!��sh�m��6���$�{{�8ry���¹՟����2*|fw��O����#�0V��U�x;u�s�?v��3`)��;>��Ie�F���e�n�Ņ6C�ª7�1L2��;�W�բ�_c�a�0�^��-U6�l�lu���Ю�?��F�1*Ս�'���s3�T+���}�kz\�j�߾�^���o���i�pO$TM��x|����)���)�:h	������:�Ƶi�\�vTOk }�Sk�n����,��j�(�+�����ݵ�Cqw
��^,��Cq/n�����ݿ�3�9��k�g�$�&�qc�`�@O�^�!�=|�j-�6�m{ܱ���U�L~�*yd���28ß<6���rR�8�� �X���Z��$K�G���83j��o���Ϊ��7���8aQ�0�vj�q�[Q]���U�ʖ����H��`���(���c�n��.R���z�~�N�ҞUb5Q|��W8�zYp�r��ß��@C6-W"�fֲ�b�4g�=�!t��qS����"(�6��8���Q�.��ǿ;r
���28VL�˞w�V#���M�zk�#x�}��1l�#k)]�TY��UM�p0Z�F���Uv�)9o��9�&x|P�O99?A�p1�Q�Դji:h�	�z	D��c�1\�����[��z=z��[��u�y���
�#3m!����S,�L�h4�o�$��
~}�� �0hL�qI���>k�ZI;��o�T��t/�B�^]ElD���~0���X�uô<JV4�飧�����o;���������w�s�Y>���d�;���z�צ���6�6���ۨ�jy��1B�:~��3����R��CO������Rؼ��y�7�2.�<�����Pn��sl���ə��&�����X�<�>��Q�,v^�bW.%��w�dM��e�q��j淋V �[��.���ec�	�h�~�f4p�tt�����C�4�)G,5���K)�t?%t=))>�$�+��d?"9E�W�~���7\"��b�FϤ8ЯV�L
�hN�v�]���	�ݜ��h���~*�$�@Z�PZ,�Y���Jj��W��l�
��F�hW\L�q��������3ϸx���E`Է���&:��7!BUM�yQ�[F
�#J��#��H�_�!� YS-��'>�!~htbԾ�4��z���a����Ð�~��)�t�_2ô�:�|�^*�Y���H
��F�ɫ~�PT�mi/�	mJ�q�r���IOZ|
��	�]��
n�#�q�S��'�Z�Kq�S���d���e�͹�K�!$����N��t����vp)��5���YIE�s�n�8���U~
���m�V�+�3m�5st�V밼������g��j��Z)��;�t��������g;�s!��L������|���Q�8����nM�`����Ez	�|kuC ���VjNB֜+��HR����Bog/_��A]L6�&�Ro%]^$��u��ޯ����_�R�"��0s�lUHPM_����	�ÄF�Y��S����c�b������#��V~�w��(���Y�@L!���>�-�e�}���eb�� ?9ߚ���Q)L��������ƺD��Y�r�����ju��� ���փ�婜�7T�o�|+N��LS�b骮{朚��5ۤ�v ş| YF���Ԕ`��=���GKq�N���ƛ�ˎҢ���/kF����I�
]�i����h~(iu��tg��*h]���-���Eʛ�j����ˢx� ��km`Q�MZܑ���1�z���4��4���P�<T).3)�A�)����8|8ố
�򔋮$�xo�T#��.X��8����N�x��u���%ܿ�� ���%
�V��� ƃ�T��Aܪ�C���a���j �j4<��ݑ�/���%,����'䊢*@�{HF�䐄4� �ݍ�1�J[Д/�adgơ]@���A�� w���)��Kͦt!;��4���C��U�^�i9;+�I�vn�~�qbM���K�����OU�j����(��v��R\�E �W�H	��&f��}e5L�y�tj>��ƈ��%��������~-
�� {6Su%a����U��x2I��� ?!����̻�S� r)��X�߫ٛi���q[��鹴l���(5WjUEΨ*�<�����,v�/������Z^�1�t�h{=���iP�EG��sWBB �~��ߌn���i�@�yu 0Z�-<��j�_�!nN�$�)�dҡvܽ���S�_��:CǄ���Ud�].&ߣC�)j$ЊD���# �Ms�2�¨��SʘaF�����H���cDQ�4ã��ن`8�0Ժ�
�B�^��%����T�=�;OZ��$�'�YF~�nE�����M��>���z2��׆�x�$ؗ�"�i�w��H�v�0�@:d�"~��p��D��� E8���\��z��a4J���ȭ%��aX��爁,5�gg�DFf�V�Sz�3��(��;�����	�/�nXdd�����`��k���YG3W��5���}I�����١c_�@Sz�$FS�N�17��� �)��MX��]ު\�iV���uRY�����
�B���|yM���� aP:�9��`kb���p��L��}�Ho������J������(ɪ)���A
�ʾ� �3����@�ݖ$"�P���Dw
��Hr�	�#��W�\܀v��x�V�Ի⢅m�\QΠ�(|�:����Vʽ�?/JD}���������nÉ�ym	�$X��G0���7Y��}Z#Mqf���c��fu�M�Y\�v����;�:a�H*2�`]iz��)�"m(3�u$����@�Q�'򲌪�@Y|�C�F�G��4o7h��q�5��4��`|���X঍E*���~2o[�<�D�x�l]٧`� Gx�qPè��On�z��KѬ5$��ϝ����
����eky���v̌	�+��;����S��������D!�cܠ�Ȯ�4�E��Y�� :4���"�{�Ki�ݟ�můdF�*����P�C9�O*|�z[�k�7�:I�^!��T�s��Q'��Q�Nu���٤+Gȹ�YDF�%i�
��4KB'����EV}���L��u��%���׺k�Z5��B���+�����Ȗ�V����睎\j�q�R�g	�����Ǫ�A��ɱu>U���33�� �4Ms�NP�q��f��4&�/K*Wf���8�Q����e؊_m �#�'�{uc,=m��I��UWM�5<}ߥ5��8!����23u�z����"�:���Q��[3��z�U��/�'[��PW ¯[�W�<���^��%0��K>�X�RS�,AѩB/�)����OX�oN���2���[����ykF*�K��k�G_Q�L�y��1l&Uy�'��r%���tɺt�OȅK�!V_�Q��T6W��J<��C���Gp���mZ�# ������Z(�|@1�B�|貴�����@ׄ��%fofΌ2W��8�(V�c���bȦ��%�\	�p�߹����]Q%(7�~���1�J�Uo�	||����Y\���#�S�i��9*'��H����0X��{������ą9�����6i��)��hlٚ�[ZZ�(�H2%�́`�o�OJ��:�0���b�\X-��E�������S%p[D�����r�qHf�����o(^�]N�`�oR}�;Ǻ�m��(O@�jk�:�O��������蹫��l��B�3��?��7���Π+'��A9i�y�X������	��{���An�p��ST��])�e�R���x�,��L���=���d�M�����ۚ.�ni��a�Mdft��b����\ε`�<��\������N%��L�V/�bb�0N�z�� doG��������r:����6eg*��X��`���"�d��Ĳ��aґ���
(#���9u��g�7$>)~ٜ��������Ȉjhv��y�kqcbU�0��+�+ԣ4%�Z��������o�>��d��o\�F�s�#S��q��% ����&z����6�C��(��gBM5q�ӱ�+-�C7�5�{���3i �ȍ�kzh��W	EZ��-�7��5����.�a�H����.�P4�����)Q���{���gu���5򦉧;J"�Ec���7멀�r�9w�g]n�7��")�&h�k�����U�g>����G�l����Bs�=x�Hޯż���*�!D*]�����(��*��|̍��]
P9[��{(Y��1{*w��NR�,��B�$�W�������xb��z1�!N:���e�QT<�mY�c��0��f;��&?WEi�*�Υ�g0P+�������Uu35$���M�bu=b��ҋ���n��_����hj�W�ښ���V� =a<�~Di��~
O5]�`��>�8ͅ�k������|�n�"��� ���ټ%�(��JN�|`F�q�]bd����	��U���'cg�e	H,E#��a{g-xl�i�
������N.����s�p��v��z�e@_
*Aέ��z]֞˖T1ر�lW�^��²��	��:W����f���<C��b�mvƭ`\<����3!In�{e��z�~L�e��h���$
8d.G㧄Ss���]~!��#����l��p]��g.�Ǧ����10~$I���/�[�G����C~��%v�D7!sQN��+��dG��ՄGD�4���;riJ��ک���P2`Ɗ_㽒���]��P}�L�L�5u:�����`�,Eߒ !x��C��@=�P�$�I~��i�wԞ�*�>4�OVyK�­��x��K��zrѕ�Yݕ���Ƶ�j�e���蚺l�������7/-����^[׈|�T��ݘ�D�U�D�%Ҭj{R��\���E%����.��������s��oMdYv������:�dH!*y;�j��������#����ah�X���:Wϩ"�X�����e���1���F��W
AQ��܈҈�`_悑���Z�����Ɉ*�J	I����~���'�i
���r^;>�'���RF= ��ڌh����#/j��8��?H;��K�K�E4��'v��ܖ �n"+at&Ӂ�dD��Mi�ɹ�O�e�#ž#6QÈ�`U.{�Y���R�*�e�����O�q��:7�J�P�]�m���,k�H�뷑"�z�[��%fi���e��3�uL�(��g���}W������e�uE	��B���cB�\�1�`�3�cn��U��J�>{E�b6Nhһhi��ZR��:�a�!?61AK/��H��,�I����4U�K�b4]�l\��0�9���6F��#�ЄJ)U��L�NMGi�,���Q�2K[���%'����P-:��Лw�dF�W U�DLZ7S�g����N�M�a�$QS���T�辐�>���q�����r�u�������Zm�ˣ �a��L:m[������&PW��6�,<8O�ÜԔʾN�gO�6 ��׿*�������T��CM~����f�ڎ3p�L��5h.����Ad@����ѿ�VlԜ8�F�c��bͿ�I�Oٲt"�r1��;����}'�����׷[��,y�VRe��?�vS���V�g���M�a�ַnz\,p�@ B���ϴ1+��gT��",���HfVʓ��LNCӫ1�95�oJ�Z�����]F�s�7m�ݳ�4I���pQs<s���$�?��� ��Y���2՝�S�Y� I~N��;���6/���T7�t>P������Gο�Ƚ�d�$ۣ�x��2Ѳ2��~�x.&X�=|
K	*��W")߿Y� ���c��?=�U��� �:��A��0�X��2�`5N��*���}����!E�n����؆��gU7ב��}�����f�oX����5KAЋ���Q+ю?V�N�JO��
Vk���<pT�L�%A)�,������?:�;.`�Xl�9W]c�+�y����xo�>�w�e�{"��6,^��ר�"�&�A�z��J-6i�jq7��Z�Z�3Z��n�����_�>k7_HOt�J1ӕ��bn=���32s�P|��3�������� d�{�ם������{��'�5���mC�[xO$��%o ��9���<�hI���P'd����Y�ҋ�-c���T���Ķ\q����[�a�2�{Y�З�֔;�����p����S�hS5ѱ�BJXWU:3T��`���=��;/�}�<y�y�V<[
%`���ƃ��~�_����������h�L���~�(\��¬��6P��v1�cY���E*���q� �Q��Is�+�D�R����]��P���<��}ޝ'���?i%|�c���Ӊo���o+�e'�xi�|X�I�)W�A�b����&�����5s���{�V�Cm�L@�B�����������>����6\Ͽ�N�Z��R���)�Z
7F��Z	�ǻ��oV'���
��bc^1&t+o�:�6�O78Ǧ�R�s��g#�A=�I����ۆز��Z݋�r���e���AJyA<x�ɈF-y�:�A���(�A�`{��ĦF�r/l�~v�ӝG\) ���e�:�ip�>%��?�#6���H�lo��
�?x:���2"ƷT�LY�Ǥsݐ	ɦ����1�|�|S`d̟��抖ґq��8�������Jo?/��[�������^_�+DL�""$|�*��	`W`x�)>e ���DE��w����v�T}���Գ!šdB]�J,ި63}�O�z�����t��U��;��7�)���;��^�;�U:��i;|���Ms�A�ϙ��N�Ϝ�}�ܹ�]�$̲z�3m/�<��2��W��r���wd�{Έ"]D�/��N��W��E}�*��=���[h]���C3�T�<�.S�Mi?Z��u��څ�^���lU��HF��[��O��-�4d��K�}yY.>�K�qf��~�Q��(	�y����E;.�����M����#HU���tڡ�N�z�۱;*�L1@%�� �D�I�I&aT#���>-�JC�;.UsK�<��c8.�%|8.��H���C�&y���N��4�;H�@�ʀe��z��Z)�
��?�}ʐ��HE΁�74F��%o5_4a���'R�CG}[�"��d|��#�,�pj�v���z��w��So]�H�(ȿ�c��ɹ�}!�nH�*�|e�I��?M����P+�8�Qd�P��ȶF��eK�������Rb;���i���p�~���l�.z�"ZY���r0�m�p�?�^y�l���&�/�(�:��.�ƞ�/��-9ပ�j�w�Y)y�Ԡ.�1��Z8�|�Š�ݾԢ,��8h���f�'��b�K=mdk�RS���Go���v]��Wqj���#���T��?����.�	,�
��Y����_�7�7^� �7�>�(�k��^G"sԄ`J�*��?�/H�S}����� �  q\��(j����1_��}v�H��<�Mt>/F�'^<�E.9E�w�C�l�Z��>̂i39$�,ɂ
K���L ٜ8Ǫ���&��Bv@[T���4��@2�g��z@�X���ܥ+:��@����."�2�]:�o)��ͨ��F���igE+�.��s�Qs"Sڡ,�iKw�L;%r��,���M��њ�^x�ܽ���7���2�t��\94 �%�A�dx
���;��E�A$w���� �;BOd�w���:�7Y���M��%Hˏ)���o<�G�@u��A�P�˒O�c��g���0��9G���W���9�ʿb��\7�M��,�w<|C2C"C����T���E���sL�+��RE���w��K����i���O�j;�F�w�p$q�|�����z��a��Um<�4c|�ɖ�b��b��%!**ʶ�F�A�IZFf�#��%�|�ͣB��IJ��7g�h��Yu����	����GohF{4��~�.���[];�6:�zq��������HbC3˂�G��T�ӳCS� T$�&����dhD���rQ�R�
�s���?���������"y갮�  �	�KV�&4w/�Y�=ވ�p�_��m �v�sF�?V�kﻸ�g1��x_�u=M8םT�_�<�gy��j�]�['��͊�m��:��9,Մ�|<��t�3�I�^���Uy��Ero�m��ʲkN�c�C�&-	s@G��&Ǜ|J��{xc�{��!H��t7�^$�@C��]�$��V_��s�>��>���[Z���G��%�,�u�%�r������F_wg��-�A���x���]�D�Q��ћƇtC<�W哾GS&�<�D�K;�A��e���}Z
�:��uS�}ލE�}Y��y�kЩ�lK�p�	ǰ'���{��e� ު9���}��1Q����䃫��;-�4&���=���U������=��w1�I<�9ݎ�Ӯ��,�Q�z�� �EC7����>ԃ�� a�lw�꠷��ϱ�^.	�8��`J�.dM쥚ıE,v�{t�d_|��}m<y�6�w����	n&��2I�N璏��+��S��'R���ҕ��p���@�>��RƖwt��c�+b�E��w�0�w�CUu���� ��3!ŀG�"ԍ� O؉�/��Lҍ"$���~c�%�r$O JĢ1�с��ߖ� ���c��.�M�Ͷm? LR;��̜��Գw[2�;�rߏT�%A	$o�2JB�<��]�������]gF�L
T�y,�U��7���1�����ItcS�h��V�6��6�{h��.��Hj��؏B�F��F{����!�E��������g�&;�$��~k'�w�&r4ْ�!��]*AϳY�˯�^�}���c��o���M�W��"
�!�)u� �(_�[�O�k����=��[�	��F؈n���å?H����� ���H����o��n�+�+����q���\�|{�d�鰲�����B۟��<�<�H}o��V��˨��+w��i�=��E,�J��U��i$#M��ꏜP#h�g#@��#y��}.-Fm�g
|3q�+W{�����tP�B��w-h=����va=_�e�>-E�wZ[B�c\��yt�����Y����`�4�4��^��bs�'��?�q�Q�v_г�j[�{{�"ei�
��#(	91�Z�|�y���~�>Ѹ8^�����6	����O�_���q�$�7)P'�}��$�	*w�ԕ+���N�,"�?�j��f�<G�#�\.&���k{98�u�_�h^��v)(x3�$D�Ļ�������22�l����˔0�`�z7i!>�*��ffZ�f��I6�v�+)�7)� ��,��zٷl/�r����W,��yr������^�ʀ��1u�����N��w���|�������Ԟ�DB��|a3����i�?�Z%A���l�%i��x�,
D�1�Am�Q���٢%�0���s��t'�m�Cn�#���j0�<-�w3�e$X� �h�&�^[���M �e	z��!D'�sܰ���݋_�0,Sn(|�hf C��d� @3�q�w?͜�z��i�Xx�?-|�Q4���te��]�ʗ�כ���3e[O􄈪Ҹ�����X��U���8��0�汣�\aQ����6�k���@�5��L���'���H���'�d&�����&�6]Dx�X8�ק�2mH�����8�/��4$­y�2~g�+�Zx1pP��5����ԎP�Ü�)�V�Ͽ����O�%�7�$_%���(<$���5�r^wi�>��u���Y�"ݏ.�i�f�э���z�y�����!1�0{&��N��5O�lנ��S.���,e�������)��ª�w���=��ۋ��0��lى3�Η��ͥ�m��S.��B�ȏM�R�s���uC1�ǊK��M+x�d�N�{���I@^P�?��V�uز$)?�OF��%m�ݙ6Dp4���X'?��ʺj �����#����,�9�Ѥ++>��ܽ���m�#���e�+a��&��s5�_ڻ�߫`��6�m�K���gN5�g9c->�p+�����:m=����@d�gk�m����W����V����3�HV��t�IWh=���� "��ѷ�q'Q�إ95J[r���9�j��F�@�d��vs���|6��|�,)�N�g�HO�E�(�Tu��$�sX���fVX��Ɵ��5⒐���Rx��W8�y���_9�����c	�c�����	$��m'UG�R��e����{��͢�r"���cN��<�}�Q���ƿ�;��^�r?���Μ�ȫ

@���C�~�Q*��QQ���)WWW[���6��Þ�8v��F�����E�	�	zm(�I���\�9�|X~wK0��u���Q��x\�i(�VlF�=-����j���E�U;����W��a����R�rF`Ʊ�!8UZ*�=�3�~!"� ���x0Ji��I�z� '.�k���.��������㙥�e�[I�l���b��m���d�>G�Z��ƍ,���5����/����A��_,0$8����4�{�z@��~���q)�u�X}���ܱ�U��z�M���]��K#�$�l��~���} K�� �F���87-�n�S�.x�l��Yb��y|�B%��~�3�����U]#��*�8)�R�}L=>l�+���bA�>�B�Zs���
� ��r+�Uߥ�¦���5l-I���]�Biƴ� mOcF�����>��Y
.�f���vM���^�@keB�`S�1x��5�I��5Ք�(Hۢ���|(�/���}a�ݶ���� ��9PW�?�<�dq�m��#St��1{uq�֕�.�y)-;ƴ] ���������֏��ڭ�`�G]��������F�.�Vì���0D������:�t��o̝�3��d���o}"�����Bs�����X۝��P�D��BX�'��{3��Rz�3쫶�ο�ܛg{nO
\8�7�^�����q�E���� K�4ĊS�B���by]�Dg�c�_ߟ%yIR��`S��l[�3D�. 	���~j�\j��N�+v-��h|L�L,w[#��9��"��������2�����v��Z�;��-cKj�l� �,azu���\��/P��p#�#��D���C�E5E�i|��P�}�����p�,.Ҷ)�b�)�{��Q]����G��
�-�����#_he�iY��=f�0� EJ��~t�BZ��~̑i���VrR��&2��z�Qf�2|�<3Ǹ��+y7լ�`$�-V3�Jj�E&��'��-��_����幾̬��s����<�Q�7�!�4��%�?���0?|��{����VW*�.p^<�뾟5���{Q�6_���Ս�}%�@��卧�,{��>��hx


 <�C��B�����G����+A�����i֟6Z�`5��;�1!�ZT�P ]��Kx��z���0��q��K�ϑ��4��<GLX�9�c�"��ڂA�ӵ�?��I��r^}ZCn6+��?`ô�W����y��,�?� 4D��M�<����~�`��A���jd'*Z�e�ѩZ*&�SE>-�"��Q!����?"��������r�ܽ��wn�4CeCX���B �t�ujuWL^֭�
ۂ�T������a��V�A�BZ2/l{��3�0*�g��-ݡywTɧ}]�|n�I��������GÐ�
�aH}#'����˨����j�NÒ�{�¢ ��Q*�m�hG*�e���b1��������Ǯ,�%\�7e�:N`��.(7y�S����������h�������m��Sk����!"/ON�{�M��r�׬�?>/vOfn�Z�o|�u]lՍ1S.�o-~��˗�IKK���j��]�R,f�^��L��O�vW��f��S�{�,�d��<_��XJ>qQ�ȶ@�UB<z��� �<<'J�U�}�r*�{��pD���߁>��4۱�����T#o2�l�%Im���7O��Uc?��+I��~dݵ��!��,�@�EC/��r�2:�;ˡ����b�$�{�V
��},��D�%�//�Z4��^ÅK��7���`�δ|��[��R{ ��=`M�{1*H�~Z9�������¥�]�*_`P.���gvV��C��7b�RC�3�F=,���.�h���k�!^8z�����<\�����}����-��U�:�R߽a"�������0(���OZ���;ȗ���/#�>^�y�/�d&��$-�*�dM*�"���x�(5�O��(��_�A��c���QO��;T��|#,_��C�RGJb��<=@��N.t'�!�F�J/�G�烒����)�©�ޒ�<t��З�T��ǆ(�u�����������q�b�<\IQ�����>#�L4GW���ZjhW�D ,�g{��L�ymL�_���q�y�`&o��f0�@�˟�jR�=������PY#�	��N�x_��鵹���I�(�������Ϣ-�!���&����T*��?���9�p++���������E�� "��fmA
n���h�{(=���0��Õ۱d��f��&A���Z*�_�ק�*�y��5��:HOc�Ԥ�n����1�����uT��r�!�V
��7:AwY�O�j�Ĳj��O�u����a�0�y�7�"����Y�&�P_jl�����ت����@u���[���c���g���\]��<|�X�p�/2��d������ᥐ��to���FQ�z9��VY9�]�/+x�Q�67y�O'(�G��(�t�^�i���H�F��a��	��E;Q-K�����!�ev��A�L¯�t��6�Z<�����K��Ȗ�ǲ[�е.�b򲲨�(�<�;#GS�3a�޶3�0��8맒b���W4A�4�A�Ww��{�,~x���X�+=��=b�7�ĳֿ���i:�DcK����j5(���-���3N���c�,JξР7��ee�=L.�AD��=�4�	cn_�J��A/#�V>m���9$Y��)��|��:Q)Fj肴.�����hT#EY�]SR����T���mW�]����~�;�~��ۗ��#���@jQ��^LΤ��7ޏ�w@�^!k�8��s�I�eB�+F�8c${	90�+��.���qUR��?���k�D���e5wl��|D�#v�]
{��y�ub6�/Ը6'^��lc��E��4��G��������1:Yp�ec9�U	J�0�I`��>Ϙ�3�)����L���ބ��m�/��������0�z���@�k�i�vc�>����-�Q�ط �-�EI�������)�c
���lm�d���#������s!-�~%���OV�Uy�u~bB��or�܉OQ�[�=��p����O���qh
�,}�IwN�SW��ɢ9h��fr'�ٟ���K�A���*��#.:?���T��|w6�����:���8��,<�}nYҝGq¹�Z�5j�뽂F^1$O�qo��k�i}�g�F������Z��!�M�x1c\Ք�C�c�`�G���a|�qԽ-��z��è��Ů�;:t|s˒D⢣�o��,������[�|5,��j�~Av�GE[�+��*2t�Q^x~�,������[A;�a���%�$]D���*���|78��tuXޫ^�eB�H���NeP��6\?..��7bm���U�s�� �[ ���X���7���W�B!�'X,�;�v�
��'����$�)���=f}:�l���f$o�+�D0Դ�Й��Q�E�� ���s����ÿ�Ax���uT�bhW'y
֟��ii�=����<`[J�;�l݉hy�_��+��;��|PZ	�;���Hy��v��.�wj�h� ��q�	'UE�ݯ�
�Pahǌ��
��QLnS�@ȟaD�ն���Q��]��_�(peX�1s�$f������r������%$f'�;ժ�B+��Fk'P�*�M���x�S��?��!va����q�����f�܃��:�U��q�VM�XCn�"�"(cW6�;����K��ر:ɘ�"҂��!Kب/��ֹAX��cƞ�p�ݟ�Аe�ŴGZ��N-
���\��GĹ�o����E9ꭿ;�h�����*hR�z{dy��#bg�y���}�����e?+�(^�+�n�nҝ�	R[�Cv7H+o8����y���ْ��@&,&;����/}?��.YV�=��X\�d���^���w}}
G4��^]k��i,���#wU%d�4Y5�a���4���F�;�<�B��5���l"�**K07�m:�n�J�h�tv:'��UA�O�ql����H�F:nAed�A�Y\���B �t�f�o�D��V���,˽Q�ޖh?0�
tp,DD�/!��w�����*T��'����uRc�����yON�z�4��s;�ff=]��UJ��t@��x����gʸ����G�'
����S���-�b��2���<��"h�qȵI�F�z{��P2T�*����D@����w�Z��X�K��T=ʛ�63�T��Fs;�Y�(]qT�$�����ËZ�e�(X�^4:���� :sK����y�ň�I�J!�[%d.C��5I	>�N�y�OMQ�B��:{S�~��S��kB�g�P���K�JT�v@I�ʬ��`zX���~\��_��x������=~�B��3���)�Tf0�Q�@�mi4EFK�~�P|<�=O�_��?{m\��xeao��删�\L�C�,ٓ���94���9�����7F=˭��җ!�bx��~աY��H��i����\�l���^�)�P�*��5��UD�p��� Y��V�c+5f�w�W�rq��uۂ�#S/��%��j���V^R� |5���DU�K���~����.ȝ��5��v�!x0���c�Շ�\E�.�(Z��P�c��d� �s�wn~������:��X���]��*�D"�!s�K໛�u`��(BV�Pb$�;ߜ�f���g���j N`���w��ۂO*�9�A��B��s�
���]�¦C��J�C�<H�m-)[���6�	� ���I���6�̛I4�N �
��	���0��$���6�M�RLSi�}�^��^9X桥,����\���)�L�{��6M�`3���6t�u��H�#ٟ��׷_xFR�|���0��F�)x������"0�vG�����h_���.{�д�y�-�r���o�_��v4|+�#ߎ�l�O�pz&�n���n�X�U�쑞�N�/��=|�
��-�$n�?�7Sn���|����%�Ų������8B8��\C��gӼB��3�I�ʕ��l��s�9��RJ)�V4�0��%���7!�'�E�q{, �IJ:dX��7���!�z�^��ϛ����%G���@U�]���<v+&�'�j�F�cH�c�N�c���9`gϥ���࣏J�p�(�d����b>�u�`#��Q���ۈO��hL�XQ����zo"tF`�9�l��di�L��f�+�M"i������#��;���]��|�=Ʋ5V���H��V�k�OD$~*� -ӯ���q��1��5c-%�f�LM�t�C0��O���R�e�t��z���]�/m� ��\gC*�{�H�Fm>=�f'�]Q�~�ڄ0:*w���.\4_�#)�P^�<��*%I�י����c�����^�5��+��XKJ�YĬ����FI#Ʀ�TF|$G�b\�`L��B���o^9��f���r�}��F�`���嗕`�t��+��z�A��8FӐ$��+�&@�kk��@�0`W�{PF(A���g�D�i�ӹ]D�{�+x�3�g]Le��J�q����o}�TE |C��_����WP��J���U��Jo�����k?B��0�z�`J����w_���MΛ ��n���f_�����Mq�'o��i�j��C�u���G-�ea�`��5���R~~њ*�����@�e��`����]����  �y<8��N�c��f<
`��z\[g�7�ۏ�u��v��`)d��U�`b���f~�i�iuqg��ۀ��W�%n#�K\�m�$6���6l�p*0���c�R�7��
*�T5�@n�q��M�;5�`��������nRܼ�9���E_d��n��y�� �=P�A�?}���7�|�Q�H;RIFp�̝֞�t	�=]��_	�H	��@9���xU�9�yQ�ϲ�Ds[L,���̷��0C��!��bF��"ח���i�����Q�)����TueAYIj�=�[��փ���<\
w���-� w�I�8�w����Ӹ-�\�1	>�����
�����G��k�|��u]���߳kK�I�ٔ$;�-�_��$�����گ���o����Mm��fA�����|7�nz?hH�)��_�d�&]�����-�x�j��`,�\3W��R۱��0Ia'�/�'�祉_GyjF��L�g��(2xeo<�]���b�a������}�b���6AA?xēxY�=h�����(~�b�h7��>@������w�%\��*.��Nx��lΊ%����}��/���.���/��7��4u%k����x�ϯ{G��1yk���tn��.J���n�s��W0��.�v^��8��s�w�=�%5m���KY��>��N<�������(�L� 7�C� �0�d��{ck��#����J*�뿾�;��^ �X�I>����?G�r��M���4|�Q{\��>�3�� ��o��ϟz��mG���)>�Y|�+_���� #1�)��=���b��!R�-=#α�,h�H0��_���׿�կy)�Zb�D�ԍ1����Z#Xg��2�h��}o������W���O|����@�VT݆q��C�T�� b�<�:Q�kr�T
�p��=�o��Y�7��L^��cxp�j&�"�]L��X2j�n��qo|��~��N�9n�>8k��?�z���>��~�k��匙6��)(9Lty�1���{��N�! &(�Ɓ��<:������g������.fͺ1��#��V�F��y�GE��V��f�~�Q�p���m��p��r�t䗿�1�{���13�Sl������ +`H��L�5��W'�6�1S��*�5|�_`����<��?����C� c@�TZV�.J���$�_GWr&�.ζ)�	�f��+�͵ky��wCx�4c����?��4o�T�e�\ᣟ�4_�������g#۠��S����ԅ�
-�>�yD8��\}��T��|AM:�%���`�kb��l�T�ip"�OI�$�G�X���}���	��Pc������u�"f�ݕRE0���?��狟�4�x�����������q'2�bw6>8�������;�0��㟡:E��9N��or�[��s��,�%t���`"A�8�F������)$듸�g�8�pMl�������Ag�u�*z��/���¯o��y�S��W!f��?l��3�I$-���A�������uw��B��":���������^���"{��.p��?��&78Sb�r����1?�f�^m�	b,����G�����߿�ʻ<����������������FG3�D�u���Ҧ�<qF�C��(���J 
�1�-b"�)2�[K$͠�j�����;�������G����v�:��v�o�f��kB��G����5!2�1`�����A�� �,��"�=F[7��|#���0���_[���8�q�>�����+F(=����9�e���0�t��g\�����Ye���в)E�%�M�h��iYKwb#���?��/~����X�c�w�5������W��H{Zzr,��_���o��sϿ���(%��l_��G��;�݈7Bpӂh�(�7���q�new��'kԶШ��#3���0�pk��`�>b����3$�P�1�&T�!���������9AE	��&���4u�nb,�$~��^j,j2��h5��V�*7���[��	�Wj�73��T@Ӫ��q�5�q�W�c~��=��Dt������g���g:��7]�-�U 4�>�y�b���{���$���a5�l�����v�5v6BY�(�^��gu�(��4�B��2~���p�3�dqf�t:�6Q:�q�����$ 6E��ԋ\�Qi勉�Q�HB5�t8Zl[ĥ�h-�8ڹPt#bs�py��[�`�<�rF�f�{��9��#v��ifc_i�f H��?���������笟�/"|��?�i��6�H����hc@#�ا���~�Ē i�`$e1�&�z�X���-o{���/�#���o}�w��[��ǜ��s�4��	o{�1��`)0�bP;�Z�$��nb�Rh��������GD�`��[z��̴�@4��2*�KƎP�a�9�E���#�/*y%�>w���j�h<^#�Z����Q����Zt'��4V;��q|�8������!��G�U�������9��H�]"%#��O��o~��o��GB���6z�F0��,������-�]ˢ ��Pzlf1���l�F klt��jQ��	���@0�GL��Y���uc%b[D$�`�rb����4jӁ냇�#�j�"������O��ř1��]��jzHRf�W��n���7bB�S��������iIZ�s.+��n���}]Ăs�r���F���T�Q��Q�����Do0�,����/|c8lF�g,�^���'E�AT�"��(�}Ǜ��A��O1�;��.b���ab������O:�']���N�$_:��8I7�X�Z4�D�ox��?�hl(�YFA�9���"FMD�K�I!�i�G�%y�P��Hc�l�����b���u��;T��,��(2���و3 Q�D��ډF�{T�y�Eh�C��`���2^�2����$Ni2��A�c@��K� �Ӏ��ki��f���^8�P���Z�)�����}�%�gz]HU��nґ��^��j�K�XKZ�6�,�1��eQbmF������Ŕ���C��.=����#t}hfXKEc��QE���[t:b�Xڣ��U�LU)��̵�1}~���=N)-�d|�[����\e�KKBA�H�]�ig�K���~�똑%���J���/���g��٘��H���/;�-G�Kb�A��GF�W�ܦz���O��P��1����HԈ����4n�V��m��F�6E�d���8�Y�2�u��a5�`L�_]`�q�X7��΀;K�%W���b|#�I�d�fIM%V�Etx����
D�6��ۋ.'�������<�1�En��V���F��ȹ�N�ǾL�8ǚ�����2�8ŝ�@�-�x��F�������G<"ڣ�5M�N���.-�j>�1V�D�^!���U�"���-�:CZ�@+e�VW�lu[�;�{E�)[Q�[�0V(��u�1͂.|oӚ���L��]�	ZAQ��v����-=H
�)5"�H��ڬ5 yDឪ�YKTm�zGz�~�cL�Ӎ1�V�N�ҷ?�-0�`K��5��BUi�j�2�T�瑚�F�Ĝ(`D� ЍZEW�Pt6��2+��&�5���1X�\L�����h�����t�H�a����E�K;�6Hŭ,���4I�,����HBH��`#��"�1^?|�۽Ȁ�ר���?�I�Cs4=J��x��,X�M�����t+W��%lL@�i�:D13���F^G��S�B{xA�;#h4b��(\}�-�p��՞�����G�ʤ�D�4�j�0��0QijH�>�I�X�������dD�y�W�*�I4)���o�(Ƣ&V���j���T�{�S�Mȿ�.�?6�;�eD�3��mL�*��e�$bo��Nu��
�����w͍1�3T�!U���	1mR�!(	i�-�4i+T���H��P�wdڝ�8�Sv u�=n$�a̗4i2[\��4��Q�W���uH���:��ʔ�ȌkQ�4	R��k�l 7�|�IA�h$�����*[hf �B��-Qs���S��橴m�؛��ؔ��*����ED{@+)Ud`L�,w���W�V��BT��Sh#�HY��d	}��5��Q�(��eC�A�7�ª�@)U�00��2 @��鋋�)�_�xn]��1���&#m��c ƈW@�$��x^�M`33@W}�� �i��S}C�\�'���N�}�I���a�����Iq�XѴ(�pzI��*:� Gu)�S� �JY��h̔}[s�6���TZ?n@5���&z�=B���1Ev�xB�r.>j@h-���u$3���i�Y�\,H�K�? ���ncj�[�D0��#2��6�?k����j�,Nr$IǟLƪ�%����+�°ax��}�ͤ.��"p��n�V��A�
��
6���k��o
���a`�c,�p�?�G�E�鴫�.�N�4(�1��OV'1�mQ�U�Y��w-i���;��c�ك'?�1,a�;�xѢf��/K�QY}�z��� ��r;��yw�qW:���uf��R����@�3K+wdVpΠ��z%�3��<���S�Ò��K F�h�NP6J�uD`0{ƫE�=G�	�O}.M	�J���F�?-��u�?Z4��l� ����i��d�����<Q0�,5��v� ���L>�j_�?�	��>�U�Rc�ͣ��p[ �*�W������ފ����ž��ǚ ��+�3t�m��Ԭ)6CS��(��a�Ddz�+�I��L���dn��"�ku ����Uw�h�I[<��<�Y�`��w�1{�h��h F%�����2��ha�=w_��/����υW\Ņ�]ƚ���q�h��k汛�R��)��n�ٞG$#�w�n��JL(�֦Ȗ��oz#�d��g=�z�b��s"��;��5(�mq���?�<81�h�35k�hl�>�F#�ae��0���ƙuF�Ĺ7U�ź�S�n�����YJ%��a�~;��nOFizdFg�?s��ko�M��P�&���jm�d���o3O;T��AGqv0j�4��޷f��v)obJś�R{�z(1չfX�4�)=����Bm����!��	Y8H������+)F�v'�˂\<�F/8�9<��Ϡ-����D4��5M��Ʀ�V���$�&���}�^y�sy���/ug��<ƺ%F\�p�l���KL�4��������R��~�>��F2-�cA� ���^m�P6�Y�i��Ɇ'�������靖�x��}�����Xi�;�35���V��ͳp������ ]Ƚ���i&��f���>�@tv(�g�H��v Xkȍ��C;<�Ч���a�;#�j���MIlJB#UʐHP<V!��%���>��?�`~~ι�y�ŔⰥk��^3��onSu�S��G�6w_�0���<��hm�bW X��3����A�Ap85�)LT������gDu�S�|���?GL������5g����
 jۢ}��6���K]z�p?>|@t�UF�>z�����R���cx�>+mB1Ѹ�M&�s��,)���,'�2�<�9�h�505+�H;ˉej�Y"�W��<�)O�k����y����%�6T�#C 1��eKi��%�h���Wq�%S#纉�֜��W�H_�&�8%��'=�O#���Ho�����ɾ���+?f���ew5��
��q�{���$:��_�ټb@KFZ��vZ�;��v\2���A�4�7�m����+y���>�쓔���7�|+�\wkﻗ|�Ͳ�K�'��%�ZB���N��7p�w��-w�K,qݭ\#�C�P�k����3"!�swRϟ����&�~��Kl�m"����YbP4D�5):�_ꥳ�ފ@#X���u�	*�y��'���P�;�Z�d�iN!�h��������1�dXx���n�|���t(��I�.-9�)O�/{1�G���&k���.1D�_{?+w[ɱ�K����g��d�PY�����v�>�Wl�� K�VSB���v�a1��7���~�%���,���C�P��(�T�~1��g�>{����Lu���d!Z��g���xɦ��������u8Rɖ��(�l�lU1V]w=�]s��Ibq��%6�11���q�a���َ!�%���U���n������	�������f40�v<�����W���,b�c||�L����TM��)/� 6������� c-GqX�O~�36���n�8눾C[,NZ���攠�ŵ3*�^��#{�)�6g��g8��i&�l��J���4C�D�� AoDv���'7��v�<�)�H��tS�q�L��"�����4]��^����3o|�*��@f��̪�/����/���?4\q�5@�����̣���&b}��+w�Ǽ�Q��9�� _p�&cbb#�^{5"ټ�We��L�o\�Ո�Q�u�L�4�a_gv����K��tKvZ��7��e,i����Ⱥu�8�cY�l	DcL�c Ɣ�xT��(*0��#pċ�`�����=��w�!�`7J��d��W��{���-�@��<[�ʛ�z�(������l��H�q�0�C�>��-�evC<�.g|�}E����c�NG��HL[��PX���l��B2�w<���5��'<�;F��@r��6��i^�`���k,�e���1l�ek|E��t03j����X&Oc�}=)�ؠ�p~�F�ܑ9�eY(��� �Q��vm�+mg��G%��N�&b��54%�|�X��R��o��ic��V�#B"S�M+s�������� �B�e�9u�Ƚ�]�F�d ėc��u�"N���X�(& �k06�[��_�ZZ��Z�䮎TRqӃ!cf�$@n-��E���?����6˗,�SؼEP�Ro}�+�����'(�`,>V��tk�6��/3D	�UbL�P���Q��]��i��Uk'i�R�XM/���Z�li?o_���"�vb=�#��8��d�Mӻ��C
�����2�Sڃ�A��2�D���E�+H>x$���XO]����,i筴߂�C�#��.ak&�o�Y���#J�,�(1��F8֑�X�YG��YNt9�:�Fz�-]��{=����i��,C-bE��ZEK�%sm��f8����x���Ґ�ϭ%xLT�i�.hڛ���)���Y�i�ή��M�{pb)����Pr I �ZKJĥ��m��#���G>s��������p��k���)��x�"DuX���x2S��׽�;L�b�,�:��y�k_���ܖ�Q}UO��k~����'ج�F��qN�c�%���𱓿���m��Z��]���XZb�!Q�Dk+n��!�(�M� bQ�q�@}Ct��E?"�#�W����7��b�a�CU(��,�(���
��4��s:����,^ �HSսF��$�Z�."٬�jg�b����`Mc �c�L�֙%�i"G1y9ؠ��8m�m��@�EG!D�:��a�����Q{m��,ʖ����:��>o�k���Y�ؔ ���lBD���Pƈh�e�i�����"T5����*�hZ[`�)}~�ƿ�@Ylk-^�	כ�.|~4Kљ42��b�AO؏'�mGe���xg�W���,��5����=��䨣��[��˖-�:G�c��ww�~Г9�ҫ�xC&����aC{5~����g�H�h��d�v�G��2�|��&�����0����	e��l�6tp�ͣ[��\�@'b����R\eI�BKKG[�l1����F01���k��X3��L��]�-j������^�`�'J�{`��#(!�Q,A �,Y!��X��D'�E�X�恁����%3ۊ��B1��+w!71��m"��R��V�Am��ŀ־ms{��A��J���m@�DJ�ŶrBP.����? �HY�XW������ /C�#�;V�"β��>x��r.��*@ȬM�gt��$��ƈS�ˏ|Əc��S��s��n����1�dh�A䡁}�TsZ����}���o��N;#b1��1^r��蚛��m��*&F���icg�5)���7º��bQB8#D
�Z4��m}��T>DE�F�Ƒ-]���`�K��Q�e�}v瘣^@�x�z��j�p��wp�92�13��6@45	v��ig�'?�q�C�h]�ݥ���%���E�2�=.o#��F,���Pb5��N;�WC�ED�3x��r7���dՔ�	��(�I�jO{t1�{�[��j_\U�q��/����&�.!����P� Zu�G�$)�> 
X+�@_u-�^qՌa��z*M:aE=/� Y�Sj^�ȫ�������=�B�*�r{�#�(�v+��u����1�4�:�ת�I��ۜ������sX�d	eY�g���/�ه�/λ�R�4lS[�u�����ɳ��(�p�2G�4�4*A=�Q�J�nG��ĩ:! �st�"�.�DQԵ�cb��E2�et�%�F)���頞i�k�,�K0c-Đ��V�4C)��.�]5���������\"�XE~����)�����M?;Ucq��Hiz�UD4�!�X"v��P�
/DA$6�6��<b4��״�@��PE@T�J*(���l��&-�9���m�v��L �jF������R�4o����yɑ/@b�H�_�a�=w'F���È�v�aG��6�n7���H�gp�E����o��N�h������'�	#P�h��?����JE�ȳ�=���1u�]PL6�/~s�8��ܶ�&�=Wݠ��q�5
&4��)�/H��u���K����+�a�s䴢�	T�o����L���Z�ԯU�k\	vͿ�#2���Wb0����y���j�����q([A�dKD�#C�m�>�z����&"�����0s�׹x�t���C#��8T���nU���>�ŋZhY �R��x��/?6|�ƴ�h��5�:�(���t��Ć 첬�Ӟ�XμtArl����T�������y�cvG|AK,������G�e����`��/9��wݭ��>�K�/����&R��6,��>Qi��g�����R�965ϩQ!���j��c�R� Ʀft����
%μ����Ť�`z���o�+�9����'�3�kf�a�R*c]��}�P�2��<|��$C0y�����u��Oӕ��X<J<��돁�
?�H͘7U���6�X(+�
}x�T�2�,'�3�
e����<��'�� �V���g:�@=�c��,t��B�,����r�6%y,h�%�:P�����g�u'�nV�g��YG�ff����b�Fl�"��L;�z��M��]� ���[����4q�Y^=]��볯�f���ۮ!�������͋[��x������Q�D�4��Կ[��kx�7!Hc H���p([�j4U��i@��3j�"�ؿx���"�h�i_3�}���@T#N1&�QH�F��H&��ǒ���!h��{��ٍ���&t�/HwL�/�+/x�����H��N��Y�jaC�b��� ���<Ř�&�dĨMbR��Iׄ�s��0&�Q���W�2Oc4� l��Ue �f ��ջW1u��T�9����T���^�V?UƦ�fj(�|�kd�sDAR�~7�K�i>#�� I~�%!�UyL9	Lƾ�7��V��!D�,��1c$�i�j�!u�׀a��
} �~�s��}ॲ�[LOZC��˙��q�纹��eE�C��d4�0��{R�'��� U�`.괡lA �t�M�9��Hy(۪�*+w����f��5kY�Ê���,P�a���_��oL]J���N����*�W��l����D�`�v��7{�nm{<�)}�~����[Z�Ňy�ϪDf�"��c���ʑ0U����.�3�d.�e��,�F�8�u�$EQ��D�_���&F�}u6�	���Þ�mA/go��OV��䟩eu��e�Ǜ��t�f�[�:��ߣ��X��.�ѹzP�#�	���ΐ�k{G�}ਪY�w�}0�2�!b��2G��/4>|u��*�Y�xє�?f��4���6M[4t��������'�2|����H_}z%�*�:qf.�V+X�����!����E��J��ED��|��鲌Ҩ�#!B_�ғ��'�lk{CI�q�U�UD��i��̰��N��ʡ��*�g6/�Z��`����I�V��k�s�*�Du�k��M�?����e�]vi�b�9�{�р�G��! VX�r7\�n��w�e� �b�HߕW^����*R#�`��ex	�b-X����%�\B
������ ��:�˯��<�5���or¢�)���
ZL4�Y�j��\,����LL��長������@�n�9)�.&�WG�&�k��ۢ�M7��y��;䱿YQ�w�)0�
��"���Ӕ�Å����(�FY�5n�X��_��eY��瞍�zD#�����1��/�E0F0bX�|9��V��w��C��!��Y��x!l�w�k��S���)5i�T�kD0ƥ�b �f(s�S��Ny�����bȳ6Ƙ^��ƘfmoJ�^k ��i�u��e�6>����q��CT�SR�ޛz�C�~z��w�'�fkl�����>���_j�;�#������
>*�r����A0-�~c0xr��fС,�No����VŹԀd�`+K�%}d� ��*��.]:5d]s�ie�cEQT�B�CQX�v��F��BӴ�š޶2��q�3�u�x�p\�P6q�Ħe�����dt�Emj�����	��gF�Qr�k1��]���T�Q�O���J�kR}s{t	����^/ |Q���Zd�U�#�:����x#�Y�������D�w|���9+c��jU���+,Y�h�;�%�����>��6b����֬����2G��v������R�*�5F�}p!P��C8[��呖���l�`�&G����s�iDj��JQ1F�����{1�NE���2��	Ƃ�Y�	�qW����Lж�P�����ԙ�������F��P�i�	\χo�L0��P��;i0��:�A+���2"��`�{��5��P ���LC/S��b{ �Qif��.�b�&58 ���m��5l��c�[�1�*ݹ���ӓ�h��B��� x2���Xk)˒�ѕ��O�Y
�U�򆛹o�$ƪ�>*Ѷ�x�us �8���̏��#��mP��[��|�g<�@��wCy�Ѵ~D{z�،�}�T$���Y���_����L���M�Ძ�����<�h�%~�5FM���E����63�jN�������W_s���Lf��5Д��{�2����-����vuJ�V�uUP���A��!�^ ��ƍ�wY��t������>��ySl�WރLkTS=�5Jwb�H��s?*9M�S�,1����t��O��j%��SOC���� �������̍������c�����*j���R"S�2oNAu ��m ��Ŕ�{dk����ch�Z� ��m�X���xA\�-�mH�>���WM
��E����ؘ��*�ZH���\���<��7Ĩe�n��K;�u����;7�ޘb�yҌn����,�.Y�=C�,���*�m�lk/��ըk1`������5�Z�\6u�3 '��D�x$�ʏ�I����g`Q�Mހ9i@hĩG��
(J�'Ԧ��!�����Y����@h��wB�F�,q�3HP?����4U�<"�(P�p7�v7��AG�x�p�*�4�F}���v���y���v'���mSM��m��$�2>>N��e�/jt��n5u������^=���ׯo@\��?�1���٬	4���7=�m�W_��|��3Xwf�ݝ�v��}Hؘ�����Ĩ�L�Cr(�R��ZJ2�R#��z+Bgb�`宻�b��q*��k�PU��_ڱ��-�Ĩ��JZڅ*"Rw����5�u�+W�FK{@�KW-��7)��%xO�:v�aV� � �1�e�ʰ_i�Ն4�z��>P��Ri��Z�x��wS82eN�o>牺f\�V�b ��j��Rՠk��&`l����k�_���f�M�[��iz�!����y�\M�r@/h���g(��"यabɢ��:���D���jH�+{5���ߊ��s�Z���Fn����7��S���To��&�^iAD����IA��t�f�%�Ò�~�a�L���Dp��~O{J�h��Z��f)2�3<�8��UD�T��9�=_5���� �Vsѷn�I�b��m����i�b�u3�K76ч�%��:�
����6�Q,u����%�͘&��KEl�S�I����FusRCy��R���L�#uz*�X������/�>g��Z�rQu׽ʬ��u���+��IS�jPW��K_6H�j�2�Z��J��\�2��ޟU2��W+g���4��oP�#�V �N}B���~�2�V��R�()�e�2���Wv����.�_���Cz�,��ޞ��p���!�)}'�4p���������{�e��;�H�$b�nH�$J$� ����t>����Mkp63|o&{��2D�%Faf�	0���V�����k8��C�"Xt�)5M�� ���>wb�h ��4��*��:j�Z����l>�1R�`��MbX��җ�e;ߘ(�B�t:g��M�q�P��qJۢޞE0�Z���Ψ@mo7��e�R�G\2V�M�W�ڎӤ��@t��<�7
y�f����Wu����m�}�y ��D5�?CC�~���6Б~En�?�㷳bQ�H� �|�P�%���X)��n�-���$q.^�x��~$x*��v�җ5q�d\s�M�I�:s�G.�RV^�s����K���e��v��U����y�t�����f:7��n5H���f����z+����0B�� p�5Qi]PmQ� LQ�H��M���&��:k2#�5Fp֑�l�w��4^���b5g�~��ѨC�m.zD_t.��t�1��c0V(�O:�J�k-C��A�%�A��`�!M�KF{k=4z?�2�2ig3J�1��3`�'Ƙ2g�hݬƦ�Z"#�`f�	������(U&�w���2D��a��7Qs�z��<�#�(<N"biʧj�P:�Y�^T,�.���'=�����:7�ЬXd:o�q�?|�n�l�O	m5,�F�5$�緟E�b�w���}p��K2�5X��.��0�{ %b���KX�x	��9K7(��6������L6/������u��/!�l�25�ezG�N�����>�3[�NJ�׵����}�4���/ ���1b����vk�e�������P:0��}nLb:)1�v�
�����r"�R�JGG��k��e@4�k@b@B$0���(˘���"�FSm}Ub�����.�/i����t���4QFUI���b�6�d�:�0�9!J�Z����7h��4�CP��ڄXЦC�\N���j*�X�ꌈ��	�����HI,�,k�����r�&f�h@�0`7�#V0���5/_���Z�	�)��ܰ��~���|���;�n c���rr޾����k����yR�e�i�Z\w�u<�Чa�#W'h1�U�V�ӎ;!F��G˕���W��j�� fS�5y��=�d֠!bbD�5�r3Ǳ�D��מ#7ș	����@���5CQ=��ӆ�I[u���^#��g!�8p?g�5�X��n(�TM?�#�B ��Z���?͑�]��k��o�c��ȗR���hFMt}��B���?―�6����9����_��E���Z���]2�#����m�_����.���N�;��\�`I�-�{������n^��C��'���9�(eIo��Y#Z���i}�V���Oq��v�����5��ܵ�L��BRcUa��W�����M/�q����yF�q�j��կ��~�x��l�׀1U�I�KS��Tg�!�%;,Y�{�����x^�o��������?�ũ��jQ:� �a4t;���RzO�EW\�i/N�+F��`Ŋ�|����ɀz�իW�l�2P�1�F��w���Ѡ[��1"�j�UGtm��orJ�SJ�2��jSHz��MW&���U��B_���3�k�����)����%T��K[�j��@�V�P!��Ǵ��(���f�)B!9m����WM_�v�`z���tM�`������8�&�kG��g��l��C��i�Y��w�!r�cW�{�ox�,�'*3S�:A��7�?��k�YW*�r��g'��Ft�ވN��	j��X�p���3��-`�=�s�Q�%7�80r6$�������<����"�x��0N�� h�LE�$*HU����=���#�s���S�V�x�}�����w%;�Y*P�k������+���͢8��T�ZE��kņ2m�$�H舍����o�y	����F���:�����>���D~}���A0���ds�l*���S�����o[ͪ�o�i���q��|��s~���9 #0�-ie�	�VtDɕ��O���}Wʲ��,��t'W�t'A�}���4�ՂԘ�%
!$�Һ�3}�f���6�H��?�]u%f����$�R��jĦ������:�+5�p��w��/}k	���Dk��s߿���eW]{���.E��"�jHSi�V�:��_���p��|�K���JP(c����߅:T��c��Jۦz�:
U�E(%���dJc�P�� �A�4=��!�������_�/��G��#���`���n!���Z��7ˀO~��|����R�x��|�������������c/
)Uz�Lju�o�	@P�K_z,Y	�Ϗ�'�:���%|�N��Y�1�J����o�o�y,#�r�	_}Nj���7ef�SU���i��k�~���|����'���>����W[��h-bRU.�7Ʃ�����G�c�X	����Oy�[��U/x�~��Z�'�غy�����>��3N�1:Q�8Q0q�c����׿���	�2���uS�j*ƅ,�����r��Qw�H&��V[g;�"��Ol�"�w�3&�!�D�K��=v۝_��l���ƀW�OF�׿�;�&�>�W˙g��B{Ø8l�Xp�yr�y��m*Ϥ����k}Ƃ����
_���X�<��ް��u%�/����MX{��Ұ���kC��Y�����M3B g��<,��}FGF�J{؀����ć	�
�,煇<����匟���oY�cw {�"� �ȴ�����qV]q%_���.�AZ|�7���^���/|.�1S��/���܏���??���qO=���ڝŦ����5xj
Q7�g����JӜ�AY�nq�ӞĚ��p������Oz<�}̞`��ϭ�]�;��v����r�x���H�O��i���u,Z����W*������P&��(Krg���������)�9��V#�3�)��W�et����������&��^���@l_��Zg-w�u7^y-ލ1���e��{���{���z�-w�up�}�s�w��r u��k��o�w�\G�=ڗ*\��Jq�F?�A	��0Q,%���[�Qbr��f�u�9��[�	=�mۍ4�r�e<�Ѓx��E���o�}�:~p������81V=6B+F�~��ȁ3�48*�Z6�����W ��/EQ��oԲiH��3HQ�:�H���z���޹��U�y�SU��K.�&$�0�	�$�\%���.+��"����,YPw�uE�Š�
���u��<,���"	I ,�&�1�'��6���>��z�8�{z�$�����<�L�=}��9u�������e�hX��B^z���>�|�94PB�~ m�o��_�������G~���_
"�ŋѡ�O��`�
<c��j����t���}�.E|N��5��7i<բ)�9zI����b)	(�T���=.�NL;W�Ҏ雕�4�p@�J��ϔ�:���Ͼpش��
�&��e�"�4�!�r ]�|���-��ʓ�(��	t�J:��Y������/�O+d�<)u�y-ZDO�o����*%,^���1c㈁P��|dqZ�z9��m2�*�Vyn�Q+��~`c�ښ�Qis�0׾v=�j�g��??�O�#<�{��\��r�#?6er:���/|R�c�Of��A�`��)�[B���5"�T��VGY$��N=f���'��x�����'��{$�Xm�HD� �$��D�j�[BFSR�"�
�O4sO9�x ⱅ�P�ϣO=I��s?��	�NP��~!�K���>���c8�#X��zV���TʈMh�:@���I�4Qx�[�.=��59X����I�H-V�6WM�w���Rc�u��v!D(�K��n֦+�"�Ǻ��y����K�謇�������ׯ'�����[gY�~bҤpk��7�_��Q�#0X� �G�Fp�C�x��n�
R�!;8HZܠ�����kk����!Qt��a8xAH4���Ǭ#๕E�>�OhV����_a�C�0e�ɴe=���xB�ŎN��$P�$e�5���HO'	Z'DQ4l̫�-�ZKb$��(�g�A���)zd��H�/�N[���<��|�L���
��b�J��h�1�0V�Ϛy�ϛ��$"�e��s|�4�k_Â'�!(��c�_�����7�|VN4=�>�P�X��d H���U1!��q]�	«���f/���?r��)0��#
�n�N� ]>�KA1�#���D"�-�:��������0���E�EFwC$2��ѥO������E)�^cG����ڵk����y[LF+�O'bPֽ������=v�ԭ�J���^�g�T�%O�L9��Mspp�c�����6��G;�	#`�cK0 ����7Y�d	���91�k�(�����R�1k,����'1�\�:~m�R���zee�$���#f1a�(�X� ����xf�� b.8�r@��CtA߯�H��$FK�r������E��VP�G���%�?���y�%�KXSFH��+���
hy!���2��I����s�/���	�IZ+֢N̞a�Tt��"I��]���S&�\�	���NY�+&+�R�%Q���g����<?�o��Z[Z�&7<�>(G!���u����kn"�6*�I�ȑ�<�쳴��qꩧb���l߫h��
kX�p	o���M���>���'�������W�����ڂ�~��nS��m�8���.X鰽�y9O!�G��B>ϗ?6���\~1W_~1!�v�N��!~:&��~�BÚ���5����c�=�4JJ�T䄏@E1�R�O�7�J�h�
k�!S�<�^p	!�+�]ͼy��A.Ȣ]��Ys�0aĽ��JA,TMV��++$��
��6H|�}��8�>W]q)_��I�B��p���i�(�	V	°L�kĈy?�;W��>�P~y�B�q�| �&�N4�\�X�����
r�)Z^7Uڊ2L�^�K���SO[���>��<,B�v��P�w��������k�.��k�&lS��i�ۺ���ӽ�@z"_��＇uo�R�$:����8�����Y�l�{�f�!gŊ�u�]�Q�����(��"�r�[�˭��'=a�U�߷��F�vg�D�A=���3s�
�g!�v��b�>{1mھc�&�>	�+	�{�j0���W_�"Lb����!��VH���b�qL= @���Ҷ$@(�?��DN���IPB�H�#�)Q2�ȓ��gs��Efj��������2�� �RȌ�jR�1��>�:Fz>Q��[���y�a��Gw��k��2�FQ�/��k��=Sg� -V�T5K�EG��{Ρ���X%`��tA�K���hE3TA�y�(����6"�;0Q�U���FP��T��v](aY��F� ?��nּ��"�V�0Hr�z��{<���
w�q.d```X�m��Y�S@o��G.�;�`�K/�<~:IR�Pe#�~��/���?�����z2Uu��(J�T�V,f[$�Ԙtpؒ���^;�y�Bq���0� ?���L;�&6��G����g2�#�r���%Qu�x��	E.�㷿{	�p��Hm�O�V���t2Ȁ�/"��<�M�ldũ������&|b�������3�p�'�:�Z�Ƥ�O�������3}�'Ԃ�C|:GcL�N�T��Ϟ�����$G�a��p���sЬ��7�t&�<�I3?ɤ�-s�u �{�ǉ�2�@h=��~sǍ�Q\5����;	�as�H �L��Dj�-�³�kwE�toh{��+0����0�I�F8��c]$�� Q�U��Zx������#gN��.�_��[(k[郕�L �![p8�⃝ɺƺ�^~r�ݜu�i�<pu�%C��xR`�d��&C/^�˯���������׏ ����>�}}���uz��`�e�ȑ);f,B
bmS�f壅��K����������E(���wpppؓ �$��+N<�x�(��E�Q��O��	�ϢgV�|��L�}4�����Y�b��������.��;�)�8a�Q|��i�����b� d�%Zk)���J��ZH�P��-'�>,~l	�*ЯR�:!=b��%�װ�f�9�1����ruH�S�����@j��<1��-�02��Ri�.�_�XT H��ēN$(�ǥK	�G��:?Gb%!9�<�<���[�2�ѣG��9����ɿ^�/\ȓ�V"ȑ�$�@/#}E�,���F��X4��i����!��JFI��6��?���}�UV��.0��>�-��ϝuFqm�����ok�k!��2�V0.gt����.�z���)�����ѣ�8�#�KC.�C'1��D�J��f��}ң$1o�����{鶋�$cǌ���)�1 T5��/��%���z�E�#�0^��y��b�����988�ӿ�$�ɓ'���+�_�/�C5N"��a���"t�g:8�c�q،�<���t��z�\w�)\>�b���b2�P྅�i���)`�D��G*�
�#�Z�<S�݋��ˋ+�cyG[��-R�5��C�|��̞�?Gr /?���Y��l���r@�Y~��7�mi��_��EV����$z�V�B
H�&�c�~mZI��]x�x
��d@��GC`�h��i-�w �͘��KhiދFM�����8SbI�� ���˟��K�F�F��y�b���N@C��R	/���Կ3G)�)J��x���gNבh:<I���ZS���?6��+_�B�G�:��+��KLa\5�n+$R�^�H<��3\���yj����/4�A'U�
��i���1&N�q�n��ZjK"<b�S�$K�Y����ǟ]Fh��$F�5����L$q���y�}xhɓ$��H'	I�$��X�yp�� �{�E���#�殻�沯��ʗ#���uop�-?��o}��E�(��5s���0�(�6�q��s<��#P�#
�>Xk�ė	>� ��O�{!IbH��SլB��P�a	�5�iB�͒O�Yx|��><��iB�Hk�e�@a��8������9瞏�K�?0Aa��f�Q
xd�U�=+"jݫ�"a��w���k�Gz`��L{NQ�N��BF�f����gH	�� ���.�7qY�����j��BZI��wY�Y�٣'+�IB��o���c9�9�9�C�{��� �H)0f���1Yb��02 �`����W���x��^�Lo+ FTm<��b�����Sv��A�]��;l|��� �M�miZ���I��
	�h<k�lV�e}:�[P��� �%D2@�J��MR�X�a�D�4_��-�ќ���=+r`=�IId,%C`��I�S�9�4T���mƳ�o��J!RN�I�{!��e�QKS-0R��g�'y������6��2�sZx�e �l���B�Rn$v߱�r�uv�|%�q��I�o��M�-�t�#���(I�3*�?"Z��H^��M�\���U/u���'-^��
L&���Չ���
�V��!�8E�:f4��Ĕ}' u����jZk</}���Xݹ��Y��.o��4@_#�B��[�V�6N���#���:쉨?�K��8릾��\�\�*�|�x:%XFFh�T� �5C�c���� ����	"ʸA �՗�"�T�"�W��gOUȞ�H��t��łr�����#+s��F�R���=e6h�������'Il��3�>ʤ�W�'w�~g3K��D>�T�l�������:��F��-�-��u������TsJ,2��ι�ʉ�wtN���j�.2�˯�ӕ���(���ؒ�� ��i~�T`�|N1m�)4�=����r���("�"�x�u^�z�εk	���Ā<��$�2��v�N��*IGDu�c�e�c�b����i�!Vi?��P5��\zi$ʤ��D���Z�*��HUu23�)-(�!��ʊ�(���URY+�/1�̎c�4ʈ���~O�A2]���hs�F�k	l�s	Z&!����Aek0Ri�И`FDm����_��|S-M��>�;�t�\Q<���;����t�)��@bdj�������i��Ȁ�J4�w��m��Ҫ��b�.2��QeR"Z�8��4J*1�"�G�9y�@�̠b�0��b�%I4A�3�(飱�����F1�i��~e �ȉ9"�����IDn��hU%H�U?CreF�M-� �4"�j���6���Ρy��9�s�Q;լ��mH����7�{hD��01��hx���Hl*7e3������M��[�]�Z"j�h��֒VaMUWUY���%-H�S��EM$HJ#|����i;���6�9e�B�":�6Q�̩T�K�/�BA���3}e�S�WNO��*��E�j��Ҵ9�u���j,j���؜��!��:��
w�͏JU}��f��c�yG�����8��J��F�5����m��\��=�-�R�w�0�F����d-��"oz�2��uC�J]f��F�R�
�4q��х�-�)�:��څ�M*�H��r���}!�U��eh:�ү�>�|ek9�Ū`�EN�E�he��lc88888��^��!��.ҷ}�����\"Z�+�ͮ�Z�9azZ>���ӛ���2�qUN�a�M#��j�,�Gx�HI�^_��IǷ�=:$�h�Ȣ��-߹!6+
������!�i�j޶����|6=�˚�`K�0�V
i9�}�A����MOMۧ�:��-#�[����Ky��Q���~�
ZZZ�7��S��iյ�g+ uppppppp�ii��wL$-%��$��sWϻ�'Xe�$��%$�@�}׫M�]�~/w*��14<��ʉ����_�-OUA��\.��R�&)�J��������aGCb0�`�J�[�-tX�gtS���s�񳦮�a�¬��2P�6�	��]�mBD+�HBhZ���[����Z�W��&L�RM�����q�Q�!-R�(*����s֌��o�ݚ}F��PT���
u�d��TD��2k$	����o��7S��k�B��a�����uppppppp�A���ǆ����\�տ����3O�
k
�n�S@��rj�����U�H۔�V�� �ҔZ�w��k�����x� +�T+�D��]Wpppppppp�>�$��@���l�ܣg���U_^�︆U�4�K2X�J\�0����n��,L|��L����:巏,j�j��IbӜZA��!/���opQ�f�f�e��6>�|��N{�۩7�翻������������;���9�o�Pf��,���I��d�����.��d�H�j	���ȡ��[�%�]��v[�d�h-C��g����~p@�ŵ�&����X�<0�a"�Flލ�4uD�QGDpDԵߍߎ��D2=�J�2F�HLYjM}!������K?��5c=�.`Y��l��݉(iqRC���E0�{܍?�u��rDbh��ID7��<**�qg����m���,翣�]��w�������?�~7~�zdT�&���|�RKV���dy^�O�r2_���5���[��a@�t��t˞mm<�݉���V��,�-4�43^}+i�ɿ��+k������dTm%	�����ﳍ��������{�.~��{���ۏ���n��i�������*c�kd}n���}�����!��2��
���:�(o���lG"�1�W�[���ݚ7�X���������a'DYB�H���?�� !� `W)�    IEND�B`�PK   �i;Y�R�� $� /   images/179c08ce-6e18-4019-8002-932a24469ad1.png�z�[�a�>XJ(*�"���� A�P:��0�]"�HHwwMb��Cr��l�6`�o�}�?�w]_.v}ೋ�9�<�}��|X�k-eJ

JU��:$$��HHn�ݼA�S����p�榠�w���w���wrgc7�⋴�NO�p��������{w���	�s�YY:�8�ڦ�dHH���|�畱��s7���8Yp+��~b��x#�񋈻�jIPH�i43l�q�Ͳ�SĚ�4"^6^DRd+>�[��:�[�WJ���=I�)�C+Ocy�;?(���(�x��ZBD�$��#�e�0,Y�[曽�t?'��|ߌ�D��Y��2���I�o͕7`�6`�Ü	�����`���C(�͚ɀS�@��2�͸�H���j�~2��g��s������n���������:�#���9rHC4�NM]O�~Kˌ�S8_>��C���d�K%I�:���*E�J�<��:��1�u����o�}w1^��o�gx&d�/7 冞��S[օ��*�$�o�}���J+m��1�b���~�`�Q��&k��#W�;O����s����X�tyt�P�2D�DB�Q�ș�p)�R�!ߙv���ZJtc�.����}��4�e����2w�(*1�l�j�['?Px^�h��WD�8�v��qoJ���D��e�IC�g-��'���VثJEVX	8�����d�Mj�e��=/;��R_bK)��u�x��Q\�[W_����u��PόH��m�w�!#dT�}�N�hm�]����¨!��`i��� ��}����{h�9�a3�eHud�u�4�K-@mɩ�����]���I/r��Q��V�tb엑��>*�O>_;tT��̯�.������+mD.�H���i�l�|���a�\{���U઩<���Z��JC��
�py9D��h���=��R�h�_d��_�P*2�e;VE��iڠW]�
C��	�QF���7|h���A_�>�s���m��i�P���s%N�/Ūj�m��h۲b�-�Ώ���t$3B��v�q�z��w�H7	�By�y1�i��v�S������ߺ>֟�Җ��Bm��gx�I��$�|~L�{�[R�e�G��J�������^Jo%�J~V~Fi�����������������j�vU�+R�����v�k��/�	�0x�{<�!
M���T;��t����P�6�+J�6�Il����Y��ρ�h��O1��#/�ݦ<~�H}��^��(9���OɄ�|	��j���P0c��t���4J��ω�#';��s�޾�7&N�ط58�IB~@'O�l��<S�4�N��1����Z ����Jr�� B��DlR��a��`�}i�m¶ַ� �g�!C�d��N�&�����u�t�������[B�|ȷ��6��Lb�t�ַ[�ʀ��c		f	��ϻEfL@N���qx�~"��4�j����k�n$#i�XW�^9���!��M��S)?��RP��(����a�Ύ�*����T�4���7:�e��š�[ܶ�4����FP+���d��{�"�$S��L��3�󿲋�s����g�k������	˦Z�||�ܕ�k�M�7�����?�Tj>�}-��������@����?9k�<\C.O-�X��E��Sc�)�8G>{�x�D�\��u;7�14�N����U	b/���a�)'�q��"�[�?�}����謁Ow�7�lr��i�����G��1�������]����{?ƏL�1���	?��]q�Ͷtω�#��p����(h��:*I�f�W ��3���ښě��݈:��
�$��̿}��k�4�g+G<�������y�_��4�Zz]�y�$� ��Y��Fk�>�Q�-7봃5Ph�Mg(��(�@�G��ݩ& �I��S�Ҭ͠�U]kɒ&�X�W�����Ͳ4�֎7��O�lB�|鼒r�m�]T��M��z���jP�dx���35ǚ��郁{�+�C���L
o��ezC��&�0�z��B�"��}�zi�r9���H����s���EΧ���Nu�B{�rV���4C�,\��.��)9!�[���?.��+��?&�B����w���,MC��f�_˞����<�8 2^�З��S-Y4��[����;Vk�Jl�9�l��Tͦ�z��n5܃�����i�(���B�/�����v���[h����C
���m�1�JGӃ�-�= ��Ԣ��&(	d}��� ��_u��&v�_���F�VDox���^*��_�ER�� 1�8�O��y��+G�>��lpq��ҋ,�۶Y�2<?��>`$������s��[4��eC%e��{�0�m�r*WB^�(Zr�CFk��퐶�=}@��j�ӫk�c/���3b0|�>�7��n����z&@@���5��ڒ���*q��;���e�7%2>!�1M���:�O🸈�|ƶ"ĵ��:�Q���ojV�F�!�Q�m�Xߦ��砎��|E���0����8�Fx�<�6�^�cb"���/�ώ�-8��V_�I)?�rܒ�p��W_/V�.�8���9<�����	ƒ1�����]�:9'u����f�YD�Bo+��wwz�uv��x�_܏����_L�&���L�^ -��Z����D�[�ˈW�	��n3��5��@�n����R�9�����|_�=o�9� �~���+�0z3�=��9m�Y�����K�W�HHb���* x�݊�5��N�(�%��l�{-؏��K�A�rb���v@r�M��c�l�i���_�Ħ���O�Gr�'h܄Q<��h?�I�(� y�X��8@d9���~�/��]C6@�,��ko��A�u?��cUA맆�57�@�y� j.g$"�$� ����q�����Ib�+f ��c���C��̽�?� B^�^�2˯���`ׅsMi �2�����XyFԽL�L�s�g��潓7����)!m�
a���s��|���eNo�*(�m�{;�Ϫ%�?Q�ǭx�g�a{����	=�LHg# ��$4\�^�sc�cѺ�*sgti�*0�A^^�3���Pm���������%���?�n)Uگ������Uku/V���B܅x��@}�ԶWQ���%��ZJ��3�fe�@*�&v��%.�r��]��F�SmH�m��,<�}/���F�-�ukgV���6�Baׯ��U����*��j�]��o(�I��$Z)�����jj)�]���W��z'���]&�ɣ����<Ęj]�8�p�K�SSS"�p������4��V����.I�4�oZ'Se����%�7?�"W���.2����X}xSHƹ�Ъ!Q��;��
�L��F��Z���Z\���N?Ӹ\�J�,�)I+˴�*�4��ſoJ(s��?��V��I������<����B��7��p�A�͟ô�������#$m�
F��g"� �����v����>���������#`�E�xk��+͹�U�%����Y���\���ن����~yY66�MR?p�����V����r�t!TOj��ه�ZoC�وB?�Zo ��?m���q��������l<���DB�S�*��2��B�;!a!bS�-[��(v�Ԕv�VH���5he��k�O�-p�"� i��X���풏���/˟�i�eVؿ.�=�x=3#��ŝsK֊�O�Xu�L4oH���E&l��X����b�*�}����"�Ù٪�GzhS�E	�{+S�ƥ*�1�_̾o$J�=�I�ıE�n���jI�r)�g1'\f��ޜ���@(��
��ɤ�*w�>O�)�-B�'��C��L��ŕ�&3ZY���2�=��$�#ގ��|���y<p}_�3J:S�mEE�x~�Yn�����/]\R�s����ЍMa���&x���4�x�	dR�߰y+�կ#to<�1���L��S�j�������
�ﵖZ�iFr:I��G�����Z:��P �["�����{;q�%��A��"������)w��%�h��̎%��k�:13F&e�m��>�tBnn��qiԖ�ƍ�P��g.������UUL ��i??b�g3� �*��qfw��1�ٽ]�����
dx�E�C�O#��D���		��1J�+�a��Նq�L9���rx����bRի3t�Gژt��
�����N����6~�� g 軳sF���.�:ߗ�xN��[�dM����@�>|��;l��Z*��}�V�R86R�ȇ=r,[�J+s1���~]�d9�{��V-��㞠�+V�S�D���'��3Y���>�e�������k���,�T�p&xf�oȬMı���ætAoL)�e`0G(�����c����j���뎽��� �4�����^ws����=�d(+��Mē���+�n��M _ȿ�u"��g'�ʗS���V�l�p�k[r/�iA"���1��Ϭ��o.���Y���(�	�R��4cc� ��iPP��45�o�[�B*A2B#	�t�� �gs0�PAD���:n�j�:2)Ll��q.��/Lk�fR��;3�3�������*�zO����c���.�ߙ�e�n��{2oMH�n���^'�'��8���[�l�z�3��Z��4�-�$?��P�ޢ��Ym�s�-�n/�z3��pi[��k��@W�����������)e7���u�Lr� ����ǣ\H[)�K#�9��%���m��W��
��Ñ�m��Kb9��˸e�bJ��K�qIBJ&�r��VG%��ilf\>Re�mKX)D���oS�W��1���MF^x~}�V�k�h�x�`���E��I�T�Pl����{l��br��կ[\k'��;�h�&�ۓ��\-���ĺ����#3Y�·��kߪd�q&p�ff<���O�͏���3`wtB��lEG�"[Y�/��p[��4�}+.��	����҆���TȰDE���y�� ����O�8yl(C7�e�/��(�l��/�/�Ko��L[h�aK�]8�=��7�^%�o!bx���챲�H z	6���q��O������y�}^܌�[��L��E^ฎl�νļ=��9� ���L]��=�^���J���+�&�����f��hY�%�n=gRP��	'�vc������1��b=@F˓�;��'
�};����$�*f_��y�֍���&�~jvˡ�o���ml�&:��� �.q�g�s`�Y���K�o�掉��s���..?	":^�석{��%�>F�N)��1����	����|O&�Rqd�D}��9�V��3W6�1�;�������F����G�\����Yƍ��l]������P4f3?)��T��z�����ƪ��m������;�Hxy��W�e����<���d���g�z����Ŀ[�"fDj8Q�g�=�X�	�����`�mfh�����^�v �_1�@�Ǆ@s����&���S"�r��� �>ٶ�*nw��i��|��������-c*� F���ý�*f�1���)j�Z��u#��i�l�����I��	���)z�\��ޭ0��b�(�|��w����w}�,��,�Epl��w]u�tj� >"�޲HB*no�_ ��۟!�o_۱�43md�8��#����Xկ�4����;�v�{mcY�a#�M@ek��O��ʴ���b��)�L	I3�N��Ģ�Ed�3���))�:�؊0d)�L�mV���6�m����2��cآ�V����*�'��Ɍ�ꏈ\�#˸t��6"`�s\��D��x~���+g�<h���HԻoj|���J�0@�[�,s�j�Dtíy���B۸�m�pLV��{�[�3���/h>�&�2M��/!�>�|^#4�YqsJ�[T�TX�� tgh_[q���S�EE���N��_�P�Vn�&z��~��Z>�$?o?m�lO8:t�#}���2㏀E��T�@��F�'F�R3�eXJ�@MߟY�W joJ/lr�J>�/h0���>�g��|��#h�r���9�e�Qlrz�Ι�j v@�AN�P���=U�jc(S�}k���NJrϩ� �cG�/|��Ouԩ��I�'�E���DqLD�$�����Ü՟�C�B���=x֒�K�堟	r����s�Z�cɷ�#�aPxy�@�5+'�?h/N4�c2j�"��H��k:F��N�i���J��>_k�p��A�T�]���wW=� .-<P�L�%Wa�	И+��}6��ǂ��g��*�9��?�5β=J|���7�蜋MH4�]f�Ԫth���$*��*%��W�1��A���3~��(���Oެq�=��R�51�)�y>¼LY�q�K�U�$�K���^�*+Y\�e�*	s��|*5�6=� ��^%��6o]��؍���aOsy�boRB�F@�e����B��$��~�����0��+�H>?��8U�yA3���˓� L;�xn���r琟��s�.�3���"��1^̸rriu�A��w��l�	�A+To�c��c�;҃������]9����%_�V�^�|&��p���#l�w��k$�?ܓ�[���!m���X�rj��#0�X��|���Bˢ�ëMF�!ι�s�ܨ¿��]a�.��B�\��{��44�&�����l���|�]0��Jrؑ����$c�rz��D.�MB��

�6T	�����1Y�3_��� ���K�F�ŝ�}N�R��~�jQ^�&&�-8�|����K���N)�omo�>��-��G��X$ob��@�`����n=�}=y)�=�j"���A%���//*F���pC6_�N��yPf��X���'1�}�3S~�w׿��5�����g��T�\�[���_�+6K�|��"�b��U|�B�����?�~�
�/l;�o�|�-h�D�H>��*L/�)\F� i����x���\͈D���xzs^;3s��r�G�)Y����K�+$�/Q�!�p������}q���9-M��Kk�c��sG�i�}_i��v	]/�G̏��L~�(� �h��W��:�Ϛ��\�(�8��r���#�$���4�04�%av�cZ��jq�?�k���ͧ3�9̫i��g�Ԥ�Ot��-�߰��|L�]�!i˗�v��gēe�[I����;�����n�Ph?���w��f�bE+�y��ch�����9�!7Rv#�yW�.����P$}t$q-hN�QFu�,�p��f�U���jnFѵ�ٺ{���o�4�}[{_����%�-6��1�]0P����N�c,�߽Iv���?�_^L��@�:%����'t�w�?~	<;��_�`Ys�
x��ӓ�h�O(-I]��i{OO��K96�;+��sVX���@�Ǣ4��7gc���:�@�'������f�l�Y��w��.nLv�?�s���6A����� 4����</&h}��3�5z�h���i;����V�mQ �S���u�y����Y�;���jE����ư̿�������{��b/�w��[t�̀�xb�?h�)~t��+���N�N�a�g2�l�ڥN9�҈b�(|�MФ����la{�������eIY���Y����T�%�;7Ь>%�~?�3-ϗ�v���2�=�HH։��2g�P��p����F�r�Ys���3�̉�3�����f=��E��z<�V5q�*X{s�L������W��2����5�q��D��r='02|>� �ڈcP����V�	�]�
���T�z��ޭHQA{�'m�4���&+�c>�n��(;Xp������1�v�m�iIH"4�	�9����}R�����a���;�?�'H/u��(�R�ꬲ��d�p�>���3TM�X>4���g��U\ⶳ-dhO3H�N���(sl��<����~ ��k�:Q�E��G)��`O�b��H�XIP�H�f�:���~���Ox>�9�OQ����Y����K����o�_���r��6�� ��K�mZf���xq��:�o4��gd�i��pD~����;i���{�u0N��=Zy�[V,
�"� 2u�R$8�������N|~�Fr��G�0��ar�A���5�|�<#�2D�ͬ�LL������f.���Y)o�{�ڊ���;c���XQ."���LЪ7��߾8U�_��G����]Y�Dc��D8�׵���VY�Z��K�Y�A��X�R_�;�>j�K��VT|_�m���H9��y�J�!�L�\���7k�ݫE��ۢ�b��;?�J�0����\��ۖ"�\���N��{ypd�nx���h��3�yJ5Eg�)��VN����{X�_���3k��<?L��w(e�BD���S�]<�cZE�Jo�:��jC��Z&���x>�Z�����ǣA?r�Ի� /�6�ԁ�,m�������_�̱հ��� M	��� ��G_�M2����+�J������e����ڎKe�k��Y:��@*KT�\g/�7k���6F�;��*+�777׹o��ԩ888؃@� P������TIR�U�d]++����oz�C=��I���_�WL��Y	� R�f�n��~��wTK�������(�yH@%w}�W�/�����SWL���?����~�.`���ݱ�Z���-&,�6�'��5'�)�o���)�Z���ȑ��t4��r�"2X������"۠ʬ4�����`m{gG����0�t�D��ۆ�b���|�@��/�_���{��O���f���)��Q\�M��=h�y�'�*��K��7O��Bt3č�Д'y���JFC�Qj��H4;R��L&�ԭ��H�k��+��Rg���_6JJ�R#�0#�X&�}�r���}��ƵJH8~�AN���CCC��W��;��m�p�q��,�ƺg��o!xg@~w�H�A�c�r]DkE�wZ��³�zE#3��[����~V�#X��4R����۴�oe(�*���������ǡR��s6�R��߁lg���_rs���߾�'ƕ&J>�gv;�[/��Med���������R�L{Z��bNC����6�#��{�^�L\��z�qn����\C��F�߂9MV�"��[�L�ڊIH�dJ��+�GSEl��ٝq��7��'&
��I)o���bt���՝�$M�6��8���&=Y+�>R(bS��ȧ�U���EC9�	f�O(t/�r�|!?�f0z4C�b!���)��啭���ܱ6���D��� �2���-s%�"�b��-%-u�}��fN(B���a�J�͠�L˻dMkj���'[I���jΒ{fy���f����A���|I�×cL�
�W���bf.=�2���L��ܞ0��8�� |�=�Om���u$$��ú�n� =�۰P%��mN��� �������Llvƾ���6_ؔ�����;�cƻ�Y%��Xd���i�1��A��IB��"�d��</��_���cF��>����+�g�i��uN�;SG)��;M�����O�	�w�5ݷj�����|�	�R1+�5����C:��:����HE8�� w^��$�]Mn������H�������<]j#ݕ�yac���,�,?,���
�����h�j��P ��ŝF����*<��7��$`� ��77q�@_�I�k���� ~�f���aQ|�EGfYEnv�y���w���;c��E
p��(�U��!Ov
=[�q\��#t��&祐,_��?�0Q�[�,P�!TAٰO��\P\�L8�E�в�)�ʘi
�^��^���]���i'�dm�f���*t��2&C�~{�m/bT�HP=>f�����U�<�h7�1�P�R.U�5��>�*'ҝ�J����3큁sk���0m�W;��}�����f��_�ո-^~e�X}�1r�v�K��c�|�2�����ϜӁ6K��W~���[ِ�C���5�{�x�T�@gy��V&{:MF�Y��	5@�Fgy����5��\k���o�R�Y�6{ �:�^6w�+$���t 
��N��*8.�p#%�,Y����zB�o=\{��,�g	A\
����R����_�X�tೲ����V�e~#�f8p�.�^j��c�6I(|����͹�w( ��i�w�g7?���Qv�evY�@,��r4�S{3T����c.�JJ��S�L�f�� 0p�4l	]�����$v����lbf���&?q��vN��$C��2cw
�#k
��6x��:�UT�б7Rq���47����S�~e�����״I��0K{n2.�Q��<?5&�!�J{E��dd/�c��Y'nb��k!��~��v���-u�P���Rއ.B���W}b�E�]�8W�8��^1��#��7/�@	-!!���5^k~�!vq��7�SZ �s���"�?F5-A-_�[�^�gZhz��4�M�9f*��"�P��J��g�X�Q�;���ĥ|������*Ͱ�і�M������]�eJ�q�\G��80���ӟ��H-����RSS�%��xf�Yh}��b��N�m�U���0C9���;��U�m���ڸV�5�p5��5��������0N}�A�*;������8�������)fg�+h.�����2|W�(�|Y����<�g�P%;��R�
[�p�����������;^d/Z<�H�,6WD�ͧ�>�~�K�uZFƸȰL~;�>��j=�Vp�@,�fJ�`��c��{�e��׆t` Y��o�6x|���ܳ瘷���:��	O�\�(��W&���ې�>��q�n�,����/�u>yG��y!i$a���٠�j���!K"?0�O���?3����%Of<f�W��y!o�
T5q�K���p�X�= ����|TW$���A�������أ��|���t����Ψ�s�˰��k��uH����V�d�:�����n��0ú���l�4TS�,U�5%�5nB{i�
Gg�R�tR�`	N٧���m+3b��i�a?���ݢe� ���~��_<���ɔE���aͭ�����&�81�IU����8+�
�c�ȵ�H��h��Rn
��=�,��:{����z��?���}Lhl��m�0��-�r(T��<6*Q6o-��c���@#c[��oO��~q�*��������S��Ui
s�?���Vl)c��Ǥy���w��Y}���ċ�����ew�3��e�7����R/{���D=�۬��㬭*BO��y��9NhpKW�:�f��?5�rq x��p�m��Ż��#���E���i0�~���A��q:7�Ct���,�l�&�����d2y�5���WO�k��c����o�zE?���9�O=�(fƼޕ�#9��x��]�/�GÃ>sIE���t��\�<�ǳ��Ke����(������@
��eU7�Q�0�H&�5�)]�o�g���t�[q���@��E����Y������ѻ���1pU��(:樔GO�#���)j^����Osp��/��k�:ں�� 	r�g�l玌���A-��9���k̡(7YG���k��5��6�1�ZT��&�˛��>$��i	�~���7���2��U9HI�<Γ>y��H_+7V;,�~������z07�Q\�߱b뤖c"�lb�o)�Wg���Ò)J��+���0>�3��&>��+����K~ʗM1��ù����n6v�p�Mf,���r�4́��U�Ù~yeR�_[W�S�ŝ'4[B@څ��"}���������/,"7�].�m��,t���X�:X7G�]��^#�76�'�1M��Z�I���TyU�zn�C!���x��9���'N�H���gq����7BZ�R�[~	����"�� UC0'�O�r7���;�,�x�<���c98�/�r����O���fV�r���S��!N)?��`�'<�cX�@K[���/�2I���vB�8@��K(`#�������s��<�(\���'�EjoVE	ک�O3(�YS2\�����?�ҙ�ҳǣ�ۙ�A\
5���syƌ7(���d�,r�ʰ��E�cH@PiJ�;�Z �����Zv�cwVcw�-�#ئ#V�� T�Y�A�E�ak=�>�Оr`��Y��aZ��!��[�i;t�N��"���)� �c�r�oZ/��1�z��wC���Rp�c�^�.���ڦ?Y�%o��Zj������+Q8ʟ�}�`��P�^eE����0�����[@@ ��㉻/���ys��~tq4M3aX��s�"���U-��J�#��Ƭ�E@��^��,�r2�4������Fa2p�~ᡩ���\���qUYYy���-g0]�ۜ�r�s�Y����]�M�K��Н7�i{�sÛ놬f�㨀�-akc�j�Q�c�z�n���J���ٰ���	z֜YĄ��7wn�� (�/�P�������t-�~����u��;��.X�	�$9�E4;��c��n�[>Q>=]�f
W�ݎ�,�'�Γ���8��t�����1������;�9H�Þ��da]�sY�y)I}�6z�?B�%��������]�Wks�����1MW0��1 c8U�䣉�3�l'ƍ`��L�X�b����z�em�+2�n�-&=� =���ɠ�m�-�r��Lm{�4�D����ҏShK���O��M��f��T~�*�9��U�=����y�&��p�4?��/���e���l,������g��ڳ,�6e���VP��d�of>��g���S��o�O�T�KZw��Yx�����az���3�`,e���"���+��|z9��^��k��,� }�{� ���hP�Jύ֚%ͤF:�E�j�q������,��)��3ulz�����������F�/�^�/�p���5R�r�����Q���r����<Sסp�ʦ�)�Ԗ32�D�v���m�, z���π��J\1d��fj���<��ڨF�;�adDXk<Bw~[&vc{�w�ۄ@M���o�qpx���w���ښ����d�4�AV%�L3��I�)a�ih��OX����&�J���p��'��}�-��o��5��>Mop/�\�&��|�mՓ8M4�9�{��*V����<;�A�U�<[7�����S�ǖ��̡'�a�-b�n��M\uL�l��F9+��!���ǫe�UH���Y�aZ�7�T�Nao���.ޘ2OyO�Kw�3�R�5ͅ��.���IO}!U.9�FZ��17%�=�������,�� c������u~�����W�H�
֝��[V�lC���V߲��ɡP�V��q���e�ǝ`�L��S���g�tu;ٶ�9d�t	4��=��G�xܯ)�yم~u���<H3��?����m�0�Ur����@�����#�öK~��֤$rG��,�:y�_������ ֣&o�ң����~m�x&�K|_�*����f���s�X�X�Ywm��]��i<S���O�&��CE*o�X���x�l�/L( ^�&���1�p��8#�S,�l��qo�u�Ot��M]\��4��jeV=m��9�T�����[��~���R�rxV��{�/����y��t�L��u׻�]ކ�#���n������?�����@co}��N�O���[n�,��+<?�5�<S˅����Q�2gۥ�B��}��{ukV�����7��>��v}�Y��B�aM �y��ܮ�8��'\#q��hq6�a�E����%�Jp��C5�P�=����qq3#����TN�����u������=��	��f�]���n��ƨ��&t���.��㌷㞺kU���)�R�n�>�6��F�߫7lm�+�xϣ���7���Z�����[��C<�O��<�7y����(C��'dni���I��3�W��e<X{�M���yx��q�q��1�^N��U�U�<A: ��K�,�v�uJjj�n9�b���0�����5T��q3%r^S��j�1�i�����]zɧD#Wxx�{i�&���_&k���QL|
���i�Au7�nf\:?����7N=�2F��2Ř㜍��v�����,�����m��}ZT�%�+�K����/������w����'(���!��追��tS,A�Ҟ;�.֝�ܹ���5���"6KpSJ��Y6+{��Բ����5C N*ך��x��ڢ�F��1VIS�B|%�rZ�n��!�{;��P��m*���� /t:��26��8�͵�*��'W���=~�u��̧#�=I~�t<~�^�^�\B^{8�5��Ű���8����{���*��ۀ�����[��Rfւ��BY�z����?�}��P�G��g�7	�P�zr&c:2�����Y��V;e������!'a���ϫ�N��tb�,a�5�u����t�x�ݶ� '�-�������C�i�k6�I��4t|�m�*@�����.�r\>Lp5�0=õ�L�:�(�p\�6��A��î{YU����_�x��͔��-�ž
Y�=mp���~^�î�}s�\�cQ�ٳ�������q�J6�R�,X���{�o��&�£�V��#�Cr%㖕5��� m���T�j+d����?%k���?I���C��d66��x2���f�)֘=��L��ϦB@u�>}�"�Q���vC
�����ʚ�n�pB7V�3Z@�y������<h �@ō��ʉ�
���P�X�a .�8`�w�.�XA�����H��ǖ�4!��1��(����Q&�PB����|�`�K�;��gw��נ��-/�G9ٶ^*ޜ��N����#�<h �q��s/��ϟY��^�O�ޗ�4Uf�Ou	�8k�*�LM��,���+����X��0�h��0��ؑ�:��>Z��]���Y����!��U<��j>\��x�?Pm�S0[�M�1g�On7P�5	�w4
��Mb��I;���*���n3�Ά[����mN�N�J�������V���qZ+��}am�] �mi:@�M�Է��ThY�r�L��c���g%Ir�_����b�+X7~�PvJ�k|�#߽!��a�>m3>�<�ۆ���cn�V��O�$O*��=����6G�`�恉c\3���ɚ�S/�G}�ǯ�F
���]�	�����|v����^���\������&h�H�J�ox�U�v�l\�A^e=">�A�mH�$�<�i�5�}�wL[��B5��
�8�^ �K���w�ʤ��:���S�[�:+Bհ}k��= ��U6�i�ъ����Q3TVM}5�%�z��O�K�!�j~Er�{��mp�5q>`	Kwe�g��g���b�����,��OD3�=�Ҵ,u�D'?XLT���@?�zw`�5ͬ-�W�A��a��_J�������]Ǻ���L�~_�I��)����i��ֿ�1��/~��r
�����{ul�m�V���>�I����,5����*�O��&k������`��w��L8��e�����
���ȿ����>}M�h{�?#'اrɇ��W3�����
]��Z��Ms�E�N�c)����S���ק��*����R`��ǇQ���V��N�M�)!�����OVټ+Mm��2��BP�)���@�ؼ�B+�$(��z}��Y�vV�0��."K3����Yߩ��~([�,)pU��,�(\����1���,��ۏD&ݙ����R�C>]9;N-�rU�5�"j��;�1�kv{���O�.����8�U���^��vL�U���tS֭�d���
C�22��]�)��y��
��K�K^��&�>/8�����b��^-4�5T�1ȸ���,��U�6��Ń��㐹<�*t�b�ʡ]�eb�������<�,i��p�W{,'���,F}^0�␿>��e����;"��^/hii]�uy�+ך�m�)lmv�7���:�@c�ѥ����|��Bf'��/�3�%K3����L]���e���k�%��"�v�e�R��5]�'#�cx�z�e��S�|��쎒��O`���g��pw)-K��O=�
��n��� �(E��&���7E���Yϵ$��F�>1-���n�y�y�2��7	FN�WUpa>>�T,N.��Һrf��8I|V�)ا�\Q�F�k��G���3�������x��d�-��l���SΧ��g�Q��O������&���$�f��6�x�/K\+E������xrV%�y�q�D�O1�q˒�bD�t�81�N�+�h��!߉ى�3?6���)ei����;��*V��Ff��n|+�����鲹��51����U�R���= e>C���lA��b�܀�₆�?�OF^��Y+&300�YuG7��^'x�k�NYg�������i�$��y�&�d�`)���y	���_)E�+��H��_:k3N�m��k�ٱp�|�\Ф��ǔ��h�oM��������X� �����iW��%����~�m3ݕ''<���g�W�����:��͟����N8L�5 ��r�*M���>��4� ��t�[��܇��AE�mOM�$�S�,,@y�}���Bl��@��<N�a��%���V��/�w��>,�a�&��hk������2Zۆ����%DZ����chD���a�:��������q��9�?�\g]k���JU�?�y�9&ȥU�Pښ�*-�D ;�Bd�$d��J�v�����g�x�
ߡq�wt�{͘��%�{F�ʵ���Lo�,VE���%�����������C���J�w^e�8n0!�ϵ��i��O�n�V��n���;����y�e�HJYѽ�̀����5S�c��O$���G���[�Y���d����R�խ=�>�f�O�m�/z��4�A��!ϧ{>��͕�?ܜ�{����~l�'����{y;h�L�ˎf5��u4�%p
�69ٻ������Wo/)�
9�:F�>�Yڸ�q�z�L�c������Ҡ������*�o��}N%�O{?T"c�#c�FaW����H�V���}���h�k�-=��(`��a|�o�k�t�_gT�O��,}P vQ�p�+(=�ٸ_Le���gRtV+��*˳�vD]K~������4�-Pa8!����������/��k3���t^�2��3!UӮ��������M��gj}���;�T����v����S��x9�ي��w�OC�#�68P��o��󦐪4�G��X4�I�?/�SVcy�c�����C	��1ڼڎF�i����"�t�)�J��U=꩙����O�HcB�O6����^�=����
WCf��Yony��*
1�xC��Ť��Kү��b�yE�+�o���gM']�)�PN�J����^�����������GF��Hǎǫ�a�~]C=�D(Ҫ��,�a �����K��T�i��ҕ;�0%�p��A/�0��?�u��Ms���9g�����[�
�|rj,!|x
�`�ǍV��6\W'T����V��?&�|���]�!fb�:����0{{�Z4H'�����=,s+�6���'�A���N:�Y��<~4���b�@aQ����H�:�CU�{툃��o�$���g6ob�}���Eڸ�{��g/���"o���
a�Un�'J=ɗ�)�3���A^]ǿPx��p;ֿ]��G�|�9d�9i�j��7�M����;')����� ��)LB$�de7���v���lt���.a\�5��q������$0`�r4�~{ᤃ��l\�[r�2vU6�&i�|,�����ȯ�F�:=�m�?�����x�>��{��4�&� ��jo�s�����"͋�FNwF��l��u�=+�S1qY�+dC�$�f_SB�4��u�E��~����4��/lGǳ�c.�`:�>�q�����r���_g�gQoy��U�sI�;28}�v
���������,�F�/�\���s������);쾖?Kfk�y��ZQ���j�x"��C�/�u'�G�� RB�{4{#�[���Q�ͭ����%�ʩ�8��s��������^"�xk+H�\�v�X���N���X��b��.ƞ7n]%dk�#���k?d<���}��I3��k'��}����s�+�iWKN?�Ok�.i��I��(	��Rӱw?�Vh¢q�4����Djp���C��C�g|�@T$^;�$n��>���kM������ok��fρW+#�gbt~�Ǔ�y����y�Q0�b��	b��#�����Xo�]$�n ޖ���L��RE\X��D�(	i��u������dЙ����t��oe��=:�����}s
s/��V�Ju.˯��u4�����:������$����hiAOߓ~QS�Jx�Y��ͲM��8�k*��I#\244<��;m�=T���q��zc�v<�m�ے�M�r�������NZ��PSq��Nr�����n�>�F�(I�`c��R�)���gaZ4�Y�D��8t���в=0�$er�p��,G'[x����@�ֿ��RH�놕�M9��Lc���=�ݘd" ?��Q��`m��n�U!��|��x=��*�$�瞇ү.I�ʽ[�I���5���5���s�8��s!�V���Ե�J� ;�5��U�*�!K#1;��[s+�\�[݆�p kMN����䎏��~���~��3���H&<�=����B�*-Q��\~��xk�sr�ق����Y�0�ywY)n�9���R�����C�G�:T�9��l��5,��[Ѯ^�^}<7q�k�@j�
�U�]�.�w��4Ɖc:��-(=l<pi�~����b�'A��	�DL;�����װ�QLL���&'E���o7�e�܅b���74��(~�8c^�'����@[�yN(��,=J�/�K� �� �/5��J�7�0ˇ��;, a�����m� 3}�1�։�ܚ�Q-�ޙ
;��ϑ<�ݏ!������K"u�LXZV!  ��(|��縒Х���hC��jW���*6iJq�[�.L�w�d
�1�n���a�r��Ϻ���/�ey� ��2ǜpX��0�.�!�n�y;�|F,\A��)��>���4F�x%%�"��>�&�L=z:�w���JM1�n����m�~�����M����-ⲁ�K+���1�++<"W�	�Φ�qA�O��Lb���ZY1a7�]��@ ��ɤ�4�pɵvrR���M���WCQ���H�hz|���>� ��%n<����+��:y���7ee�^�ZS��Є�Up�,��3֗ QI�I	�1�>t�>A�������>�s��n�5�v��-����@3wQ�p�g�����+�^f�Ѣ�d)v��QC�S��-D�O��I�0ON��-���_*J^V^}5i�N�ɩ�z��s� ��:@`�:�?)o��+�Q��� ��i3^�e+_`�"��6T徯����D/:�7A�������(�{��#� 4�������_mm4��Ʃ�6�,j��D,���W���(�� �"�n��6r�P9���_*�/����f�)s����m(���aM�\�M����E�(�A��֎����L�`���SD	�航����.�h�Ƥ����e%�Fa;N�oP��0�_�&&��\�&��1��8�[�@3�nF�{#j܀G���s|lj����?�(߭:�q��ыF�ef�Ч�@i-�� ��N\ϯ#��}}����EOHT��;��0��b��ܜ�xF��bH��T3&y���՜+�1Q�ΒrT�ؠؼ�B���s���xc0���xYV�+��bO�Z҇��X���P%S�`�P�?�B����mBڞ�T������xX���y�׿t2:�_WFM�l�'w���o�D���H�/��#��qv����N}�OT}Qu�T)�,!2��]�(�I��0g�>�ݳ�g��Oy��xٹFz�B3a��{�:Γ�g�V#"W����w'��"Oo�$�5���Nf��1�Ӿ�T&'��]c��m�Ej���6��p2g��hFA��d�����l	��0W�k,3Q"t�~��Z�+SX� �~�-�#� ��<����r�F��+�\�����|���3K\܊�
�g�RE�X,�2I�$y;��]�zS���朋�.�v�i�G�9�_Ŝbf��y��Y���u���3�CܯE8�����V�TV��-gj����S�fc��T��9~��~��G"4ΥK?�8��@ �y��R�6�]���g�^~^�G��~��9���qTl�{��C�!5�̏�v�*dR,��<�H=�w����{̗�0$>� (�T�;�S�般:���Ws^w��S<��ү`���HF ߟ�>���V����l�]����\��@�â�}#����\��5�Z���5�~���'¯�&��se���J�b�ܬ��,������U���) Si�杘��Q�ms	�/xq�^�&b�;y;uz�]b����zGt���@i��\�^?W��ERt��㩂�7t����מ�鎋k䕴�V���VF�Հ�L��^�I�U� {�1�Je��ˍj��=_:��\`�yN�o�x��W�fSo*�,�����4��T��&lU�M�W��D��x} ^��,v�����~x�u^���M���fU�$�)0�����h�Q��7���jă�z�����0��* 䗗�@�Й5r���*�Q�éW�Lh���4��&S�i��ǫ�)��o�!�;�'�1z��$���=�)v"��V�J�����z�V7_@gk5�+�Ƨ�Ϭ5��71"���\G�_u$'��b��]t��8&8˒�<�Ͳ�KJ{c ����"�Y�_0�D�)�n]A���+�&�+,6�����v���+i�\���8���'~zGAdǥ_�+
��C  ������a�����8�w���@"!�|�Շ/�>�����


h�x����1��@`�����K��n��Ӧ�#�M�3<K�^s����)4k��������<<����~��MA�oO���&މ�'w��۶崂��_�%�#<j��"טr3-J�C��x�"_���(�r��n��]�T��(B�)�K�_1��[����- ]z�+�;S�<����T��x�?@~����6�%�GF}�����X��|+h�yE����.[!P�YNy�!wCh">���9��@��]E�CK��E�m�'=$t� n�ӡ�pr��������x/x�>}�?����H@�J%��ٖb�����I�uDY�������o�T1��dZQQ��}����ζ֍�&�M�����z@��ژ��
c�l�����L�!H�n��R��#殞8O�]��-�l�̘���٧C��Y�1i`h���-h��s�2��UZ}@������U�v�K��Z9��څ-j��6JN�[���o�	����*�-K_��~��Q6NR*��"��o٨!��ڪ|��K�rO_������F��;Yj���y3�?�ƸH��@�2�'N����6�Q:����^�����x�J�f0��C�r�n��l�l	
�������[�Ҋ�X>#�8���F���s	�mN�w�,�!�Ζ�}!e�1����A��&���:�y���L�m�_T����N��|3��g��h2�߻]�9�~����G�z���t��$��(�x:-��&G��L�7����Yj��
g�򞉪���[��]���SU^�Eҗ���Z�ۃ�h��&C5�2͢vk��R��_�K�TB|ַ3P7�D��!��;O<��q}9(��r3@�::mE@���^��6p���$|jc6)ca�h9���E��+�Q�F#��]��v�/��<�Y����A�������c�\��~O���j��P	��Wy�js�vǲ�^�±����wdŷ,t��Q�ם�;�/e�(7��m�6!1d9��\�+���p�d^uǕճK��wH�F��ϕMj�'�D���hhp�ڥƩE/JK�tl�CEj��#]�i2]������v�N�+��N]�6=ӛr戓�V#���pXFrϰ��}P�sg�~�'牎��<�2�»F_)�Ϸy�~'Lن��4U��D�A8��E{���q��<�_�O���lmm'y��_m��^\^�-68ؤhB�LT���A������㮴��̠���!>�����]�� k���Q�-l���ypc�I��;�ni�:����X��Ĺ]K��I��&C'��#���I�<Ж�פ˴����Yn�C#c�����,W�rΊ	w�I��3T�r>���/Ge��kKo�=T�m
���5��b�ju\G㚻`DP���y^�g<�����%6���w'j��0Oq��V���Ĵ�|��g�W�t�$�t.���_�#��0�Q��I ))ys�ґ�����F=Y��K`0�尼�E���v�}qW�fa���b��hC��3�9�÷��m[�Ѕ��VT@yj�d?�!x�nQJE���$����nװv��q��7ݷ�.a_��+l�g�7�>�B�{����y�K��ܿyy=5����6F��aۑ���\�y+�笗.K>�o;K�˪>��R�}l/#`2k��Eo&�݉<D����Jk[kc�'])�u/���q띇����7�%��N�[N3�ֲV���M\n`f��5(���+������𚲼����gN�O�Ua��A����.8P(/W�P�X����	�zq}m]���tD�fݦaL9�5�Ay��i`m;`eT����\������3 p!5!�������Y�S# y���U|��A��:^ a%�dn����}�{�� �/�A2W�
R��L�A?Y�'������No �����'� ���aB��i�;I�<R'��q��]Ҳ�EM�)ݼ���;�&�|��}��z4l�)���p:.���q���`���|�"���b�$�%L����!{��\SS��UU�yy�i�ܻ�Vv����\P�C`o��a�DEP|b��e�����w?䑼	�5��֞`3a��:N`��x�u�H�.cGw󇣂ȣ�n���L5��G��W� ș�b��9�pj�p�#�K⢩`�:��<��$ݵoCo��-�,�8'�9��T�D���G����Y��8oweV��9�W�]���䁜��P���+{1�Rg�n���[�U�V�����R�JH�����J|rrrݰkU�ݝ��R3����:����Ȟb�$K)p�1+'3��bh������0�eK�Euyl�x�%鰬 �����[�>�u��_b�v@?<�1f��dH�.̢RK����b�h���	ͤm��Vg���f��1�h����'h	�J5,����"Oĺ�8ҡ���1xSڃ���F���j��W�
2����L�\�'��Q��������ϕ��y"�#���g���l%�۽��W�ڴF�48~V�^;�Eհ�Q^K�G�4��(*/�+�,����Bgm�J,Z����+/�.v�%u�sM�n/�먺��X?�
:yȩ�;9p��@�	U����\˅u
s��1��CܭO<)�ү�����l���`��I"��J���&�G��zG��{���0�q�R������	s
�t�E,��u2rř��~��'.�^���3eaf=��0*��V��]��{��Q�%�#B,��V,����Z�v�gG�a�x�m>_������i�޴6F�rpw�����]���/�x�xpL�&ùF���Ař���oK���A�2M��[՗Lh���A���3�4$�\H%��1"�k</�L]��HZ+t�����y�[<���@�zYD\���8���� f+Q7o�:�<h��X�n�6f�#�V2R�sנ%?o�9�gּ���b!�
 V۠Ôk�VࢻFz��nY͏��_"O�p��f����< ċ�@��O��E�|�����U��1c�Oa�?'/mh�.`s_�\��Ee,�w�g����z����w|�fB���i���~��ax����R>��2&MQ��ƕ���+�ֻ�Rrrg7H�F���׎�y��E���lA��e�֜��2����Zq�#Da�(39j��[|;�S��l��P�(��w�Ǚ��R?]hՙԼ4r3�Kd�^�+KD�t�������r{�!��8����,���Hnj�ғ��h����� 3��Lŉ�w��H�3��~�`k��K��v߳��[���,{DZ/�$'ȴ��N7��}^�#++�H��E�~��#�K^�3���$�k�ʐ_�!��]�;<��L��W������;�&Х���Q"~&(Á�V%2���P�(�ϼ=�	s��n�>`�}�+����d~�M�䉌�.^�&N�T�a��l/�4U`-z�Êz�i��ZGy?�[���v��B.e�V�k��Gs����B9MpMF�l���	��{΍F+���Z���j���E��5��i����7��v������v�)���#a0�U�D飞�q5�
�K�T���$�`�U%5���}���j;�����i��T���6T��-�p��/A|������ǩ��-���=�jk�j򹏖[�ү:
b8�˓�
p��"�5q��|�^L���ȒLx����5��Cl��͊Q͑W�@CR�o�4#�4��_���
@r��* j��]���I@�o��C S}s�>zP�nYګ51Y<}(�_g��W[���I����'�����m+(C�㳟Nv�>��c�t�?e�7�(����{E`��&$88X���G��������eg�����O���[�w�,�B?1l�i�G���k�Je���h��w�`>	���Q�G�\�c�~#��9A�C���nf�@�0�\� ��g ɬC��J�#�ט,��8�@�Ӷ���q�i.eΫ�YVZ�������l��zɷDkԊY'&}!a�c�MCk�x�ƈf�"�x����-��n�yDp�ގ6�Pe����Qk��l�� �y�&��� bi�´$߶������?�`�7�\/((h�a3?Yi���Uy���)2�$P�}E:��=�eR/X#���N�4yo`}҂�\�{�@�;��@�tݩ�b�6�^�0���)⁇
{���29�&�ߧ:�F#(�Zp�vF�;5�h:*�Z��Cdmדm����W����r�G�85��ſ�G�%g�]�njڕ/q�l��,���E���� 4��1�8�:�ܖ���@
T3�,�qGR��ppp�^�z5؈��fy�y�.ԜY�1��{y�<��גr�d�S��3�X\j��hs�I��I�%`�ώu�0��}"Z`��aǀ�+}�ž:�����CǭtҮ���z����G`9j=�}��4��%!xZ�����Z�e�@v�+�s��G�i��JX₇f�LbEz����U�<ә^ON����7,�X�g��b7n� cD<Qd+ RW�%`[�M��1�kt�[�h���U��\mYƊ�yK��ˊ�bRy`�U��ܨ��%_�Lj�/E�����5Gr��ǈq1_v ��Y'k��Ϣ��K���ٕ�P�ﯭ���k
�R֧_Ϻ�Go�U�HIt�������N4f~�5Ln1��C�d�.C���:�GC�֧��w��#a�Y3�E��oM��(��Tʦ,���Leg�*]j(=�H� �N��^�o2�� JH�}[�ކ�lO�H8!����Lk{�®ɑߖ���U8U2tg�X���Ga�6���L��}�Y@��?N���ד�K�s!�vܰva˽t�9����ZcccWМ�Z�+��RӾE��, �NL|ÞT�����F ��ys֟<�S������K���o���L�- ���d������FKr����;8����{� ���m:��tz��{<!����=�]��L�e?�&�'��ʦ�OuW�ڍ$���:�E�쬰1O���B�����9z��Ծ�����ᝡ�� T��Axt��z;CØb�����_�\����6#�k��Y�������n�9<I����D��	���W;P���7&t�<����u��ta����-����Js��9Mk��GtIF�7$��~���h�B���Ǆz���-�M�e��~L����G�9E���,�b$��oN�~�@�)�ad� ɸ�.���[����T65��87� ��9[?@�TvL�>��nq38������h_,�����yKG����y��q"�a�Z��JW���G-�$�".B<�x���"��(�q�j�㗭��O��<��RL�;�;�.��lR4�ɥL�D6��5ioj��^V7(ћ����D�zO�3=����ui�-�7"L��}���s<ĳ���V��-,�����d���JJ ��}S����%cN���[��#�E��d��xd:��l��L�hs���oZ�a� Sߕ_���_N��_��n�!�Q#�D_���i�8�)��zޢ�r8�p7����4��o"P4����^��Ru�&뿹9R�ٴ�O�r4���-		�f�����k3,����l�!Z���(�)����w�w�?$��ɉ0������Q��b
)��?P)ּU�KJ�Cۗ4�0N�&����>=o��?�`��l�w��d�?�u��s����S�X��E�c�+R�%R/�R�7Z�R:��˫�'�����K�pk���Y��tU��C
i�
{! ���+ާ�ermpK�����E�����
GY9(HU�����2����+��t<�.��sɞ/ԟ�.g�����������9���"Nz�	�S�M��
�[��jA,�b��Ud-KR�V�q�y�̎)�n��`�U$x~�p^�\�=�?	���_ iFD(���2���{���#1}�k�~����m���s2V���c;U:us�P���B'Ɇ�@0���Ds�G7r�$h�8��%x���p�fW�E�R/�Rꜞ���+���i� �c��j*���h�I��a��ᚿ��I(1�3�%^m5��4%w�wt%��/�(�j��X�(x�ۤZ�?iM�/X;8�e�����J�I�I�**�3�ړ�|����S���z���g�l�N�fnO�InPQU�GZ�l�#YX� �4�!u�C@� �� � p����),FĄ��
2�暺���g������j�"}⋳c\2���s�뼻��Q��9ћ�7�7���0�J�Hơ���4�>��q��#n�9�*��+��B��!�'����[\F��q�m� �o}7(�J,[aC�_�ՙh��S���l˦ꪅ�,�	��$��,&g��j����[�:O���^t�.}���M�M��հ8�%b�7/ۯ����^�u,r� ���X�8|r�	�pߑD�7��p�Y�+F-ᅏ'y�ϭ)@���5��xNB�ۮ�R�˂D��E|���}�F�!?�jG n:ռt2���CkV����KM�N���x�,Q�y ,f `��:�v+$����.��uz�^ۀ��b���*�
����E��!}��/���b�觺@�h�͈�7	X�d0��w	A����}vT�IE�UR�"ؓ�	�#)M7�h��>s�Ya<���]�w0wi�fp�.�fׂ��?�ym���o׌��=e���t��'U���Յ��n���2�D��������M�eO�X.'�m��'�H�nqG�t�0�����վ<��I�f;#i6)k����s?�	H������|����WdA��1)n�h�v��X�N1�|������TTqޞЅp$��������T�B?i.q�""�?*�s���!� ���`lM�M�}�7:w2��h�ˤ�&����s����C�;���I�@��c��A�_ʖ6U)��rE�5�l��!ݎGB���P�����R���?l�AS	���M5E
�V�fң9�A�G� ~f������o�il�	��ʬ`�sf�w+ �w�F�F�w~�B���E��4��~(���<�,�_$���Q�#@.s�9�p��TUU�o��M�V��&��D��i�9��hLf�x��r���N�>��K9���_��߿HĹwGA�]=��F��R��?K�{��Wy!%3�����Sf�C*��vwzu0�S��KG��Xh)5O^j]	7%�q��j���C��A�X�H���x�߮u�o3K�z.�=h'�����B��POe �80�S(PE��d\�E����
2U��3s��w[�E����hN"�f?Ju�jn�XTvv&�gސ���P�Zn��S���g���I���=g��;�������eNo�?�6Nx������6g��/��4�K���pU����A��~G�"�9�#��e�1�Q}�����$>���o&��M�>��O��K���n�gw̷'�1��-Z���@�r	˩�:w�g��nt`�hv�^�Q�\2� M�!zfV�\�J)YK��*���FH����_W��c�5y���Ǻ�O�k��o��0����}�|la��4r��NtLG?m	IT2��ܻ̽7s��kt8]�1��P@YlC����h,I�ƻ���z�3��>z)Xo�n&:u�;"9�����������iGN���D��G�J���
C�͜pe��i�a9��D2`��+8�k���e�ECV�W=�TѓXՁ!�����?ֽi[ZZ&y,�?�gKz��9�U�)�3��?���3����b���֭��{�lzr o��À�ȵ��Er��B�*oء<�0���~����b�Ԓsq6鲛�We0����f�"J.�	.έZ�*�[V㠛�8,�t����n�V�ρ���`\��E��>��ֳ�FJ�}ܨ����}R	���݂ՏZ$1&Wx&�D3�G�ٚ�O�}/�u�o~�3�％�,��.D��: �e9�g���&X��s�&��WyϬ��t��4L�q��޿�ߵ"G���v�<W���.u}/�������������oT#{��M�z5P:�n|'	"9����?���8F�8�����tv"�ZM3��\������a������%	u�R�6)-��2�[^X�a�f������A�:s,��S�[��lG����k���Dq;��,xRSyf�Q�����C�n��p���?��H�):��<9� &�I�J�1��@���Y©F�"��H��}��Π��Q���B��]q�Ӑȕ�XJ%�Ӽ�T���ت��=-��EȔxd8>x��|뗦ο�qބ/Lu�pr_w��utG̻��пO�q7m��%k�فxTr~~���}������P���q&־[R�g�>m��ێ���_��-tZ��WԢ�LP�ԗ����h6_�����^j�k'S����s�"��<k/�/l�M��*��l�.0Uj>�0ѳ^���:���
i�AÄ���(�nY��]�'x{P zȻ�|t�ΰ�#�5b-f>DF�e���ʑb�eaq�y+���u{6��W�U�N�S�{x���eJ������ĨKJF-�:���r�N
�I�U;(����Vm����"H�U�̲J�ߍ��U��z��H�*�½����h�.��#Ű�^�����V�|�N۔�/�R_��yEY�h=���P��;nG���N�����E���Kf�_\\_�&����~"f��-#i���=�}||`�Hx�����,xlL��n*��b�}h?i��ť��J9w~N�y~2-x����m=��������K&r�a�m�3\��E����!�fFlt��T$���!�c����l�$s"����T,.2v��T�+,��Bt�l����Uخ�*�yA�S����6h�!݆c6:��N����T�8~qR���s�X /�ֿ^'#�8F1�b�]�B%���sጉ5p��Ǜ-�������W2x����l�	�Bf�&w���M+����r����f�'Ϳ��Y�<���Z�/������y�=\mއ��:3��C-,�k{��0�dy�&ؽ�W�l��M��dXu�?s�|UY+�~�F�pA~CX^d�d��?�i|�q2ƒ�K�ڰ�0��pMScC?{I)�a�ӵ�T� ��m�x��O��gϨ����y4�+-ⒻL]�t�#�f��7�k��w^��Z|
�Z�e�ծ=j�c�a>Ԏ9�錡� n�����:Nen.�4ĞP�%p~�e�Ap��rq�nY���C}�m���;o�Aź��tǙA�Dv.�����D�\�^R������z!�`2�M�tL��q�,���:����䧏?a�Nnd��V�w��
���/ �;��J�z��I���(�鉏&����{�)bB�5�����2�֑�6p�oS�4�H@�y�
�B��L���yOu�����
pjո�![Z��7�\�T�c��h1�ؔ�e:&LYj��dp� c�i��G�6�qMn�-�V��!��;�@LĠ���t��gC �Q���Џ�dl5�����N�E�Y[6�fX��3|��,�W/�[�y�W�����0{�æ�?f��T���������A���� �E�+�r\�j�U)���Лɔ�w�
��S<]�M�جM��t�{
s5_��b�VW �݉,ǳ���*�@ "���\�� ���	��FF5k�q{�p)th���>���&���p%l2V'�Z�9/��>���p���Gڣo��W2��3�2|����us�j�"m<;��⭄��.ڟ�`0Ե�uF��E>O���YK0�M�u��a�-,���c�^^+^	�C��w}z���q���gk�`�X�|��]�K{&|]�F�$%0�S��t�+�����[��rZ^)�������ۥ���'+m7w���1�>�εV_��S���>��z��;�7v_�g�����V�m&Hg)d_�3��wi�==�1����������;[�"��k?)�j���Ύ�ׄ7ՙ(Ů�y��/�RBa1��]��6f���XJɨ���S��h59D�Jʨq䃌*R�VzH ��-��Ր��iJ�tr�s��:˲��r���(D~�>�e�I���Jq�]��l�_�����6_ z{㜃T��K"��{��5�W=�7�nP$T�sB"���U�l�%^��(�2�hTv����c�%7��[�����lEbh�B���XV�K@����[''ޙ
�9��%�����5)�r#�Q!avɗ[�/Õ��;�p�W�&��O>���8�l|%�wk�.��[�V��}8�ɉ��h�?ο�n̝p!��Y�9��8�­�^�F��#�`��ϪDI�����v��P�#��J����G8�_�-A�K����q�@X�D�����f��,��<��H^��gwj5��\&�uC�y�8�Ȟ�yB���\�ׁ�`Y�+���,S�v�{�:�FZYE��e��Ï�\DH�<:����d|��7'�?�����ʂ`]ht��3�̽M�ӝ�Jd{�1i���X������;���^3���q�Iݼ��-VoJ���ʺYڕ�	XG#��0jB��{J�`@/�f�.����4t��M:�R�ŃqT���i�EI���r�ܾ���6`j�D+@º�b9븶�x�4�0�i
p�5�bv���Q#6r�Uh�Bx���O:lp0�m�-XS~Ȟ���ʹ�/�s0g�&��~H�a���Gq�zh3<��X��N��^�̯]���k����H�O#,{�\b�dہ|�S�@������j����~�����W�_�\��9r���v�=����������94�i72��/]���i;����t��r��w��M��R� �E|`�V(���8�x	Ε�f!d��VQ�f����a6�d�)7%�\j[���TH{Z����7}`��k�k��p���]�Y�w�6��������0����=*���o
lC�T���'��"\Kw��O��}�S{+_Q�L���˲>����� 1Wm0���h�I�9]��K�zv�
3��3
�Tx����\�5w]V�:}�Q����[�߹���="j��v��)�8ߖ�W\���X
p>p��h�0�ZG����x]��-)1.++������:��F[[[ ���=��y���Vy׵����O�v?�@R=�Pu�;*���5S��`��B�B�/V��O��QuM��ݰaʎ�۫��Y5Ĉ^(0�hm�<&6Q쟎_�z��G�yb�.�-H]?��wZZd���ű߹��@�=�zu�T��HCҕ!o��80�����4�Ѫy�*dDk)���_�\��f��GՎ R��R�}�kY����`�s�=�3K�(;�;�IEs�x��Ip�l�޲M�����2�̯q�X��'*��22�Hy��*����� '�[P�3F���4�a�.�������G���Vђ 2�6�L�4I_�1�g������w�x����]/G��1�_M�lD����A�!X.S�4i�$���o�lÓ(���~
ϩ�n�!�T��n&�C;�3&��8�q�7c��J'J��f�C���*���'�(�r(��֙h�����l�T��Y��a�,�m�jm�������=�K���-{L���3�r�^�ʀ��+��M1n��>fc�?�F�m�?�v�zHҦ�:G�H��G5��w%�JFOV���&��e{�$:�NbU����w?i��h�������0Zd����q;6� ��IE��բ�SC~4��X����Ug�@�.]�&r���):��@h��|\���r�FQ� ��ۀA:;��
	
o����m&i�G��5��Y;K8��W c6����'
:{�jd*�+�.�H���6'�h�,�p����z�|���R�@�7tc��P6o�qGA���U�A$��!}�J~�
��Z_��ob�Z�C�߮Rc�<Ē9s)AWs���Gr��ީ7��ZO��'���,��þ���̓[�J�sH��z����=7���^���V�k,|,�7xv �����!���D���T�
�?�VI ��m�V{_��yu*PT'���lI�B��>�	��v�/7c�vK�"���P;W�6֠������cY+++[���K�K.�,�f��"�-�Y���1Y��6��P��,N��<X]U�^�&(V�C��O��e�u��Vz��ă6���&f�Ku���_�m1��.�2�CEt[r����T�A�H\�Dڿ9�����?0�+k�cP����_D��� �H�" �!�!"]ҹ"���"-% ��� ��H	,]K�ұ������=�[�qv�3󝙏�sw-mW�=��|jG�O���V���¿��ZN�ۦ�=�=��[�۬��!K���	�������t<A�o���XX�;"wKn 1�7�	]�k�=2%w?�P	z[�6/�-[�A�e�l������'x(�	W�S1�~���~Ǒ��_���	��-Dh#�I=�,P��ڝ���M ���K��#��b�����sB΅)P��5�����E�1 �%���<n!��2�,�q�c9��W	zV$k+=D�ݨ���E���-6��'״�y_-7��ꏐ��fu}qu:����1=`c�U[��8�Rַ���֩�ǒ��s��.���u�-��X��D�}�7�kq{��4�^/& �R:}�
���U8�?�*�dE>�������!WϞ��� uTT��X��nA!�s��);���\=Ǥ*~�T�����;�I~`I�?>�]/_�!@��~?(vzl��`t��0�� ����d�f��er����w�36�-��A�����'�����G��91��D��!a��DX�S�xZ�vu{V�VZ4�n�|�{�1�K�[�7#�#!�
-R��P�j��ɾW%@A�c�J�W�п���@ѻ<�%�%���G�R�O~��o�+�نw���?\�)&]�x���Er�8��TF�)�2j���kk��0	Ǔ@ Ժ 5BJ�[�ѿ�����toUh������u�?y�lQ�b�!��es��q��]bo.p�xA��;f�Qj�Nɥ���i�z�)��R��1,�"d��؉3/�_���#�����!߸q[z�6Um0�m<�Z�2�?f_D[�߈�+���_�d>U�6��	��� Z��Y{¨n����9.	�����o��t�~�C�q���i�W�ITǻ&��8�uDA��e�?�,|�?�4j/��3v]����t�,K���D�ReX��a�����Oнkm�SnsK)y���J�T,$�Fٶ4�ԝ��g��5�܈�'��oؗ��Թ��H�
)�,}��S� 𥆮iD��2)������?anm&`� )�8���4�����ᘜITG�Ɯ�q�O,��B�����"ވ���e��S�[*�R[��GٰN�OgO�F�X�G�iFP�۪�z�c>�V��o��D���&LV����
-n���L���ֱa�lKa�2
{��%�����NMX}q�?��f 1��O��f�hV �ɧu�%�'餹2ǃ5���MıCؽk	=2hX8�G�j7�1��k�(|iF=Z�7ĥ�w�������Ės^E~���!��h��X�� ��q�ښ^�^��� oSv�r8���r�i�F�jKH!�t}�]gt������13䵃��n�񃛋�xz ����p�@ą����k$t�����v6������/�g�j�W�����+ou���@!�GK𛼺2��Q�>[�i�%�)�,jN7x�:���������!�>��໮�Eѕ7X8�T�%�\w�1o�ϸ�=����e|_'J:�j��+M��6?c��#��8�֭g���;�aC5�m]�� y_����C�%����ɞLt�Wz�tB��s�ns�|g�W�;f�2~�jS��o�3�F�3�-p���>����a����ك�T��.�N�) _��w΅��Dޕi�����m�*}?i8/+cY�ZʡX�qt�%�؉�/~����� ��������)r�ga���A̳�y-b�������&r��u�+�`_y���w�h�hp�[咽<L~�w4BK+s$��4�"Y]�ݱ�Գ�����a��/��Xpvљ�:+ٖ��Ðǌ�°�V�[��"�f�"ӛ [�ٲ�����>߲���?þ�X�?u�F�/��i�^���ȠԮ1����T6_$Lu����)�[���x/,w�&��tU�kr�[B�NR��i)�h����zW34^�s�[{�ġ�T�y���k��?� ��e�����jA������z�����o�b�Lt�6��C������j��S��:�g�V!�@�5/Ft��ܝje6/��!Q\�=��a'���h�#6]����"^7ƛ''1n��5�V�0��y��u�r�N,�Hv��mP�H�Rt4�.���&�`9ۛ_�*Û"�پ��c~��0ؑ)��|�2�DD�U���B@D[����E�y�M��R�-	�=��ÄǓ��6�TV��r
xT�7���2h�x������;!�<r_�e�7�CL�|��'��H虈K4V̏�E��wW�]M��eS���n������r��؋�so�f������5�H$�æ�#YMsK�CS���Ck�`J'�y�_荊��o#��T��z`]�lj!��Թf��1�W��9Y��&��l��,�
��$���((��q����y��
"��u��zH�[ޠW,#t��0!�D���c:\�P-��-UԬg�����ej)�o�Ι~�ER���s����oʢ�������%�6kf�ڣC
���1#r񻭈ms�����)[�[Ǫp���CK�n�[@�k����x�h��T�p��S�Vя+�B}\~�ѕq�<�v�3���Hk��������p���<d�d��[�~$�V(-��Ȟ
�l���{��%8?����Σ��W�pd��K��:��\��:�Hom�߯��1Y}�.S�҉�?�?%-;fg�8Hf^wf���Q&4iٮ�s)ϴ���Vyo��r%��Ā�ILǬ�{٫܊@��������W�&��|��Z�R������טQ���+�0�4�����[7;vg7�3>�1�� h���j�m=��1�5�R��h��}Q�&�a� � ��D$�j�w��� ͨt��L��W@�Xؾ|�����1���W�� '9�����tc;ZHX�kz��X~��',M	裳�H| Ј��M\;����lV���N��,E&քw.1��r�ҫi8�Cr�95q4V�����V��Zn�3g�k�iV�FL��q������˽:��>����4*M��o�����E-3���hR鹖��5&�fD�0CG~d��֣��"_��[�&�E�w֒�Y��SN"��|�!��;)���y��D�b蒡U^�	 n�R�5��Pc�@��:^��c�ZQ웣n��Yէ�+��J��+ɓǎ�Z1SK������1���\>���5o�7��?-<�\�'�pmU���᭦*z��ΙE4[�c伩��E�����ak[��O�m�/'��tXǪ蹭zY+�}Pȋ�q$oe#����^Ѩx)w}Ѡ�ӂb�e��H "��i�ɋi��T��KO�Z�'��q����G�5VY6<��K֌�a��ͳ��iՒ�C�^�ȱ��w�c	��9p���S~�~���l,�He�wf#����b��'���+eR�j�S ��L7`;��ųU1��z�*�O��'J�a_D���K�	I`v�0wDG����H������pSw:�!mʦN�#�o"UÎ�EV��;����KOJHטu�^2����0/��t�>k}U6���(,��/T�l����W�Iq��~X�ϗZ>�N:>1�h��1M��g����&.�jA"I�T����(����W��y�.�e�Y�-�Mx9�iDt��%H7+#* .Ir3q4 �� �̲0|}�#��A�L��y�m�MG�Y���Ij���p���>!�F�V��r�[�(;M��]� �	4@�[c��⦧��)l4Ĳ@CR.X���qRׁ
 �4I��RFu#��fL7��|gwML�v6�h\���f���W��&�6�x2ޭT.N��\(���Az���,>"�����K��~���E�����/�T��������l{�I�	�@��//Ɵ�ހ�c֝������X����1������Xä�L](c���Hu�1�0 ��Q���6�����cx/�C;|�k��yv=�)
���iS�]�~����+�墥��9�J�&x��a�h/$*U�I�>�D7�����P}�x�|8�W��a$���<Q�ٌ��[P�?�G���xC�a&�޾�ɛy��� E��5�=}G[�Ւ�"�u�^�=}!y�?Yq{��)�̅�~t��1��4���Jr5�;?�f��a?t��ܐhd�w5�����!���Y0n+OЖ`k���NCմ�3s4$�A|BL/Z?�xYj�;�Ր�W]hc*q*ݳ� ��C(�����m��0ʵ�-w��/������SE)�\/o�2�$�q�S�ֵ���O�����F��^+l�Y��*�6 '���#1[#?����5����U
W�ߜ)K��)#��^_�Dа�kJwO��
ҭ��-z�7V*�����3�
֠�H��#o���L���n�@��l�����Z��A>_s��>��9��!�a9�c�ޯ����A�I �]CG�%�!.�5���	BoB;�R�c�g-瓪���獪�nD�H�Ǒ�� ��X�6��,���*O:���ps嵙����5�~jN���z��;�O#:��B�=�|�g{��P�.��%���{4o��T��za?r��$H��jCs֊�G�=���Ā�'�V>��E8�P�q+8y�:��@�뵞#�X�^�~��1�m��4)���J��q�� ��M����S�^�,�döe#P�8g�dO~�	�F��G۔5��\I|6�e�� �f��hzL��2t�wja�׹ҳ��n��[PL�$@�d�����W����e��ng��|��7w��Ҿ�y+�����h�=��AN4����C�;;;�:֢i�gg��4p<B�M/1>j�Ư*�9�p�6y�Q$��-�\Qʬ�bl������浌��2oIk�CU��$费��6y�^�H��P���=Nm/�cS���<i~�ν����,��2�'��%lm����j��E�ל���m��+�9��'���v�D�<wN��W�M�U2y���O� ��?[��*%��ӭ�����^`���;��x�/3ц
�3�eEy�o�500�ɓy��!�r5��/p��NV���4�z	U�xߚ���w4p&8ۡ/��d�*�v�C������>�l�ݚQ�^��y�N����Tr|;??_�P���?�s]�P������R��l$������kX���>al��_K�W]��`�/����h.7���S�8��\�F��!�}0��2�i>oC��1���Fs��w��u)��*��&)>o�П�׃]x�����?
��v�x���!,�AUq��m�ZQ~��L��g��\'h�b�e�/	k:�G����[�'�ƈK�����)�7�{�w��&6�3�4��M�?A�'#"y��'$lt���
-�fꚌ�.�ӊ��� �S���9�^4� o��[���؁��0��#�ڒ��{�!n�R�$��1�)�)l���!7-�69IqZ��:�VVR/��������)
J+~9G����9[e�4OI��s����l�Ih�tP���RF桎�ϔ\�g���^`����d�Cȃ��bmnޮ��Gn��qk2��D�Rh!�fZU���-|2�o@�q��t/I�Z]�8��
v��ŭ7P�h�����K�2�W��8S*��7��+*��rS�k�̻�5�'S���f1:�"���d�5z�}�ӫN����$�W{��ƼK�J�s̮�o���b�eBmK9�~HR�t<�׸/�NŎ=20��f�FqAD����X����=�<�T�]���/Y������{�q[����&&$����4����LƄ-��$�kD99X�^N�?^���R�OlR%�u���3�J���7��s3+'\J�6�f�n��.$�Ev�Ŀi]3�l+5���Yd�.�򧴷�(˼�C�Q����� ��z�B���8]�Q��0�Q�������6D�I/XC��X�v�_Xg�m�nJ�5Y���+�K��܆FЖ|aE�w֑R�@��*�m�KFx��t�E�:EQn�x�V�=E&�|�B����M��p���o�_���/�Y\��+&�O%21=����bY}�nk#O2���"���<ޯؾ�0?_�4W>��2��0p_�}��0������ā�U,��o����1�r)�a��s	�8���D�c���F�n_��ژ���
�✪i�%Ne��u���K�0Q���ʤ�\_#�'q�u$�c'�֤��&ӥ~&����v��0�*�����n��H9���g�:�g��pv�[e�O^�Ps���޹��OH��k��v'����߼(A����~Z��z�ş���6�����ʳ!�0wn�b	Km�ڑ�k�G������.|Q��qG���׎u�?��\�	�-aa(UF,yP3_��-ď��>3NhI�f�<��|_Q/������Ў�S^�W�ƆX��!9�=������K�C��h
�c�Tʸ�/+
ό���;Q����Ճ�MQ@���ۍac�s�ؐw̘�"σ(�#�d���\�Z��쒺y�?L��kG�_Zd�&�N6�pt��R����W奋.�扷��<�
:,k��(�����\{���N��ެ�|wݰt
�YȯSh�Å�~t�6�aybA�.2��G��<M�.WC\	[��v��dN�K%�#�p8j���yc5�<�÷��e�����!�3��*����ӕYK��Ye�rX�^�懻$��'d\���._���x�f�P|.+4� ��j7�̍ʮ�������n���q�Bv~TA+.f��?&��B��h����������
c�>)(˕�I-l���8&�a��'ς��6�g�J�*x�<�(�������4�~�3�o��^�D��d������<��G��1i����p,�������I֏S����	G���k7���K�����t�wA�v�����ʇ��G��Їųj�&��i���	���v��@OB��3+�[��'��9VG�Oc%�j���A8�8����~�F|?�<���
?��$�(���<�"��:����3�(ݖ�S\�!�T����݈�P&V��^�Mw7�8>��"����io�n�H��k�]�����Sܚ">kf�pdGKv-�'���n��-��]�w�M�21��M=~�HF`�S���!�Iz�!׫�{F������0��0���'[���aG�7�y���ӳ��k˕�K�OŃe<Y����[x���Q�1�kY�f��N�zn��4��=X�0�S�F�)��g������I��uD����hݥ���Y��b��=WI�B��oJ�ZL�:B�1�(l�C�O�3�������JRDw�F�7o�|@��B�2� '���1Zb"򽲿)�A:���9-��ەK��=h������+˒9��P`��o�����8��]?O�p��H��o�����F;GԆ���2Y����ݣLtNoE�Xa�N^SBF�?��G�U#��3��X����߹�b���w饒s��e�˒x�!�yv9z�7Fm5����Њ��Y��4���Z��ȷ�0�_���*2	tU����(�ڹ
[�^IrB	�v�����La���.���O2�j��5Dկ�d7�n�z���(�L@O�O�_Z"�f�㒸���_�QMIS����)�V�͵���o" �����Z	�Q�V�b���[r%Ha�|n��{��;.�U�9׮�i�A���J�4"��/��G���p���vhBXʃEzr->�P�Ah�y�^�)��Ũ�Wu�P���bE�ҕ=����U���X��80qߺ]�W�e�5����-�5�ţ�hDX2]���$�=�o���E���(�>�,|��W�A;��:+;a�V@���8:ʧ�<�Q��A����F{K❗u^!�H� y���������b���q�1ek&�Q܃���:�MmP�(��HpXGB4؛�ζ�����+�XXLO�'�_���
��{��*�\���I�G��$��\Q�K<5�0t�,�:�/@�ar�C�}��q���37","��T�8����x$����T{;���X��3���E���~�6����n4�b;��r�×�6����ζ��"-�3$K=3��$;�`�:��d�L��U��b� 4����!��rl�O@6#k�/��tz��ǌ��^����b��������Mw>�J����&f�CT1�"�u�s ;�8�tPo�.����!�W�a#1Cd�[^nn����SX���'�\^��~��N�T��?O�������T@m�x �53R���<��K!���fkä����{>�Ψaˮ�h�>���J������΅{¬W���tiS����{撶���d#��E��7��V_��E����ް�X�|b���|����f�lj"��U����]]�U�IF^1h`t�F1���ZM�e!�Ipԟ�k��6B硎�!�@��̧:&�crJ��i8��1��L ���^o�]���r>;�^����%��N�2�b��D��*Sf��m2�_I�؏�����N�ŗ`(*�GI��/X���ׅ�7K�*&�w�]:��he��!<����)��\�d�/iLq�~�I�o�>jc���wx��agyZ,�b�x���{A�p(��xu�d``0_**�[��Y�D��������d����.���_���S�+�@��	x�=q0#�"}+mݘx )��J�BQ�H$�����Bk�D�`�����D����VBgA�mv'x�r��3Br~@����~��f*0jw?q��桢�S�:zx�@h�s<����j��&���� '��c:x6(�ABT�4��)��0�,�Uh�~�V������_��em�KJS��\&A�վ������?�V}2Ƭ�7i����6+]��W��*)�D�JϺwa��׵'�}bh��W�����a�sZ�Qgռ}��mo�Z�|��l�s�3�K"?�@"G��!H�d'�/.c�g-��/�)�[f��#d�EE	`�ܻ�x+r��������<d��Q�;1Nq�_�7P6Lx���\�0�|�+�GO��O�W�`d��Y���@#� LS]�,v�����b�t��9�IZ��|��� �v�J��	����b���ox?@�v��:u[?�men4Pa��wٺ�A�~(h�6ۙ�����N���
�`V��r%2���Lf1]��)y?Gx��}�DPn@�=�5�֣���gh�r�dBO�+��@	��=Dnd���GAJ�gK̆B����3�{rm'y�zz��a��/;�vfv5|,���Yy���m�)R\S���Ǘ(�@�>�GѴ�d./�K���/�$S=�؀����a"b�?D�$��+R��A\�7n�ϱ~��^�q��?W
�Jt�Kd�&T�a't\����X�f���Y��s��odH�+��l��@&�r���x�	�:�E&�#�����f[�:$�4Cw�ܚ�����:�[�J:hM��O%��?H<~ם`���VBk�OX,�Q(Zwd��0����|B,��D_�K�u2��._̶l�<9MMB��{oS���'��7�&�H��܎w�>Y�r����L�__�����/�>C�!��a�?>iY}�F�3�>�w�i�o�-��I1�RC ��,gI���� |��(:x��?��	��=be���y����,AY7:�sغ�x�	�H��ژ��w%w���o���r������v��ں�<*�d�/����s[��|�4^g��`+��Q������S���.���l]yW96	�b�Ǖ����!��}���<�^����|����h~��8����}
pbb��&�ևԑ�9K~���j8�-Ol^g����B��Tq��H��uzn���Q��2A�,qF��`2?�	_�bn]N�c
����N�)�JP��2B&��eE�~N_�¸���g�T� ��d]\[l8-jTe��:d��i���PXGX���|��h��|��G=O��xf������[-�I�/	�4��;z9OW�˽��P/�=��t4	K���'ȲH1ݦ�`H�����h7�����_��VO����_fI,I���]��MK�.����Q"+A$�k+���I�~+�>�#�J+�@R��SyL��jj}�nv4@�c;"�\Ph����'�XeO�e�?<t�w��ߙ�K�MW^
M�ѯ|WZ��|FK#�g��kd��;gҵ�+DYik1[<��&�U<�X�J �2�K�3s""!���X��:�g�ځ��PS`�ؖ�硧F>�>h���5���/��_m�<&�Z��q_��6�`���J�䯡�Oh'��or-�'��y�:P��7#�g�$�'��z ;��'���=Y�*����ܴ�yP{��a�Y����vi^�:$k�x�u&�^\ u��U�d�&O�GvEy20�|Ur��Q�?lЗ���o���G�z�-qS�GL͚+(�$?u�f��܌I4vK/�a6󩈔��{���,N��.]m�l�W��b��$/*5�����؁U��K>4y����΋����[�����f�-9��6>���V6�f��_(��J��,�
�zwh7H̾nhz}���QZ��%��2�[��*\ĿQ�n�@"!c��ⓑ!U��ee �>Z��t���I��7)����V��׽S;��صQ��p�v+ʁ[�3���9�{>��y����M���=[+���V�'Jl?
*��M%̆P����H
K���((�~����<����8��d]�i�4�X�Q��\�A���C'�m
{�(�'W|��j�M������pG�	v<��u>KM	�P��',��oɐD����1�A��	��HT�>Mm9���x�����	陋��1����7���Z�j�8��Ua��?�����h\ 7M8»�����ڱ�X�2@0�=|�u�#:}N��#�n6�Po�:\:.��
\�qX$����L�����݁�q!#ugR��q���9���b��G MȀ�D���n���ੑ���t��z���з�K�y$��T��[��dR^��4��	�{G+�5VT�ku��k�T�ReĆ�!��Բ��ʓ?7���OB{���Ax������wt��a�$������ ��*�ܟ(�ٯW�\�C�!W�����`�ۮ㮻�����2q�1���NQW9k*'�&u�����\CŎ��Z щ��-ߪv9+�����a~��˲�uÞ��+�w�+��S��<�/?�b��g�TJ�H�[xK&�o1����)���x'.��I�\��k�kl� ���h�Ê�Q��V�E��ւ�BdH�h?�M�D-2�nqNƗ�C.��i���� ��:1�g?d�l�M&:������3����^�c�|Pa�mH@9��h_�e���=hO�С=��ى������%����1Ĺy�׌=rT�'p�μcWݵ7Fa�SMZ��םD�|���">�=�0������c	�R�-�T��Kn����S�t)�p�;�f@ Z]=p!�v/�a�)�[`B�{�d�0�w�[��[1R�o��'�'�d<R�+��@�~��iOe:S��a���(���*%1�FJ(ߤ���~����	k%Q5�-C40x��cT�Tx/q�pw�X:��fE���z�?�Օۺ�x�S�a��{�=aT���P�L_B�ˆ�E�an��pP��&1�lW3��&�n���������ߘҟ�%׉�_I���}��FN�z.��j�C@�����������A��:�z�㈃cV%�7��e�F^����^	�ZR�*|к�e�g�WÜ�1��Z�Å��+���& "��y�v�X�(^��:ڝ�*�v�����ʣhʮ�nt!Ao�F@�F��O��S�+Y+��ػi�1��_����V0:̒����'Ԭ��$�'M��`<�_Rd�S�ym��mL�iR�Ud�R%/^~�5�<Wܼx��i,m���C�h^�~��9�&Y��?��!�]� ''�'�XK,&�	�=��$`���^�F�t���=ޭ�wl�L�D�]�t�9��osu|�f'�#�Z�}	�i����l��#��ٙ���Ϣ�B�f����m;q*Y���aM9�*���S5�2�_�W�-3�?���.>����B�E�C�,~�|D�md�ڔmhR!���������")����]jM��L��%@��(
ſ�����d���TӋ
�����UO�8�	2ݘ��;�2^�-eY�J�WJ�U���6G˓�T��S�+`�Gx�J�D��SX�ZدF��
(���}Ʊ'x����9hG����a�v]�؟�I{b�cN:�e�KW΍�r��YlP��V����-���R��x�V���g�m��g�˺. �LC����'�1P��4j��Ax���$��������SӉ�ϕ��;ʾ�%m��:	o�)����B��������u�n�CӝrA�������LH�~ʴ��4}yM�p]��Á�"�tS��1��6@�V���ۯF��W9yh�ʯ�Gz�v_a��3+4�zu#f����q�g�o&�;����:�l�Xz��x�����~{n���C�G���A�|�.��ڭ�/5����R��)��$"]"�fŸ?�y��庮l�);~�g��b�.Q�St=_���&�O�B~��SD*ae�E-��z��G��L"�ymC�Z)��a��Jm�Vy��\b�ѯ?�1�M{�{ϑ�E|�HK�{�"���\�����KH�����]u[�jרC c
�.1C�WX,�K��t�gB�}}��Wo�G�i|�
ݓ�X"�F���hvV��A�(�9 �L�#�\]���G���#OQ��W�}��A�{ �/�8h��p����`���Y��j��h�����c�j�m���p��SA��X�����a�q����l�ʲ��?��Ћv�ҙi>ȬJ�|`Gg�����:`=?�+<=`ѓ{���4KV��3�W:���dL�k��,jR��3i�LQ���Ӹۃ�`_&+�D�w���~�ڿbYW/�4���T��´R�e����- �<�o'��Eo�~\6�j~��K�:����YxBᗜ𩬥�;�l�ҕn�ƚg�-O��d�F���T�ŹXt���\�C�L/��^ltAj����
-gE���J�u�v�����[oL�p��8��Z���;eP�:W�͚����}�0������$I����3>���8��4�y�{P<+?�p|"l;½	D���� E�s|D�u�?��W�lU��x�ט=�K 06d�6�$���E	��O�(]$�V��w����D��板%�j��B����طv��z���痣a����\���p�$�{S�a
�^�f '�j�qX�>-4$6%��K���g��
ؿ����.5����
Y�<p�� f��>j��K)��N�����Zu�鮊L:)�}2\e:����"�Hx�
�Oz�1�K��n�	ZP�g� ����f�v̺�?����L.�}��`�&����©�*����i��$����߰Z*�)e���НZ<��r7���h� v=��g���_�˓�����$
��:nҩ��H�NK��C�9?Q�,��f:��c�,�� ��OBQ�5\GVh}�ܳ��e¤���n�f�F��J��
�@CA#�:j�"g.���m��X�p�#Љ�3� ��F5 ������������%�oG�E�^��&�!!���-���I c����7[���~V��&�Uړ*�JQh�T?�8L���}�kJVK�O�n��gM��%�u��$5f���i�a�9���t���l��wG̣����%�f��5�$�(�����g��f��N�~l�E�.����� ~cfy�52V�y��'1v/���_\�~-����Έ'�#)�)YR�����7��o�j���s�q�(�J� ����$-k>�8��Fak��mR�?p:{A$�A
t/"��a�5U��s�;-ʡ]��S�A��H��zy:w�ې7���&�a~���V}1�|W��Owl%����؟Mvb���b�3�X���A��\���ǔ^��%�<����(?�!�k�r���4��v�뀰b�Qm��ok3}ۺ�s��D4�^?��
\�u�D�^�a��Ѡ��'Q�G>ܤQ$,s���5�����=�=�1��}=o�%3N��oCy�M--쬀B
�G}��0�%�\ω�Yom�ٽ��m#��8�����������%v�ի0���iQ>Rg��J��vQ�X�����+J��UȖ��Z�oUf ɥ�$2�o-�U7�6�4� GZ�q��ʐ�[y�"It���I����
�Z�ͼ�<~�R�=�B���*��y�ɝݷ�w��K��3��,�`5�����0����(�u��J��Zjp�k�!���<W��_���1#Q=����t���˛�'y�l�n�a���7��b�͊f��̈́ٗ���]�/;�����%� ���$�N��V�'y�R<"�������f�'.���8�����ê�FW0Q-�Q�6���G|R�F��u�z�7���!�1�M)���F%}�z�W<bS��W~�G��y{�K
��)��#}�j�s�|�j�""����S*]=y���\%��f�!��B�сiVO�j�>[(� �4?��t�j�����A��� nPR,��HF����~I�O��uF���2��^-��l���^�s�ŧ6��	 �7��o+5�s�x����<7d�D,̶�^ׇ�� �ϔn�JnlN��e�7��a��^V-�M� c��r0�L�p�i��:[�$�Ч5��""x�0�Nc���m喫��*A�Z���'���������~�� �P����)�;䓄��{�R��i=���n�k�7C��`@'����8��X���;z�̻Tn2ei�Si�+�4�y�o"����+ڇ?d�|�b�v~�$��-��Fݯ �����N�;��h���,=	%�G���s��1�{�M��s}��ΧZAV��m��;x���l$a�D	w�h�B���50��o�Bo���ҙZ��� [��~�y��h������S)�<�^��9�C�SE#��OP��(�}���b�q\��a������j�{�]�=SI��ajM�W�}M�@�uƾ������_�5��t���p��(���ϩ=I�����o�fo����\��Xչ�<!ݐ�&8M�v䨐K�d[�!�Q��W.��O��OT�w��wv �St�V<@�Ӓw�n�E�x�S�� �P0#�9�q�GX�Y��B焷c�4T�����6��)ah�j�l{�}�ջy�Qo�T�k�'�h&�A��bI�f�;G~m��4l���et_��� i������2��,��������p�9I:Ŵ�O�f�����4%�I,�9��6�Z0Mu��"Lu�w�.'�Oi�a���W��XT�2t��,�*A.߂ǐ&���	a�B�/�݋���*p����.#�6��ʛ]$_������tm��+�K����ª���t&K�-ʃyr_}�nDB���_�G��s�+<e�	k/�5��֣a�������k[f�j@��
��:Qƌj���{�ݹ��H2�����~JD�b@S�c���~�uwԤ!׿vVv��ڎ�М�@�	}k,�����3+���Jj�1�9��&|@������A����W��.q��3�<)"� ���"vHo�t�LSA]Z�HS�zF�2�'�a=�՟Ĝ�҃�)�چÏHw5C3�ܝ����q�xA�=xm(�D_E�pmw�TЅ�極`ˑ���H�[��ϙ�Dvs��&t�C�w�&��-y-b�o+l���+�Y��҈^rT#�ĺ������w����<=))��M���IS��PA?��Un�����S���z��o��*���mlC��|,��_Ȥ�]p��C����Ȅ��bi=</�1�c���]w,уS������O�ʻ{�s��'kUu�|�;>�;�Lo� ����_I5�U
R��v����7��n��W��K�`^���%2Ϳtf��7��@���<ۃ�%&�%U;օ]sMc^�I�}�+��kc{�\h�9	M*T����x�J�N�E_�c�?�]�3�S#hr�0!܍A�/E��KtT�����D�������P��{X����5��@�b/Qs-�Y�g���`�m|��g+�*�Fa�l,��\r���;埊�8*��5��9S�*!���L1�~�D�x�['��n3uV2�l�K�lf;�D��N��;�W�u��X��[t�~T�y������D�e��E�x��W�a�X��ݒQ2�՜'-A�w�
T��c�{��#vم����'�Ť8�1��*o.OA3��<2�`���C��]�t"�=����4�"�Et�+�=��T<ŦA ��>a��"BF8V��pfq���P��`�c�#������Xa�C�RF�*M�p}�D�P:U��+��p����)���v� ����6�w��d�-ſ����j,ތ��[�7W&��fKx��𮞛�FH\\ԝ	d,Z��P\��k�jSA)�L:�vB�F�݅d�
o+�U�W�������[xE�}a�H* ��#"�%=�4�%�HJ7��ݎ���20t��w@�����޵�>��������]tZQIؐ@4��{W� 6�J�9��}�_L�����%�� ����:*��������A���=8'�F~�����R���O��r���Ɖ��8U���^'T ����~"��4��{s
|�'/9 >�<;oV�bFio��Q�<�G�?绩
ֈ����KtʥI�#aC�)����w��|י�u�>�f�n��<�0�����4�1�CF�c�O~�'�o64���#y'���F�2��M�/6��`[�78Z���˭X��{�_�-5qgz��83F?F{ >:e��&�Hϔٷ�.�&�uD�W8�������<�.[���s�#�scG��K��2�����^c�8cu�	6�Z2�&
��
��`*��� �Qf0� ��a�[>^�)e�N�v���YZ=�:w����H![�dU�NtH�$h��g��+���l�s3��+�'�����:�l��N�����7(��J���O�(Z@W�)!�lb`V��Ʋ����� j&�jD�����\��7�2k�͑�ݗ"9��Aρ�[�ߪ������07���\��T�lN���^~�����'�Z^���Sx�0�ۃ��NL|�':�f��t ]j^���ʸ	��W��d�;T?\�ud�L��_0���R*����ΉG$'F�";H��p���9
N���M���(�ʖ���}�N�Qђ$Y����U@O[z�z��]!��a@��Bĳ|<w�!�y�|=i�[|C��⣭��:	s��X؉��WC��<jY�A�6"�4�uMw��$�d��Oqyi��
�Z�(��0�Źݺ.��]�T�e: R���}_ �2�J�6��r�cD4�o��(�t~$x��	y�F2%i���Y,Z�V���K����f�|��9�	d�L������9A�<��(�� �ψ��S�i��.���VL>l5i���]���
ȋV����Y����U�3ޠ�|!�9��f:u`���i��wh�釐�?���H��AZqq���Fl�	&��8VR3AQ����{3�¼�v���S���~yjYGa�q�Q�m�saۈu�8�ĉ[��z2�nT��:^���q ���*?��^�)�PÕ��ViKm��؟yү�k�~s�v�r�#�\b-P�|�$���� � 
"��I�����a^�
9�nx�p���~�O�M�[F٣���7A��AҽZǉw�\̃������"�Hb��A��faԊ@�\dӾe/F�q?1�pF�㥞�\����5�K���=Y����!�x1�E�Rn���
�pHekzy���C3l���8�5OQh.��X� g�+�C"�W|n۔7��+�y���|�8�9&�$2#��/����=m��Kst< ��v{�;�33�fP:�E�<�OwW�����z����m[��ц��>h���e�}���Qt#�-��T-�
��k�=v��"}��F6w�~_�@�_�0b�?�z/!������7Ǫ�`ǝFV4�\�����;?��Kue_z=F{�2U�C�! jD��OX�oH�۰,�"S���]͐�(Vs���Ȏ�o]$ǿ1��ʮv45CLJ��V�^��^XS�֟}��v��yyBzV�������I�E�
[,?�0��"+���&`X���2��CPU�_`���d�M�!s� �;���c�H��6��˞y��.�&�C{D��69���;c���p{�ո���C�A<�T�-��;/���i$���N����˫���b���`k?�}m����}��83ԣ�[)��S�FV:�w��*+'ɗ��&lyl�#�� %3?p��	��4�9�pѰd�D�»�(]�3�f���_/I7ӈ�J�q<�z<��Aq���oC�9Njӌ��۲�o�Ө]��-m�A�F�r�r�=�Cy�.������c��h?1�'b��׬���O��WF�/ńC�ܗ��#��0R}]l���>ϥ�j�򵟟` П��prpg�� Ņ��>��Ҹ7{��w?儵� ��w���:*�;3�հ���ɒy�M���U��+�*D^<6_�y �u�i}#E[�[mKOA��i�Y����Q�U�geV�k.�h���H-���>�4�u�����&���"G�u~���ƅK������]F�>��h�������D�w1�\�+�#�g������]t�-�����x//G�pi�ң��`�f�/%����r8nI���m�ʥ�/�QvP�:rM���֓��%��]	&�]���4q"z�������<� ͓���y���K���P)�M�\>-�U�C�?3b	8&2��F~���
M�2��ZI:*5����'S�1�]��@�y�xቖ=�n݊�~���$6��]���v�.���!�[�?�׆�j7I�U��m�4Q�\9�c��t�*Os[���Aw�'��խ���={=�Y��n;���t�%^�^����E�J/��ŏ�H�K�`���#pO���c�`G>b�l�KA��+�y�/��~§eNv{iB�h�i��b�L}��3@;'u�vBXGq'j��5O�T�Xhn����,���;�GW���4t�|cU�.��e��������;���������9K`P��~.z���܇S1pp������"��8�.>�mJ�lIQ��J+d�;��X�����MF�~���<lt�h�ap���oP'�
�++�y��5�W<zR9�1�uj�,aenE�@�W��i���UMv<�3+8H�Pn�z�T׵QT[h�<�����ˇ���o�K���Z3�/eI����4�=�r�Z�"0����_&ɼ��b��PJ2����=��-9��[��ͭˈ�u=6S������co��ɌT=p����e��0:�5�4�䊡~�e������8��*�J4�����-�͞˯w���g>�~��婀���{�,M'x��B𠪘��|���T�/�e�<�y���'�Y+�Ś�����KMh�`p|��o�G��~J����z�����Za��f=J��x��v6.\��~���]Җ�4�����'q�B��-H���H������%��/l.�o��y�T��7�_�p�5ݙ�u�y[�r�|��A9���r5�ӥ��Y˟�|v}D|9P�O�.}P��X@O��K�T��s����h�O�l�u��Vy��I��������nvYY���DW�Nw��y(���"�WxH�bԣ&��>�S.�0���JG���꽡�r�yI؍��-����CLڪ�׻��e��;�%�ӹ��f]yu_k��� �S�?�S�}��|l��Q8"R[]�`��$��Ua����=C b�\�)?������ګ!_i؞����n��v�ab�-M���s�:����Gp�_�)?�(�	��#lo=)�c.�ؓ
��C�-���k��!=�/ɲ�Dݰ�Zi�de��������h�7�U�$Fs+LK�p�׮%Y�>�<�i�`�W�O'ߖة�f�r��w	�?��}�n��r��uD�N��3񋛇Q5&��l%c^]�~���qĿ3�G�E�-�14U�̋��Kĥ</8��;�\��H�wGL���d����!���=�����B�kﻨ����ca3��Q��G��n@mI���F�iO|��cY���Uv��~?�޷o�=�Rh���ˊƭa�`vR.��|�ÿr�z�1kV�Fc]�v�/��Z��]LQ�m�Υ�ߴތ5e,�m6D������sG��Hy�|�z7�F� i��e>����v��	0�F�ްj�q��t�l�%򦟮��W�<���K(4�Z?�*7����>ר�<��$]�����?q��[	���O�����Ĭm�R��մsC�ݖs`�\w.����O<��3W��TV=1�x�h���[��r3�7;����=h#;�|��Z�B@Z,���[;��T��ƙa=&B���+󢌔�w���[�&���2?v�g�u��)Pf��;�\��HH�A��I����wn}�ͥ�<�w���_~����ר=�DL��5����} k�-���%��6
�����<��7^�aIp!�ŗN�M�Û��׻�C|�9�;ą6sY�^���DG��n�f>�}���&'DC+��e�s�q�>��6r����a�f��+����m
x��B�U]C�]]iŝ�Q���v��y���>�ۻ���ޢ�ö�Q�>�udP5jͤx�,��',IaT,�	O���WzQ:��䞑:���ø7@��#X�d �@�!}"Y�T������}�)��V��u��1��w▝���Q���_}aH�G ���9�\|�!���X����r��F^�i�c-��w�!�q"p#�n0'����{��0��i��W&9g7ǒ�K��Hn�.#8�7\9"��Ȃ���S�0/�.u�o�(�_��<`�r=Y���je�"���w^��@���]V�0��4kHDR�����ݸ���{�<�ѱc׬�A��X(�@�:���xF�7`|;�D�P��2���̧�7��%��C�3��QM1͉q�|���Rv�k\-|��n DVK� 3����S��q�����#]��UAL��0���c9����?xD<�d��b_�Qo�E���|��7/�[�����ڼ6�P����L&�~��'e��-5ֽ��lc�!�y���OiL�}ص�s|"���:tK�]A��x�n��XZ����0��t�d_0z��^E��W�{MB�
)�^���F��o�
���]Ҽu;3<S��e�&�,�n�
���e9��[k{4&#�l�-v@E���a`�I�r=#H�k����e�H��`|� $ѤK��B1I=4����J�T��
<�u>�T��Z8�6��N�_ ���
�҄���Jꌕ�iQ���a�Q���<��J"��2v�>��G��T�ޏ%j5���q/���H?��f�CE��]�[2�zzL��M��\ZN��LHhOP�E�s��c�dT���{��D:eJq�$#���W�D�$��*;ޯ��Z���(��(2ɪ��Q�<	M�{I�jǈ��s��+E��{C�j����ݥ<2�-+��
�l�2�4��W����0�M*Zӓ�П�UK��6���0<�Z;���ΘV�I�ˣ��c{ȩ�T�|I�|.�/��~�#��k�k�+�r��h����$��2��-l�,bd��I.�^0�#���ɖ�J��L����fU=Β/����B�Yl��Ps�g����fj�=H�`�N�:�ᇝ���Od1h_���ɞ8R h��_���9���b��i�I�8HW����|0R'�-]:�!M��5d�(�iI��m*��Kz#�����o��H�
�U���e�����W���r��8�@�Ŷ��E����	�Q��ە�$���/ɺ+�w,���y��t&�I�=6%`}�_@"����y�-�V����\�|�	8��1�)�v��(��I^�>]<I���+�=O�h��ֲ���DH���ۊv�ws��ö.����Ӣ��l�6��y!��7��^��D0�gZ_wE�_-��RN.S�P�EW��oe��������°���M�L`�z{k&���U3W�(�m/�D>*P<�8�V'֘�����/����yC�6������]�e�yXs�_M�^���k.&Jb�2S/IX5�tt���-*�
ܲ
C�D�l�C&��~�+.%�oJ8N�[�
���g��h���_�Z*-��џ ���.��G&�V��-��[,L
���U	x��C��{�S�+,�7���Y�M!}�m���y�~�N�����:�����y��:e*�� j��5b��{��-"k�Gz��C��4���A�w��«�CBR�W���Nj,׀V�-�}bS���8TmD+D�'��(z�����
�N�.�IE`��W��Ɋ�9 ��ؑ��I��W�f�,O~�m��825è@>¡s��-��ֱ:*Q�2�`Ӵ @�����q}�'���!䇈Ta�7���E�~�?�yn���q�Vh��g�\�;��^��DN�d��c߼j��kA�Z^L�G�L0������]p���1�,���Xh�Ρ�v�����mԓ������Ԏ��{C�1mJz�nF�:DEe@�(�q����IǨ���p�۽�e�~�Z�U��׎=���6�!���d1B:.k N�[��+�^H�Z�Q����a�Yu6�\OҔ�}'���Tܯ��Yϗ� �^�ԨX�>s�}��)s�b:�v�݌pf��\���<t��MvM�������%���$uCX�9��k?���<�&YY	���xu�7k|u]ɤ�֗.e��i�� ����^����42d�[SЭ��;<�o&��郺��˨ފ�cd�e���'G��b�X�c���$�r�ku�s���e��y��u��~��~�ֈ�`@��.���pa"0����w�q���1��ix$�:�[����Z���f�o�����OEt��7�D��H!�(�k|a\87�������~�8+�n�n�E�E��*^^�z@���������d�r�"ć�T�I�X�>���=�l�1��G�k9c��^�Yd,4\��ښX;ʧ^�E'����闒�2=q'v-V:jF��;�Y���|䨼Gs2�M�B��r(|q{SZ�J4����auYZ�TP9�+��?��5�u�����|{�����Bq����+˰%�����퍜3�V����|Cim�^���k�s��镛n�b�<Dza�T3�")��Tq�]��
����[�+5��ӭrC�˩��/�|B�#��
��$�+�	I���ߖU@;z�#VN�=�9OJV����)�2�M���j�_�Q:z��d@g���bX�2k脵�W�]W��ep�ا��0���]��Ӻx�P�g��M|x�wLV̓�{�+j0�����vJ�փͿ��ٍGh��Y.6p���.�i���,�GC㕽��:آ�P	<0M�}�a��X�#.V�"��8BkDK�?6� 6�V]�l���T�&��/��h���=�s�����TXIݬ`��[1쳆�T���a஝���V��G�>
�zt�`�g\G��o��7�ʊ�ah}WpK�j|����yS���'=���ɱ�[,H�NW%YF�eke�K	���-!5���	�繖N�h�1��3���*)I��'ަ��W6�����vi��H���W�f~�O�����dv�����lEuj�b̀�.�UqPur�_
ͼ:�^4G��Eu쿶���<�"=H�Ɔ�Ol���~�Ã����v�D;�ja��7�&[o+Uc���Z��xdA���Q��n9?�i�t�\jF~A�[��^Rѯ+n�f��2�e7�|:�Yo2��%{<_��TalP�O$&�N�� ����"i�W [�φ�\�i��.ݕy3�&�P��.K��Zr�� <X�4���P�6��u���#wߙ�6����D��i��;{����_n�'�������%�J���[�y�\���(��?��>�@��b���E�kKa����V[���s���
��cp|��F����OQ듶g���,����96\��	��p6�;om�]@��K�Qq8� �{�)Z��r�5�S������kw >�P�֞���z��Qd�<^KQ���}�<1A܉����Z'y�I[�?ΓU�>�?R�շk��4�ޫE�$ӭN����ME[ C�#5`6�'��� CW�${��[��i=��x@E3��z;wn�%C�HJY�#�������{ �C�M5q��RԀ6B�`3�0	��"|��Q�_lYȊ��E4�]y'��K�H��k�����,����%n/�p��'��{kx|f��/�x�E)��F�cc��4�qȚ9��5��'����r��O*��]6,<<�6��?#���+a)((�,�ov�d�h\���3�N�I�!5�xA^ ��z���T��ϔ�bX���PHc�ue�u�gơ��=��>�а�m��Lb���7��7]�
{���L�����T(KO�t�s�^��N��?*���zR�,�]�������e�����w�N�N��n��-�Zq
�V%}��4_2z����7�B�-��2B1���m����A��N�y���W�μۇ�G[��㝆1�g�Nhph���g�l �㪮.EE37hntFxU���K���#��N�_!wm��WM�>�ƀ�CD/'}Y
���_���&
��|<���hQP�((Ko�!0��x�P���8�D�,���\|sR����L�a�m?�z6k�v(�H�!��=9�2�BJ��z�%�(�)'eG��nj��YA�F�u;����S�f�>Δ�7OQY98b7��Ob����<���1�y�_��?�u���?�%kV�L&���l��^�mM��Q �2Vh[�P�rn��,�T9-�B;i�W��	���Ѓ��[�	D�uԘ���Z�_��5%���"�� #���..bMH��)N6*i��5b��d�����긝-'\S�8��3�˼�BqȘoQܶ���
��?Ca)�ћɎi�wj���M~׏5+�M�꡷5ܞ6�|w3H�}��!�c7��aqR7��>�ٖ�_��7����C�_�+�4V[k1^����C�j&[�Y���#���ѸC�z�.L��<�����Y��h�a�a�����t�JI�su��u�������z~�H �@�ch�ݲ" �|�vI$ٍ���MzG�y����7W�aNb�+�j'1�^��S�Ĝ�r����9��o��VCs.���F2��+).3����g׵�9썌��^�@j�/���K�p�I2%����:�����|���8��,��AU�?m5�ȗ����@+*�)4��PMnk�E�c��5�ߛ��5bѤ���  j�Zc�۷4�#��ff�&Nnq��x�G�dN
c��@ �6�2���?�nf�N^��2�/�(���{�l�3OSsO�x|-����=gd����̐qss緼h�)@�.���5�	�kv����Wx���m���K�zMfVHF��$ŉ�]�_�n_�D�ʵ�=M�FE��r��;C`��ͥ�B��U�[�ʧ�����@i�O�gMY=��ݴ�/�ÁJ�q�I�}X���-��:�=׾}D2���h �D�A�N����m_~vxFWJ}ʓ~����b���!F0}Y��X$?�b�3UQ��?TP������]Bh���p���񓺤g\�c;��lH�-B6S[(�P�;��x<V ������Ps���p��e��뼗i�`��_mI�C�ZC絰�5x�[`W�M�볞��|�������j�<SOga	���Y�E�k��9�s'�"�=�|�#��V�yv��.Z<���A	3f�~�k���=��¡�xH��H�'I�e���;[2��;�m���$HcoG�խ�+��\�����T_9�ayl�X���? �H}>A󹵂��l%1W��(��Oj�,G=I�ZjÀ���]]��A�u��QݼLo��(��M�.y�^%a�?I�ۘKC�ܢ;gD\=X(Ш��Ο���b��{��'�o�Rҡ��-A������f#�;n^���<�~��Fm;*��&������ц!�{f�8��WL�C��3a�O����׸�T��)�վ�Z�%�N�M���i���D�9(�l��f��9v��������X�Ce3_��or�7�+�ʟC[��s���Ở�c�������f��T�	Qg�8-9ݡ��&:vf�k�&�Ɛ���`�E���V�le�e��k�bRgGѲ��B����Ј�ac�nx�^^�Vg�����`�_8��O�#�r�����;�1#��'�v���o�|�G+�&��F�Y�.,%,��������㤆�(\���)�o��$j^��W�7��I��4#Y�tBν��0�XKt�l���Խr<"]~w��^�3�u��<)Y��n�{��F��>����4�[��i��>
T`��8�>T��E���\T|od��I�����&|���Zφ,���;t&�"�uC�m+�ϭ9r���Oԍ���t��)me}�v_-O%���槩��\��R.6�B�j�F���"���rM��;�^� �
��[����jR�	r�zۈ���s�G�\L"�D#�;\�M�d[�n��.�D=	)��f�,�b�" �=�vFQ�IB�Ƞ
�ÿ$��c�~7O6!�&����褵Iڴ������!��p��O�~pív-Y/3��ea�N]��STn��-!A���h^{��h?�Q�R�d& �`Y�	�jk��������Wr��KU^%���n��b66m���5�4��t9.����g�C8�6���d�Nˤ0�R�g�N��b�
��C�(�\(�ޭ8���HG������B��}Y�6��H�ނ|�2<����)�m߁�ܾH��oF�t:]���E��7�]���
�\�rw�*P�$�4��[r9}X��7=���Ы�-��y����a��9�dt���D
 >�3�{����0�7_�@J��TN�-�6,��4�G֞]�	}g��p����Id~��q��&`O0�"Ae�!�|�#A�\p�hB��\~���H-��|*�Vf'Om�N��e��e�>�i?�9��ݳ6V<]�P�7�@�}��FQ��M�g��/�'Q�/r�}�����1 ��S����8�P�u�Ȕg�N�0e�5�? o���ҡA�o����,��<�!���'T�������8G+���V���=A�S1`�٨��ԩ�ʱd�\F��"#/���!�_ڰ8�Zz��3�s}�>|�y�F�f�r���c��gz��V�
~���OE  ����aRjK��7(H�ᔲ��s�H��q{C!,����I�������Z�x�¿�*h��r;@l譋�7�'G�D�{�2�fַ�ć���j���`fe�٨y�q�Ə(훖�t\U��vTR��P��?��s��1��r��U�HnN�
,�����{�uͰ������k�>�z�@e8�|2j��7M�����a4i_j?1^���HҠ\ҚB����[�#��0e ��55	����/���$^8�<��ҕA�t[�����_�[�MGF��v}6�B^Y��xq;�Q(�(lt�wb��#�
�J1�j�α@!,�)5�|�Px��'��\f�W��AE�P̑j�o����$7�D����V:v���h9iO��fA+D��p��f�r}"����,�0�����~=Q
yS�ST�M�V��/yf��"1>m���ѳ\G��H����F����1��/�N��{:������n�$�v��Rם~Y�i&��g��+�����(9��aq�4�?{����$��v*�����g���N���K/o���� �Zj]�8�(?@l���:��a�D�4]&>��sE��Ms�HZ;U�C'A�ژ&���(��J��t�M�CM���"�J�fI�����;�.����fS8^���H�<l{��<(V3�� �i�����-'>�E��P�kf��O*Z�@Mc�<s���L"E�+�K�h�[E�-���vCC*�hqi'�3��]Ɇ�8�p'~�U
�����ˋN�1���m�5E���7�/�%:V|��;8���J`�	ҕ��:��.w^T\T���:*Q�}���-�,����J)k@��H�IJ�x���D{K@�����"�\��{�`�����3B��?i�u"�^�:�+6q2�\�]��3g��%�K�i,�Q��ˎ	���GCi�����u��I'��v��Vhߤ鍅n��@f����F��m뷗B�Q"{�+�*���%���T>�L�ʘ#��~�u��u���B�G��}jG��Osp���nݶ.�aU@ZI�3ܝ2�c���}��&���U�G0�V!�����ħ��7�J�S�����]�"��r<�M�YI�p�:�E-n%V�ͯ�{���r<��g�M|��ԏ̓?���ǌ�2�������G��U`���Z�Z�l{�#�_~uF�{�����j~������N��;�"�����-u��!Of�Wy��3���V���=o!__�3�o��ف�?�+k�]��a822$<�J���6��c�e�K_����&1��_�3��,����1�	��C����Z��*;-�ËaJ�������@z��`G�H�@6�]�7ep8<v"ƈq�YD���X.�KW��$��9?1I�TCQ�e:v����惜���0�]��m�X�p��n m�dH�+��a6�/���>l{fQGC����$,��Z�K����bR��*��@�w'nF)$O�Ъc2�O���xS4ζ'tk���)_;{�÷�C�A����v�ga9�Qt�+�D��qw�
ы�awn�[�S����b2S=�gů�V�7q��o�6�]�,�O�BL�|%nZJYU����-i������/���g�Qԓ��y�::�ꮺj���>;���;g�V�p��G����`��2Zҫ���E�Ya���ƙ������؂%.=܂� dp=�A� i�^�E'� ߝ�Γ��i�Oߝ7t���A?���5��ѪǗ�OHnL���:���1�In`Qps��D/Ğ1߆����6�?��X慎�ݑ]�������.�����HU=���e-���}\ۀ�抗kX"��ԕ�0ֶ����$z5B�+�|o����-Y&aźԳ�� ���z�z2��uW��QHL��/_Z)]��@Nn��E�=up?ؽ��/����k�5Ř7�N�#7�L�f���`����x�:	�v��\]T���￷ P��ne}x�F������� ���>��;��2�_�9�Խ�S�����q��[�l�j�aҬ�:]�a�C���$���2��g�t�B&�5
�)魑-\���q z�X�fȿ��j���cwď�\W#�p��R���I!����|�8�˟�"�x���ˍ��>������S�T�MC�~��
���
.�E���](:�T������׳*�q΁k��N�&�p\�����%���<&�l�)5/-�V~�l��5��i|��\���zF+�C��d���ޮ��x���^��@��H|��X��#|@�d<�����u_~h�ʹ�_s8u��X�o�yu�[R���������֦u�M��v�`��f7�O![ݫ��m�����bk#��'h�C�����J����n92�l��N��#�4�[����_A�����ϙsʟ�8`��J\NuU�f']�&-}Ɂ��b:�����������zN���+�� f (�x�f��D�ןIX6@�mbܲ�� �X��hs�#���i� �(O��9�\�|,�W���
��db_Þz����.�u�G�Gu�����Xf��$f0`�2�^�dw�߁+zެ�� �����;^lܼi�/L����v����=*���P��-�>'�/�fy�3p�e��~hGQx�ǈ�����a*����Id�+J����GjN.Md6c��|SE#˜�	��>i|��V,����!0�������C�j�,���W�3��5y��4A�CA
��h�j\Bc�xB[+֑�\�s�t�Nz�BZ� ���c�V��]�ʿ%Y���V�!���(��8	j�^I��!���!f)���敘��H���%ob\��E�%��^_ڇ:���V��ˊ��C�X���w�v���(aG���N��-��A�+� �W������ϸ���r�MVZ]��G.�M�st�h8tx����%��&��Y(�0w�~����#74',G�����PT e�q�d�kt>�Z����;LKy$#�g���ؙ��yRL�p��zW)��":S��5�X�ل��Ӂo��~��ڠ�^��� �n�X����� R��Q}�� �&����	�k��ݕ��N�(�Iq�d'�C:���M�M�^o��b�L��S�B~��﮲�W	=5�܈07�������DFH����~1�kf�.bx����%r�L��������i$����l���`��������q�S�f�QȖάcB#�|,�.�auh��GmYf�'sƀ��̘޲��VϿu�+��������~	i�jm�,�]�
Ԗ�
��'�߁����٨S���t�j��|��]
֙$H�"�e�A"�.�g���*BGh"w�_�,��p���Q���o���R���A��"ۆ㶋�l`��gP������N܀��0�ҩƇCkE���X��e��?�^�0��s����8�8�T���O��jm���M��pW�����pf�t��r�.�k�%z�"2�C�?����d8J+(1�TQs�w�}�k�+t:�de� ��T\y9��bC����\f�Y�u8c�}t���y�p��IIL�+��^i�^��Q'��H�D{3�����+ɾ�i*z�;��ޜfMVCKO;�q�����_��S��%$
��
q�5T��q���3#H�0�z C�{'���0'b�AZ%��7��9���yVWP�تKhG��IL�`������v(]���qN�T�q����WuD�Gz�k���t�9q�/~B�����4��)E~���j����$��>_�:v�F[jSNj���%'s��}E8�1��0��p1�J(��Z��m���%�����Y��::�0x˭�n�0
�a��� i6F\e�G�U�0��;<��7?iꜬ�|�����Ȍ.��9.*_;g�#�ߓ�����ff����i�j��qcǊ�-(y����'��Q�3~I�S�5u7j�Se�a/����z��XO<Y�$gh#�X���h_4�^��܌�-2}D�jZ��tS��;�j@��&��2���&�7�V�x�Ҟ���DM�Z[��lh��|ۉ�� &ΔP �_p�v}Px��)?S�7z��Y��z	���P��aÊ���.֧-��X�ߑg0XS�~O��}ف����D���������E��Y��v�1��p�vql5��6�5�	Vp�##!!c��G�3�{��kIF:Ϣ�r�Fbd*�ur�{Q9�h�&�?��-g�{�{�ԁ\���'Ea�q"�	b�Eἱ�=�!2�>�B�X��;�B���ⅰ-��' ߝxg�|�����f��Â7��~��`�x���0E��W��4�?���6�8���Mq��ǯH���h�A����l׊�����V�Ƃa�W��k��P�b�M��5Ԗ�F\�鸁���N�(���vx\�V�?�&A�b��R�1k��e���oR�e&�3�m��,ؔ%���Vs̞�65z4�ۄ�ܮ}��<�j�ѯ�@�|���;��5�gϲd���f�6��3QU��9�ʰU��ģx21D����	T�xa��҇�)LhV~Ve��Q.��g�f��<�߹Q dӘ�K}���QiX��xH[=Yj�����?����到��-k�9ŖܪU�]ܚ�=�ϵr��5�j��|��2T1����Lʅ]��t���"U�U#���~�5E�;"��~�jܴ`^Ə����m�њ�-d�mUx�j����si��ف�5To�,��`���%`��Q�u�,���O���lV��1��|R%�t��T�W�/�V�I$��OJcڋLsv�x��D�#X����xK��	��&9Ari��5�[g�Z�ܪC�����+yYՄ����H8����M��p`7FGֶ�1��樨
��υ�YʾH��O2�Q�fY1��Y4�I�x2v��D2�vY�| �Y��5�k2�F��*(�" ��x;��j����>�ۃ���2k8�Ze�Ӱ��,�
����e3n��Q���[O��2��T���G8�������\�L�"������O����ս�^/I�y=�[˄�.��x,���B��C�41����iK/	����&�)^r�u��췥PN���:$p�y����$fGV�̛i����
Y�>\��ۺ|+�Y"����D�뿩�v�UVsȨ��#�ݬ87�Z\�����H�=4t������8l�����ֶ�0�cY~sB<�3����ı_d-���x�)ٯ�A�d�3���F�h�&�ɬ�*���z�F�����@�gl)�C����ܱT�֚��ϙ�c�G�4��V���O�d�+�~ &���/1Ü.������ʷ��x!0��3�L�E<�$�*�&5�=36���t�*d�+'�ٽw}=�8>v!����+Ƃ���g'Zg��1=��v�O��n!���C�� �-����,���o�ц�Չ�>�ptuO��yL
H����OMˋT��9�kd�� O.l�=dkHG{ jUզxt+i� r���Q��ҭ{m�{��������R��Ǿ\iLջb��^6��s�#��p|$p-O%��`��3�tɏ��C8�u�`���ل�uؐ�@s��Z���2z��9o�I6��!�:��X10@�P�'!���ÂN,�\cE�A�w!�k��A}���u)�i�b8[Q��X~���˲�u�	�y�^����g�d��Vws�U}��(����t��+:K�n��*�kXN>712v���:��l6k��u��Y~NK�B����v���T=-vf�p?�����������r�Zz�J�<���\V\�M#�m����Q��F:��V�_˃�=�>1gF��#%L�X^��s�n�@��~����4cs��R�H����h�C(_I�C��'C��m��ez.�XV�4����J�g�k�je��_�ׄ޾m!*"ҥ���t����HJJHF�D�.)���"ݝݱ�	l0���y~���kw\q����t��]N���oI�5fՑ�Y�ӹ^������_�����83<S2"�0�z��_ϣu�h��Ok��K�V��!Y/��gf �8���D"%O�5��k��%&cv�-�y�'E�)aF��b�8hZ�`/��+f��W:h,��#�8-i�����yF$,�C7F������/��;<�[l}]!��)��[5�$�y.�2�]u��{���^�h^�X��v"�+��ǧ�M�V�8�M?�h�b���'O�W,�,��ݷu������x��,!�_

	�~�i�qE[p�x��_N��=݉�I�S�����b�f��h��%�8 ]�z�L�/"^��*u8ZF����(x��囗wh��(��A��n�ܐ- ��I�Ӫ�n��M�?S/�?��c�y�s��Z:b�:�2��Z��3ّ�[��,6ﰖR�m��S�{5X|+��EF=��y_w*�}e�v���[Gc��XX�E�B��L�C���\ԡl����%��z�l���㤘�{����ZO��£ud:G�����'(لpΈW�N�e
 ��_��h�C�.��a���e��I�g��t��kW��g����o�@o�]�o{�M��R�_�x�=+T��'��&�ѼiFF���
_�b�e'���D专p����$�7�������e��.f3-�_$�l��6A>�hצ�����&z=�&|��Yw���9To߼;b�C��#��QM�H'Y�O_��J�<�����[��0
�G�|�������Ț0D/ô�d�~�/�5G�^3�z
R��1�
H����7N#od�Gy�y>U�@�|��"�i�5��yY�䇆qO��~�eQ8�;��r�	s�sR�y+��뽮r׶V����&�:m���I=l�'�-p�nUu,%��f�b	%�uI�/>)O>����{�j�9���a�����c�'�1�9o��H�t��Y��2�>qE+U9���z�r-����@M�O�q�ˎPB[�����l� ��Y#���iGk}�[=b���U��C~ARU�CZ=���&K�h���[����xE���r��$����1u�e �oك�(�j���'�����D6�c���J�l��1����irC8_�N �U-�4�;�f�	˒��p��m�c ����'boŘ�i�f�0O�B5تJ���Hb�aE�;�	z2�?O�5LC�6�:��ɣ�ɔ5]�>`��H�b��r@����O�m�ܳ��W�fW!z.�mx�����u
�C���Otx�����=��v�����l�Y^Ș�Bi��DR�/w�Fi)�$Do�����>tV�y'����590ç(��録����肜�Y/�卂���Y�];�V����O�G��V;�Hd����C)�4;�l	I%Z��Q�qUc�HLa���?�_�e�=Ah���)堋��HK���Ep]�K�5H�Pd<5�;�k�I�J	;;qT�V>�j!��;��}��!��o�c�.����w'C�Am;�h����c�$.����|��1�kxr�C�l~��w]�ֱDkV:��)��x��Z�����慪��m}�z4]������9�5�j�{���dmHOȄ�|$*����ތ�]9͸���"����d2�+ck�I/
xK��A�w�$t}l����f����������n���Cq�7n:	��g�O��=R;�؝�ʹ:Y��1v�|W�T����yx�Z^����xqs�d��-������]j�7#�������S�!��^z%N��j�ٔm���ڥ�H	����?"��G��j#jp跥��2�L�QM�r��Yy>Z����va��Eb�s��9�4��G2d���u��鏭�ą�n����\^�;;�F�}6�t+���E5Z?jTJ�x�`�K)�H:'�(O�.��7y14���Ι�*u�ԣ�W�JX+��L���k7�޿�JA�D�����@�d6��h�`�Wj��b8:Yݶ&/��4�$����gdWy��>��%pV�����\��BF�d	�d�j�r*ҁ��=9BM�s"y�+�L�Ҵ���p':�T�O��8Ɵٸ�)H{�=��=��E���Y��͓��Q��w쬼������4�"[�p �O�VoB���#V<9���rPf�����y�سT�|1?)׬���?��������[uCc|tc�t��K�ŢX����lX�Ω��P":�"���yHL����֍Dje?���0������$�Ug6ٰR�aR�|,�֯t,��ӧE�ku�-���������QN�7��3�����&b�o���x�����h�d� w �2Ր l"�/�H֏�׬܁�F����B���i4S��n���i���������\[�R�y:�H�)������B8�Btwf���>6�K&�譠�jF;l.�������֕�n{��fz+�3��*�����#�۩�\>
 P'��h�Ͻ�s�d<P��(����>6��y��<?��n���翰n/�˓
��ͣY�0��+�)I;ͽ��t�M�����*�J ����ũ!U&K{����
�E�/��K7��*e��e[GGqy�x�Yff�N����͇<z��XU�`�4 ���.�To��v�כ6��]��ZxJ�FK�Ve2��!�>KM���.��2@N2��J[�=�ސ54��r���!����1�
���dɝp���j�=�UH]ޙv''�<�e� �R�O֧��D���-m���v�|��Yg��qVTm�����롌-9�}�n�@����I�ò�7kVH��:����صr_�e|����~!�ו�-+wǄn�]-��3v��E���'_�Ew8����gA�'� ��~�h%�QdK�j7��e�dN�XV4�ޤ��O>8~qE��6I;1�m���5sz��k �.S��r��h���'6dZ�x52LO�Ȫ�K�[�X���3�'�����[}��B�;���x�>���ى,uhfQ?��u~ߏ�&q#���*��j#�;���<�l���7N+9����J�|뫄�bvt^j�Wd�H?
�h��
FF�c��n�<%۰��w#��F;׼s�q�Z���E�UL)Ѳ��ک��L��e+6����C�$�-M(���y��<%�7�����M�qK{V�DVY܈+jH��l�x�䅈���\��L�4�ܻ/x��^_o°o�?�;0�o��c<)�k�3ɑ	�^E�qme��$�k`�Ih:(�J#�V�l�M��7���L�ҩʻl�|fXd�;�Y�&��%�H�p2�a�M����=�|��6Uuϋ�P�����ҋ�s�+S��oE��@<v��\"Sb{q��OܿO�n�ݏ�r?��<�l,;��5'
�2�����6�*���䋌�2���CI���}.)f�9���x���M�`f�4���������2��P�5��������Z�x���"�^�08p�/r/d�E��Ґs1����bff�!I���=�ў��\+�S�g�T�*��˕6ʀG���^klE��.EܧL�(�R~NE�0#�ɕ�Q��A��k�w��V	�<�(j��[-���I7�ɲ��Nu��r����a˨�/b�q��l�/���)�!D<�[��=�Abk��ǜ}���I&iI�v�?�)�;'���s�Q�]6Mh��Tv��'�q�)�}*�T%~���EC,`t�f������&[�B�/�<a�;�;("6���n���!�?�oX<��
��أ��:���ph��c�3o<��_l��^	<�|�������^�5`ڣ�
cj�?��B��=���sG�0vz�q�����.fa�)�y�F��Ot� *��mU�ג�L3ʈW���n(�1y�S�;����7v2�f8�����B�Lbi��ؗ='��Zv+��U��Bz��}��H���o�P�Ҳ����=4͸?o�['�F�L@�J��2�mvh�j�fљ�����:����4q����]}��;&��� n� �k'w��iA7'��U	��`�θ՟���κØ�3�7��J+7�7�>sܸJk7�@-�v	��5k�2S�R6�{Z��{�_t��-�4lk�r��3�|��#r��(�V���E׻k�3�NO���z��I.�?U���嶦Z���zx��ޔ����~��bi}l!_t�Rg���t�c���uZD�Jt_j�dȮ��8�X��Q�m�k~��{e�3��w���:�2�]��Ӡ�쐌QL���Q��$J�v�P���\Nث�욒mP�S�ڏ�s"jN��Hb�LS�x�l;ZF.�I�y��4?3��A������g�9���~�}�w�E������?E����3��@�n9)�V������W��5P��0k�=M��Ԗ�J���}(��brЊ�t�g�A��<�)��;�A`���ؐ��"#¢��p!2�C%{�Ù��ڀ?zL�����2eP5s�y}g=��z�)�c�O�����?aR�"��	�/4�_��z��3�`k�0�;�@-Q��V���|5� ��xN�gG�H��ϙ��3��	�Kh�D�lZ�8G�Cp��`��t�\d<��trh��h���rr�[9C�$c�r�tJ`�6���hU�`�lU$����<���3�Μ_�z���p��Kt8H'�v�<8��6�[�I����֩�H��'K�PK#(�-��]��;bM�E��eg��hVF�G��S��g�MüQ2bIƐKR3j�]�¤O1^4�~���X�"4d:�W��9�r�/�d]�"���/���7�^�t�K�IOt�i!$�L��|.��C4����9�6��5�����]�?{�,r�D�!)��%��΀uǺ��D֬T?Ǚ�#ssc�'f�����M9iܢ1����]%�B�R�)~~�g��W +<��z6͖�JNԨ�ݙ��8�#���ӗ����`(�[��zqlEYk�	Gg��w��ky�wnn�V��?�����hf�pM��,�:��_ժ�4z,�$a�$��euqFH���~�RƯfĒ�������!/�$�LRy�)�p����-��7�k�Cm+?���ޚ����=�2��S�a�ޟcD(���m��z&�!k0�J�=;~l_V������ �|����U^�C�lȆ����@d��\f�Gi�iȋ�"���W��[ӎ9���M)����P݀c޳����>�{+�(V�iɨܰ��iF	��#�����@�d��}�ߒ�3���#s�Oɏ�� Ad8 ?sk����1���2#�-q۩�!����M�C��+��ă~�����%B���5Oh�j���Ƽω����<�z]m�U���e��,�L��8|�+h�9��/cB�/��M�%�Bw�W�=mY!'L,�c:��V�1�Y��i}�EF�5����wm[��ӻljT��!m��ӷf�e�Ǧ^cTLj�x�%�4A�>2�N�ܣN5����7�L$~���D��F��	J���7'�Rlށ�*pӺ}���}�(���`1�n�ɷ���/�	�یr&D~�S��
��[t�� ���6[b$�j�l��珞R��x��%3�k.�,�do�&���L|��g�>�6����z;6���4�~2q�#��>8����c�/�3 ��8�o(��Ȩ��!eu��J�o�w��]���ރ�}�߽�>�m*V�������MD,��%�3:7LX�� B��`�������Eѭ�c�y�ؕ[ѿ��V����C�����<�[��bxNdhOE8�8�׮V��Lg �AG宺�%��§�/C�,�e���M?c�hR�'>w���G��lwC%��;��<|�z4}P�<����*�]t��C�i��>����4O�V��ʤ��E�-��E�|����>ol�:C5��O�e�8j��J��HzlCS���ƿ��cA�/ �a:1#__+} �}&�X�S�D���	@�4�O�̽OL"�3]նb|DP� ��+�
�[�=]d��c>�?,��}<J1]~n���и�'d`�s����ō*J� �ou8]��1������b��m�U�_�8�x�u^OS�*uw��t���'}w�N���kڹ��|tx!����x7"EiF�bX�&��Y�������x߄,Cu#�:R7pHh��hv�� �r0�G����fx)�Y�}D�y�ǎ6rLҵo���Q3�ó���_���9sʨ-����7lV�"��?6S�}�i��	�Jӣ�m�$�:���������j���!�2%z��U��Òxu�˵x���Z}��߃���E�W!9��_�J>p�d<����<��֩^�Hj�j�@��@�@Y5%`��HG@��o$c�ِA���'��k[���;���$��!�h��'�s���a����$�p"<�D�@���X��-!ib8RX���������0��bE�BZVYH�D�mG���$�R7vѢ5;������x� �};f����}�W�Z�]��0G<]$̢C�������ރ������{�H��yP�-3����!D��w�1%S$>a���t�T��`)�� �U��˺Q�5�̯&a8�:��2�6���q���'���
]�i��o���V*��Ђ���E�.�[�@ٍ��-�o
�2�����]?p�(q����ߗ����5d��S����Si#o|�	Y}���y$��Z$q׃)�{�rkQ����۲�>s�%�?Q%�ė�
��@O�'E�kW�[v�@C
b`��]�Ƕ���w�:';k����IT��I� m�Ug'�hچ����5��3ߪ�|D�U�[A�������[���\�ڂn�綨�����k�0�A�}d�"C�}y����B�fvS��
�4~�lm�&$X�>aS�x�j��GKèoN�h�6M�\})B~ ���ƒ6Y�J�j�_`��1"F�7�	��Hn`	6F8�_Ԝ8��B}�ӧ�^�a���,��&�%�>��)L:�¤f7d'W��Ɍ��}!��o��	c����6K���M|d���S>B-���P0G�����2v�ҭ=�4jSi1�d���W,q�&�dV����q��S�Nvp�I6n��@Cr@�������<Y���"��c4�#FlG�^�A7}�)Y��1z~��ڹR�X�t�Ǣ�λc����ԝ=��W�Y�8�*e�e>~푌 z�R1	��׻)G�P2�ƨ�������N�#��!_�O�x�r�	D��]��Պ��N�%�[k0tAUo���� ��6`�{,���5����`�_�W��}CZ�prݴr��ݭ��q:]�
�� �u�"��S�;o�-X�����_��'B[:��\$9G��
���u�F�x%���Z�}8�-�]00�T�J7v��.FB;�A"=�������zc�����OŦ(��o!�z6.�0"���=py
�J�d���Кjj)�)l2Do����/��FC�HNa���vf*>�Sxe8 �U?��ס���/�#���%�'\П��e��u>Y���W~��I���,����'$��~���qu��O���RWw8c�sZj�^�Ԍw!#e���	�ת���u��՟��?s"�W�jciЭ���YP���[�-fO�й��|�61u���-vт<�B5'z}���t\�@�o�@��U�%��//�[so��+�����$��i���X㚠�C�U�x�U���#��c5цg��7e�ň��&�`U5�<�3��>�p�]("Q����c��Q�E����G�7���Y����Ao�@2�<al]�(���䒖�^1_��'eW��`{i7������|�i(if�MAl��<��˂SZ����(���}�K����bG\pJcG��E������6md�K�����&��uC�yR�B��UJ�#E���M|Z?y��� n��vM!i��3�"�!�}�#��[{��{���
��ە�� O��+����r���+JH	��GT�(Z��ؗ>�U�H���-J�3B29F��ȢyP(���l��L�.5(D�<��/�lT�_�D��įzs�_%!�VƝ����s����{�W�3�TmS�Vz��co���kɦG�խH:���	?'b��|}#��r�y�&�4��^7;p�,��m)8#t��l���kkl��r�ؘ? (�ǋ]��b~prrH������уw�k�Mk��ڻ\p���h��2������O��waG5�HJ�伪)�I<�p�p8���O@	��2��w�l���-�g� n��]��̄g!��&�7>L��fpM}D�4�6�.t�,��K0��-�+�ʼb^/?#>�ʛ)ؿʭ�<��gYx�g"ޫH���F�Z}e�� 6d�ƈӚ8VB��f���ҟ��F���-�h�VM_k9̿DH
��HM��O�i�:����3{$*��޶E�E�'`��9�����Q5h����5T6�AZ~��Z��Y�X8NJ��ѳ����ٮ��ʹ����B��g�o[�Q�#�GY�Q�a��(��u��O�L\�>r�����ٕ�8��"S���������L�_{�c��<�����A�=eb�^}�F'���D~>iM�N�CÉ;�-?$���Ђ,l��+�O|T�bdM ��ԕ������Z^F�(��鷥�$1t%�Ǯ�15�ěo��yoe�	!�j�f�	H�i�%�ڬ�+��yB����wOV���#�o?p씱�+�|ҒH-��G����a���5�w��[>������G�z"S��|߇�`ZYg4d��W�����i2�.��&O��oI�ZU�N����X�h6.Y����$��[�Wn����lKl�aΠi���.���S{�\�Ja_����$��	�ܕ��@��s�
[��o<���l@E���!�դvH��nɸ�>��[?����Kk8{�����lid�9�|a���{���t��c׾Ԧ;��,S�7�48�L� :,�#ټ��71�7��zG����}I~���?�]��ԋ �"t�W��� ������&��ETM�^~�D���c�o��B��3gp������SAh+8��'���wg���7�����B���Sm.�@���Ӣ�c���a��8#m/�-��\�aޫ���\Poy�jۗ2�D�L6��P���N��WW��y�WD���:&OQ�'�C͒%�r����s����۔�i���˯�tp��Ҿ&��>����R�}���p1��h�6���l8f�F�z�q�B�|[ܕ�mG-!����]w�K��G҇����}6���d���ګ=�]_���jN�;��@(�i�2�ۘ&�g<EH���w��2�ËKٕ��S~��Jw�ٕ�!�fE�����G�[H�oe�M'����d\N��q�S�ĵ6u�r-��=mo�V\�yџ�T�N����	;p��#}Hzī�V1��)^�&�� �uwl��0�5��1��VEF�w�l�7������&C�3;3�"$�]��^�&ď�ѮzF>�x#2_$9� �q�\5xWy�@,T|����y/���)����)�Uo�S���,����n?�B�Lu�n�����p�^{�ݰ�PEa�b�"Ta�<��8ʣN�v� ��PԮ�%~QEK;'�ٛ�N(�5�E�������H%>t��c���
�-"*�\%;lONҮ�T�d�΁ O���HM%�IMZ�>�&D��w;Xn�M7�Lт1�v�*��Z���G�K_�N��w1ۋ7�C���2�$Ք�g�0�ͯ����O?��b�kK��-�EO�VJ���̖[ٟ:�F��������#(n���,�� 9|��E]�O�Y4»�89ޙ��Ĵ$b�P� up�E�^��r/ ��|ڶ�%Hp�?�(a-3�֋�3x(Y�Ox��vX�Jg�gN-�R�I$uYצ���t����M-��(k5�����oǖ��6̃��#�?� 6�Ix=�`pI�zUZ~�����~\�6D�l�3��)c�J�Νi\"�t�L^a�M��2Z袰?3���ѩ�<ґ�ƽ$y�0��/9S�M��z�+��J�)o|`�Q��m��I������٘����T��<_��;�u!��g�ɠW�t�[N.��x)�qnn�\�=ZD�_`��}��f��V���s��Wt����yf��(1�-�wu�⫽d���##d�ᠠb4ͲI,-�UmJ̩�>a�lsy!��I��ֻ4��S̭�FD����V��%���4�,�ر��(�j�j����0��R�Z�A����]p���s�#�!՜�:�:�d�[��{͖�g�V&7�P2q��a�L��}���ax�Ǵ#hA@h+D :QL[�"Q���D�Hh��!ar����BOO ��R�B�Mu\I9��N2<���?t~�9��˫��v(��J�gp)0��ٔ{,��~H��o寋.o��^�o@"�����p6��v|�.+I�n�w�jn ت�_��󻰷�u_T
oX#�U�-�R�Q�-VX�)�V�g��xYGxN}�o�����$�?���y� (�f<�0�0�~g7l�Q�2�D{���8<@�P�:]/�a&g}�I+/7��Jy�us7ǣΧL�j��~޼��A��dzҩ�OK�F�HYٽ|�9��Fr!1���m#�W���C�i�5ByY��L3}���}���+c��ǲ��l��
{���/�X�WS���&<��2�Ԏ�|C(���SP#��s1�J���_p��O�׶�l]��g������%G<xE��΂�m�'5k�/,�����NSx��B�͞)�=���5� #sƪɓD���\�
{��l�ոBӂ}(�M�St/�7$V���	����hK�͡�Ac��hM��3���:C�%�@���%O���O.Z@]�/��=�}LZ�Q�n�ٯˑ���V�t���[���9�g�̀5���.)���Q���6�ޫ��`�P����!�9i/+N�~�HX�ٍ��>�¨9��[z �R�]���4O)� I�a�,��o &B���H���ϓ��{��g*�����W䑁b���8/���� bӛ3~
�i�,	`|�s$�2�<��`r.�'u�8��Xw��|	#��lOG�fV��/�Ѡ�� L~I��%ԾOy�!�
S���*i65u�c�l���}��J�LmO.��������)����$g5Kd��$7������""��������i�#�7��?���e|�ʌ�V��@�,��uEU�$�qHo�;��������z�`f7�����@���-�M�a@%�ތ}	��j�CC��7Ov�h��l�l�r���n����LS��(Ω��I9Mѥ02��r}J�[�϶��"�ʍ�d.�D�Ɉ��;�b�������^���]WU=C�EL/��g�w�]yi�:,w�������ژ�`<�����>BN��TL���ʏ�9�%!#q�:�z�py+���4��|�u�/�]�$"\�����.��4S�߾k� Θ�^��p+�r������X�t�5*Ư�r�gDx{P���:l7��%���[���2��6{�Z�3.g.�%VQ{�>��[���s\ж�0A�E��{�vj��i����s��\����/�?���d�o���ߎ3	S�-%���j;%,݇�Ps�O�6Q�l/���>��[�D�ڮ��������;��z���˵�����:Nč�h_�Ќ���#t��$�^��4�s�y��w��]��@9���8�ȜW�[�0U�˝GH��f�|b�}��=V��� �t
�G2]�F�%�#ĈV�yd��E�Q��T�a�E:��J�|���f����N.y��8�J���Q6<?�U�C�>�,"��^KX�m��f4��_��*�N�s��˹J*z�6�D1>d�AzƆ�$��oB}CcNtv)�?(�W��3(�_i�NZ�'��Y�� m��ۉ>��e_b�dh�MLܜ(��n'9y�'qǈ� )@�΄��J�.��`a�q���f	��Z �$}�nxC�yБ<O�.i�N�O��fT*y>:��[�x�.��3x������i�������M�Y�=S;)�	��Sǥ��H]�߸�PR+�êll��������[,��jwrSI���^����B��,���rE������K~`_�=�>g4t0��i��M�~'.T6 ))P��]�Ĵ>���\"��ЉX��.ic'\s�32���>i�� �If?����T���_����0���^����� *�~��[N>�<�Ih���p��I��i�f�6ŋ��;J�$*�O���k�@>%���O��<�q��p��-i����+�CQ����ᙈ�!�����<��-G�F��]���=��{׸�2~�-�vs��;���A'|amLmD�
(����"P�}���dx=h���Ȩ�ԯ�xq%���ή�о�N&]�rC����JM;���-��B�	J>2�!">�˛)�M]��iD;2�krt��޵�.No���a_欄nk������6�Ȃߚ-�^��W �a3���*xR��0���ڬ�����@���&�d�&Ո�p|�׊zc�1�VB�0�S���Y8��k�[��=��'���W ��\�!�'�՗I�,ZW�87���;��8�/%�f�>���N7�)"���|[�����FvJ��̩�s��t�\M"a� F��-�+t�~�:����ǨY|�Ⱦ����p����^��Bh���b�ӕwT��d��}Wo�n���aJ4Yds��u��pv�o�;6�c|�o=�|W_�{k��^��X�C_��8�5��ߝs�w~3Dߣ�I�K%U����k�������d�H单Oc�l&b����_Gn���W~�ƪJǧ��p��φ�v��'P��R㊧�E���q}Z�O��oj)��Ie/tO���X:3
�]��D�MZ�b��i���>E�v�4y5YX���<��}{Y�� ~��
�ӯ�N����[��#xݨ�O��f	͓�7]�	Z�0��>�� �Jr�^�\��٘�c1Q'j��=	�����=&����Ϣl�.��'n���q�s�bf(�,��ud�����/>e�%ŗq���s����{�wϠ��Q�z<�6��1�>KW�q׌D(�X?�ht'sGHz_jK��5v �JQN��P彰�,�OҰ�TQ���$����z�tr���jR�B��TY���&]�A�Tj�g� � +&.�.E���<��?�8��3SΑ�l#	\V�g���-��-���!nO�f��	�W��n%����vĽ�}�G@;�V�}v�d�]�Iֺ��6�G��Y�눕��;ܾ�	��6�XV�����ԭtY��ݷ�ӷ�o[�U_�pFK,�w�7���,.��c��-�rK��;����f�Y�K��B���	̓8��{Gg�@�. v״�?�����������t�W��R� �������C��#�XZ4@ԥH"���>��䤹��:QP8�����}\���5f盒7�BF����;��і��V΂s�#�í��tf�ι�ocu������,�zkH������l�$z�q�~C�/�a��̝�i!�Q����Y+[��7��<V�P����!��؇�m���X-��I�)���I�"ƺ$9�F4,���xhX@��q�l�~�;��K��N�� �bP�
ѳ�up�%Ҳ��Z�͗�X���!�P=� �O��Ƞ��>�U۸���ѡ��l>ϑIX�e��bج$��#�<���c��$��n�M)� 8��5��0Ψ�*E*�N�DQ��.>��tzO�G?!?���	�V�;xk`}:��S`u�p���β�*�R���O��i��
�ycTs|Q04�V�yT���	���3h-A �(��.<�+�f��Y���b57N��h�G��kNX�hxJ�\E"jHZaP���k/#)��*$��#�>����D������qq�t$�S�8�}4h?�\�< 2ڂ�se�(�����U{u����LsLn�@�<YJ|`�B=�Yq2z��y�h�`R�C"�/���|���q�
�[3�1�˧�����E� 	�l3���{,*p�DP��u��h�Aws��49+,�D�_o�~M��=�PX֫�	��4;݉�ޥZN5zڞ93�̯*�fВTI�|��I{!R���$�m�R(�~�I]~�(;�-$���'UK7�$��V�0�xe'���ծ��h��H��_*~9$����6Staz�h3���8|�?�Z\"�~t:�#�%�L�~pGZ jؼ�Ι"9��w����R��P8�W#i4��c8&���@�a����u3C�/��D��2Lm̜�΃�,�Jk�#܋�z�&�ȼ6��H҅U���vV�SQD���O��ψM�]U2`�H���p�?ɾ�v�s:C��'1v�.(�q�42��
X��t~U/}�3�9�sB���VƉ�߾a��xE�|��L�g|�)V�����>��R�E�����7F�ZA�8� �V�w�{��MG~��J��F�5������2VG7#�Ѓ�q��I�Kۗ7�+�Df1��Y)Қ��Ph�$��	Ԫ�kB����2��� ep|'l����n��l�B��Oo��h�6qM��[���yI�pv�v{�gk��Gl�K@�Qy3��O�4��9pG�|�c5����Pu���iP��_��ٓ�,��թ��U:�R�������$G3{�b�k.��x{~�P:7\:n���?Ž�(�d�m
��綟�Mi.+�E��?�gb�G���/��*KI话òZ���#���,��%ބM�Smڊ�3�^�9
���v��R飹����=2��Ŗvs'�(��I��gF������g~d��%�a*p�Ӑ�^�;�bh��%��L��$�4骄�+�|����[�*9�v�>�y��dJg�)��堑�t/�(14��a7M\� zԲ%j��8��4p�0���ͼu^=>�i�4��c���[~�)m�q���KF/־��U[�g���c��b�B�@p��$� �وw��:�V�1 �b/��oM��h>���vp����NS��И�#"Pm�S��^�	
�",�g��2x�p�A%<��s�/e�O��yW�Hw�/��w�?OoA���u���|��=��[ �o��.~	�����x%[O�c���*B�ښ$�MW�ı�5��X7��1����Hl��ݤm{����
;�kf1��s2��&�#�������-N�+s�����37�����O�5m
q��ڨ=SL�*I�I�jp�k(�K�1vA~�$�3�]��������Lb{��eF�����)�y�����G�� n�w��j)Et���= �r�ƛ���/na~p�L5���.����8���~�5��75�?�y�4�x4�������u���T��n��y�7v�̴^�B�Ғ�BDJ-��~m�cL/�˕U.�y����mب.Y*�r�/.<�����G�fM;��p;��
���ƥMX���Hbo��4K�͍�j�q(��)�Ia���E�*��6
�%��\����IC%���6;i��W������w���r2�|��->�n(pα]��+|$�KB�*.��HcߵJ[��ޡ��jw���*���'gk�K?�8��#h��ߪ?��9c��P�$��bL��fw@H�b�{�gi&���<�k��YD���Ž$Q�g�d2���$P1��,IIgW���ܴ.�5��;aq��ݶ����	9��@O*L��ΏD���L�t	LJ���n�ȯ!��%xCQ���Ѭ�.]�β�#+^h����d}M]�� ?R�ĆQ�t0�~��b�a3u�r�U�e	Z������e�]zX��n����b=i9�^�ްe��L�E�I���tяʬ�!&ю<�
&Eqo���?�| c�(�îA�o��7�^>���b)�i ��<�X�I8_~�[�.�J���|��ʠɜ6<��|>�Y���7V�+��َ|T�iV�=z�S�F�����j�T�崛��b+7��~z�F}ىwº$O ,�By��3sj�#V�no/��2��j@�o��fM�S�
�gy^����[�TD�/v�!=���
$أ[�\�H��~uhm>0�N���sj7W��0aH1�	a� 7=4-�;������r^>�����ghx6��Y��k��`A���<R��J=�A}��r�ѳ���!�%�ˏ9�9^�:
���	Na,�Z���J߃^��h_vU���#
}��u�.� b��m�>���4/ v\�d���@ +�%��4B���CK�e>?�����zV֤arQ�����}8����X��،�*��_��)���m���,b� �ȟ�9b^��'cu��E>(�?�ӓ���P1��4�,��yG�շB���y,Hj`��)'�֪��l���Z�e����<��	�ޤ[��a-ӊ&ߵ�w.�$�b�j�Us��Z����@�o��R�����ҵJ>vx��/H9������_̇�5��4i]���u	 =r3���O!Гv�zs���H��~a�r�H�ָ����_hU�bF�Q��f9��,i��,Vi1s��g/B�|��_�6�q�wk�'9�xy�g�\��q�bMq2NuO�ɩ�q��Q���`eT,l@�R���u3-��6<ٓ �\��T\�#����m�RU�RiըZU�v[�vmJ�-Fm"�^EQ�.�{o�7�C{�H�������~�{��=�9�s����}�[y/�����M�%���'���t��'�k-��	��Ա=a7��k�kT}�ۛ~��8�Ƭ�����2v���z�k��eMf��To�f�[m3>,k�c��x��&}��-�0q1ٍVk����Iqo"�CÆ��κET���F��;?���:5(a���������~[6h/��!�Tx���#"Jbt� 3TG|�����0|/�0�SRw<i�<�5�L�uTC��_� �L�̔A����y^%\㝙��ݻ[������Q��������յ�;dSs#�k�J%��q�:\���)·J
���W�AE��|��g�w�4M?�Nm�L�찥��T�9��\���Br��w��/@9���uQq�xV q�Ǽ3ܗK�� ���$�et5�vM#����]�
��oT �4�@6ng���l4c��*z(���W���/+�k��gؓ�]~!��1���'z��8��I�\)xEo��6�w@Q����ގ�}/���)!���8��dP
��H}��~�l�����N#�jT����P���hU��0����V��B���{���aB6t�;���#�D���u�]e@���]�(f[pq�^���4=����&@X\mj����u���S%�*{��{o�Bָ`Gna�ȴw%�ؑ�P��G�6'�mZ5~U!����h�6BdǢKzP��տ�XK 8�{�~�5�����OP�r�������wYq��	�N��k�����zJ�9H7
 qaWZ{|vXs�#tď�F�h��B���֓��A=�����P���]������Y�V����K�M3	��)��Ry�)���J.:���2~Xb!�wk
kE��~�c��_.%QƊ��I1@m�TG-��j�nR`����o3KA�K=}?�z�E�|�Pua��!|%o6Q�U��tUi�G��a�:��I�Gɣ��yU�'?�e�*(��+�f���]��܆'����͓�z�y7��
�,�%z��Isr�Kq�s��(Բ��f�N�����ҷ������I�5g�Q�{]��Y����e��ғp�V�P������ѧjlxe��&����:����"ę��ffODF*|Y�X��`��d"�z|�}�=Ƈ���c lv��՝��G���z9�/|�����4r�w���f�
�L���f6�lLA�X�ڤ1��3R�aٻ�d�ڍ��.�{������C��n�&5ayY/o��� !B�{22��g3D�"���s�Xc�}�$>�@��� ��s{t�������A���&��c"aD�Ҵ�(�HʌM�C����]V���4��w�����Fu����}�؆k��l;>��T�,�S�e�bպ}"08���K��38�{S SB�/_��֬�����E�W�h�#�� �������Y����˴�֊�:�o�w|�5O+��*��~��JU�=<��#��*����)=޹: 8��ý}�4.�q�s왮�?��!��jy�G�"*U��-3�9�Cz��3d��
Z65v��"d򳰫T�͟��	�<���=l#N>�Kz��,�>'1�'���I��aU���g�%"�o�#Q:�#�"5��#�=嘼�9z��qNd��Di������_D�]UCw TS(X]N=E�>.Z}����+��֗��p���a �Z�5��q�t�b��CM1����q&�=�^9�dD�쟂m�|1C�Ǯ�J�a��e-ǫ-�̞������'|9��s�ΰ2�F2������P���mS1;�N��ȕ<���!VU��c�������[~��I����_q��Q[�8�@:#h�:G����������|��C����^C2��iV��<qW�MP��I�붸»M�L�9�ބ��f���]���>�(��e�S�6�d���z��-��c��B�"-�n�3z)�֗Sg���;�d�[�/>'~8{4&@�[��>�[�ҽ�q�pt��I'�N�'�pV��-͚�VT&4F_8*ݱ�à�'KODh��s�70~����j���/Iј6�����g%�&���0�fi��7A<���jZ����<���W��ȭ2�L8S������A�%b�g�'qTH�]V�i&h϶S���/|T(m�����>���ϵ�C4*N٤����u[�y_G�[���l��߻P}�ԅ)Bꌱ�U)z2 ���*V/�f6�����_�&h"�+<�!�Tԏ�j9�3zf���el֜���E�[��ǪՋ��2��t��ج��+W)4��$����<��z�ؚk��rX� �bOO�+'��鏻�O9B�P_rB���Q�-��[L��K�K�����k��4`M���2��嘢aMo�q h��c�l�D������lO�طQ��	z^�xR�ݚ|C��(X!a[��������(
M�(.��.a�Ǆ��Z��5��_!siq��@�x?&��;ɉ�p���L�R�{-�q���|oA��KǤ��Z4\��=Jq���~�G-:�f���G���@얱���q� {��K,^�s��?m��ө��r���X��4�J`�-+^�PT��;������M��O�}�}���!�Ƒb�;���K)���p5�y���3�7���p5��f�K�dKM��k�Z��H�^�rL�շi�v��Z.�bq�w��&GGz[���&O4m�WURyB?�UYi�R�(��m��������x+l�Y��5$ ����ûX.7�������Gtew���&�-#�=�<��#�H�cL���S?����(J�)��j�z翆s��Z��5��)ɧ�n͟��&�Sr�cy�*UW���*�L��p�����e�5��"8�{��I�ޝ9��<�N{��e���S'�}���|�W���^�0�*)ʨZ�̉%ؾ�U�c�{$�xU�BX�z�1��޾t��=+��E=��"���?t�L�8|���=�~�3��i�����L|<sO)��_4��,z�cQ7%?�W�#ł@m�v*(�� J�u�_B��n�E��a;�w�H�:�&	[T�T���z6<J}�8������BSG��<Oi��E�:b��T�z��{�r�@ˡE%\W1{d�9�@���(A>6_�ӆS�������Pg(yi�Oʡ�2S�v�DT^`�%j�ۢ�h�Qg�U�W=_�>��۞�z��6|c4�HZbY|�t88K���.�nEⱗ꺲b�Tͧ������(,�3��Ju��푲�vկ���i����w���	g�d'�����`#2�����m�u�K� �������p9�q<4���Ra��) ����O|�2�ձp����J���ns�*���<�7f=y��e�܈�h���g\4�H�e�--�6`�����ᨴ���ٞ?�Z�V�V\L���QTM_D�M�0����@����H��kigIh�A���!vP����ME��fYb��'`�˟"��ֵЖ���:��rً�ߴ6�V�>40�����]RZ�p�a��;�jZD��t���ӲO۶����vjޤ?���L�-$�H��Iĸd�NJ������Owf��C���f
^�'v��_�+���b�^��p<b����1�{Ty��������'�΢$Q�����E=Z;��]�g�v���/?@�#��w��J�.`U���� ��o~��j՝�kx��*í�fw	�>��x���y��ꤥ��)'V��hy�sHe{/�rb����/�R�4_�K��ՅZ�]0}eH��ep�9JBזϫ�=t�P�r����b�B��v����1�7ǏQ>��J�,S�C0�K?�4b���s��K('�"Q�X抌p�jO�8�#�/a�ގ���&d��Q;���R{K��(�$;q&���$�57�Z�'N}ܳ"0�ּ����E�i���܀�ͼKҶT��|�P?9d�'��ER�EDm��N�;c��O}�No�m')���ި�{��魥�l�YiA������36����wN1��0��P��iv�A�\lf�Ǟ�[�J���ؔ/G�.����'���Ӊ�S�2S��uG���?�6�u�Fmy�	����a�� Gd��q)�ձE
c�"�_/���m\߇��������o?'�܄y� ���s�pi�z��,�u���&�	G�<��k�=�ۤf��])c>���u��/q�/��f�
��<����@��/��q� o1r	gD|�d��X����dm��~Q��&Yu��DZ�t{���ֻ2�8P��V�XW$���\�w��cG@���n�^ր��tC��ܕ���E�^#'�w�Ty�n�g;�h�9�0�2S��8Ʈ�Dv҉r}�\�D��-�6s�_Dv<￷��C*~#�� ��4��x�<ظ�[w�J���Y�� �V�9����I�b�X3�K;s�K]Pp})~K?^w"�����~cA�S���t�0+�,X�sd��-8Gm�v�/� ��-	\���%�g�̤+�6Ʒ+ w7���D(v�1t?���1a�[��Q"F����"��-2c&�̻V�߿�>3�a}-ЛBm���ۭ���"��!g�]�E��f��d�eYMo��H��E����E����9�YU����P1�Xׯ�s2����K�
���{h�J)k���t��>�P��X��G�<'83;<��u��y/��<�$|��	��K����MV.���q���j��k~�>��C�]#T��~֎%hkR����$��s�p_&K��PW 5��"a���i���F��b?^����?0�,e����Dq�J��he���ʾH�
.��])EE�mA�S|e��e�T&V�[G��)�~���@Sו.S�ٲ��>b�Al4�7��+���e��L�n��NO�ڭ�G��Sa�$sL=xfi�C��o������0~��i��9:0�ծ�t?�9:�z�z�����=��HF�0�9{��y���x������w��iH�3o�C��w��K(���[��|ۄL��M��w a����ЂR�j�F��^��k����Iť�L���e�&�Vf�uI܁-��_ƞ��N���qKĊ�#^�_fM>����y�c�©ڧ�?	�Q�HFn��x� jF���wA,~����l�Y+ݴ��%4�B���TY�w�RH��_�I�ʚ]q�4bP�A�P�QL�z�w�! ��V����3י�����߉����uWhN�c��\PZ��^�;g���\Qd��Β��
���-H�eYJD���vwQ��t����Q�.6���O��q�[�mC��r}�r���kd,�f��\Ѽ�Wひ��f�|��6��8~^����R_7�!���ґ-=���p>��uA�����Q�7�T���;Ӭh��#aQ�r k:�E�r���\!����F�-�ܞ5���:��I���m+̈N�*��'���>/?�L!)��r�Iˡ5�a��8�=4<gP�tʮMܝ��+q#��7�T�d �(M�z:�4�����H�*c4f����t��
�Nݟ�#I8ˡ"s9ۀPyE`�Le�d{=���ʁ5ړ:�w��\���>.�0fq�Z8�BFm����#����92j�d�����IL�B ݁�����߻�� L��U��#��l�Ǿ �1��]��̧��)���'.��{�O�]?p��;�}<u7I�+w��8m��.U����}�{TG���ϻ��J�*�9�,�t�qy�ZxN,%���9�҄¤���>G�����%=g3\��pyT�@��B�lyZ���'U����D��w)7Z����������VRė�{@��k�����f��O8�
 exM���RSR�i�۸�1!���^�)���?I�w��o�JM��*��/�]�/����(��RѦ����Jz<��`u��X ��&O�h`6GT���.�d��ޱ�3��Ui�K����V��Ӈy b���ŤV*�FH�Y�q�sP�j�co�ؼ��l���?��\z�&KiP��M�j�b�)vyO9�Ͼ�̑��ɖ3?���
_����ңBO����ߺRm*� �>HQk�-���tEg)_�M��8��!k�=��2�@�l$J�z�vھ�P�=t\AD<	c=zb�?��~Dtbd�)�3�L�O�9y>}���-g*��ï8ӂj@d�H�A�ص }_��x�FoU�����ͅӫhp�Ur�g���N�2���%tTS�LitAj�<v<"e]ms��M�������TFH�#Y��;R�����>xP@�Y��c�;��0N�zdm�ڶR���s-��כ��y�8��%�,�ڕ���r�u/��T�wJ%U�_�B��+0�p�!9|���繀䟴��bvg ͑<�5'�"��?Ns���y!���:�]%�ty�$\�����>��; �Ψ�3�u��s�O&�#&����-�`��os�R���ߒfukS�#n��5E�X��-�^i�/�T͢�����=�E�Y��t]���Ol�Or@��=���k~1E(�/��ׯ�F#7^f'��B�^��� �_${bt�8�i���5�����U��xtJ�1[����A�DNG���f,s+����z���|�MtN��d�E%�E�ʙ���
lcX[�Sir��\�@��΄v]���J��Z�.Uf�]���(�\�X�vL��QrY������{�<�@w��tʔķ���O2��"�Z��&�7Ѭ�l1��F��S�ib�8�	���,��ȧ�)m�d:�)��ֿю���mr�ԪJ�5D�����hA���;�p���(�*J�?O
[�>��)pAˑ5-!dУ�ԛ�E2�|'�f��PD^cqNC���YX`�g�����<K^� Ak�iOߧ�v��*9Ĥ1Nl��lmb΋3%�C��1kzV�F�ӎ�^��ؙ��@�3�����}�6�4ԋD��c�Dce�Y�Q�@�G��R�{�/�t	�5�5[d���߼�^)�q �TX�kŀ�w;�[���7ʯs�,⃶�e�N�v#�pe��	��P�� 3�@{MQ���N��ƌNuo����fP�9�"/꣑���~f�Nr뽉\K�Z�{%���f�b
=2>�V�|b)��q�;��9����?��"Z<�D����[�h�~��J���ݍD��Au��]�2AÃZ�B�o�7��������c���n{9�l3��937�j��.[�N�_�U��v�?Y.˖>�Q����+��|k�����V��bO����>Qқ;�I|�S�@cS��tq������AS<v]N-�E��+�5��q�<���nq�sDk�4Jg�ц��f^�Y�����`��#|K�K�Yj���\�?5�M����q��+;Y~{�۔��$h���� >����E�9�eK�QI�Y7�.���H�ܓ���}�@��Il��e���hH���2�98-vƴߟ�mc��,��}˥r�O�4���o>��I�э2A�鈅ң�
< �G����k�_�q,������ې�[��7ۯ��u]�~���.A�s_GKW�:�W&їƄ��OZܺ.�Wv�X�~���uߍ�H�����/�Ե$��yI�{���@�����|�5��h�"K��K�E�5���z�����i;�Ӕ���#�q�{G��Y����HR�1�-�
3Q1�kB͏��Ț�2���Ws	��G�o�"R���k��1|��j�P!&��:�l�b�)�����^���［��-�gQ�dx�h���ې�����fb�c6:�.ܵ���,�T��.�y�2��!��A���GC�m����R�l��a��<TS�G
�Ym��[��A������["I�~�i׊!E�|�Ğy���U�.��K�۱�p�I�Z��ol�:�4�+7�r$|E6�����o�*�y�!��'����6������o>�I%[_���rׅ��7�q1|v20g����)���ŷ����D��>b�T[�1ϑ�����m�˸_J��b��9k�n	�&0����g�����J�Y�#����ڃ��;�\�Ol��^�a�*� w-3fi�^�4@�5����:�?�"}����+��h�[�Ը��)�(8�VH�cI�8�εѹ߯M��R��)q�v@,yn��|�@��5�h?g2��8?�}��T��2�tU���n�C��Д�!N�4����y�冥k1@�F�;5�٤ZzfG��wJ��o�Ҵ��
���z�gw�U
��Ql�/�5��[jՎ��(L������ޙ����7����ˠ�v��wA�	����fZI�]]O�M� ��v�ڣ[��"���� ���yJ�����NV�X?��?0<F�@�ko�z[z��|p������=Լ�Ϥ'�N�o���7Bc�:��?N1[�{e��k�t���/�Q9�q���Yg����2̰�$��l��pt����ُ��j��+k��e�z�ϗ'����¤GYj|�x~!fl�#��_�j7=�����O|�.'.|}"jZg	�X�O��%�F*YM��@�"���z:e�<x��!�����OZ�<|�����J\���'�jnnP���(��� ������3�sƹ
p�R6UI̹���+?�\�6�B0�v4���d�䪇���͜��%��z�^����4��`��@���ܩ���1���F�\Ub��D�&�Γ��׏�'�O;��f�'�cn��[�����I9����߉L��P9̩�]W"|��1|�Rt��׷��r���[����k�]�����9��wT��_�Hn�w�XW0(l:^�k"#ׯ^��:������G�b�YZWY�j_Y���$��բl���QV+�T �q��;$/_������;n�
�#�_�Q�dW�.��z�Ɛ�Y�H����<��$��-Ƙ�"�K�Q���B���d��/y��04���ؒ��ez��0������xG<��4�F���hՅ'�[uAb��Y�]n����=�]��s����'ډ�0@�'�		;o��<�v��}ql�ߟL�?�8��yOsE/����wVW�/�Ƣ���
�re����y>Y'S��Gz���x��|�$5z��+Ћa,��-sqھ<^���T�aQ�NlNR��?��p�M�����i���4�JU%C��x2�����}��C�׾`�����D3�3l{� "��Ѻ�Ȣ�U��q�o�Gy�F��'.��'�+
)�D�A���ɧ�׬��b��t�jD�v�	U�*�,��ïyM�B,8��F������ ~���	=бO#�2O1�)�����/�:�6���kà{9ZB�~I1j�<�ȕS����̻[w�U�:!ɬ9����Q9_R;�)rR(`-���0�o�R҅\��P�փc�QQ[ʤ��m�E���w��b~�.`�a�d�Tj[qZ�ڧΒ�>�w&j����L��M�d#K��X̍�M\�{�V½oYSL���5�|j��.JW��ݠ�A�F�^f`�?�1Պ�M�]��X-]t�#���9V3ȋB�@'u�i�]�j����'#S��`�Y��ɩq>t���hn����;��g�W��6>P�ͫ�\�� Da�L��d�

LE��MM'��px��:�ŎP�R�VB�}|f�qk�U#U�K"�O�W�{n��I�>�}�Wmay�/� 
�ଝY�(��y�L�.�R�'���_#�.}�Ѓ¢�]�x�����0d^y�4��������\�����AM�/�ԛ���}�m��X�Y���i�T+���EL����Ҝ|��9g%�n����xh��ݓ�t��}�{��%��67����k��嵋z6x���\���˱��r�{Ue�7�L����*��xZ�>dͻ�ޖ3��P.q��Uԗ�X.�F'%g�8��|VB�ؑ,x���b�k��.��}����3�^�d��Q�b� �.� �EOW��zZ[�����JG�8j&6�5�L�C�iU��k�j�Bo#p�m~K�����!�/�ʑ��a����;�MK�`g�Gi�qX�$���oV�����}�_�>�1�3m~���Q�Q���p�7/�����L�Y�.�.E�B��W	g�W^���o8��2������$�.ȭY�˜W�^Jޠ���K#Sr�$ݵ�vuvd�F��hߕޔ>кnt��p��q����= HKZƟ�v��I���>�f��Ag�-��R:�Fų��&_B?Y��@�O�}'22F��kB�b����<SmT���K��bi��5l����/�W-��ɒ,r�p�'��934%�S��#-�<�Pbg��vLo~�l}���K�M|���Y5�Wg����[ 'ªoD����^�k�!��`Ա�uY��!�S�a�E A����/��ބ�\���C���ѕ�ZU�륻��uU�Ni.��e���گ[mu��gߑk��r�	��Do�dF�5���/Δ}$�T�T*��!}&�q���?;a����)~�k�8���aX�v'��C���6:	1|�˺��~��8�vV9%��I��.��L&�h<��^sĆ9��],�D鿠ڣ��z�xf��� ��;,3s��`V�D��G4/6��n��>cD�s��?u��:I5AR=��_�Kz-Q����B�>H6/,�~ȴ��Bn�/7R�k�K��N_�Y.���φ�"�<eeN���	܀9�:�n��
F�̫�������q���n���i����}�lc����j.�M(x����tP�;}e�e��e�=a@� �q]v�u������.a�i�"��_96�HQ�!�c0�=������˾0��$pMa��[���������?ƄW�~Y�w�=�uߧz1�-q�k����e}����R�Z��-�n�EH����t<i�y���5s�lӑ0H�� �+ ��}��WBDj�'f�˩���0���W�0��f��¸H����%1�_,�'�|?�B4�x3pK��!E��kn�s#��?"����z ��6�l�mX�E�����z�E��>F�����ho,޾���K~���Cs��bff��+��abwZ�����v�����(4ʼ�59t�����Mّ���j������Ldh~wV�P>�|��zJ�F��X�`LX4�������c� �}��8�������0'��+�Ed����I��Qb_��]�D^j>
���f������d����w��M��)b�)2<j�_m>0��h��bZ�^�'�(�lۺ`� (�5�K���d�7IQ�(�ʖַp�Y��)T��e���_�^�3�j�Хuҕ����ݞ֜Y-�Y�qk��k&����LK���o񠘫^U�����Xi4�f<U�ɢJ��=�]Ў���wȪ:C�ߝfy�BY��/T(1L��Gw�#�s��V�Ì���N�kId����_�������s֓���9[x��U�S�?��P�G���0ٕ ����C�$$o��@Yz><U�qa(�gq�	a�J�yg���/X�ś�F���	N1
���D�P��N1���>⡐��[Ϟ6?|��q-��A��c$������sԸy�)�6Xt��s�O�P��kAf����p�� Ѕ1�=����ܱE��MD����O�T�>�M7Js]�Zf�t:����*s�"�s+�]$��+ᛃ�׾�
K4}�����
?������e=�7����\�\fhP��E^k�~��ɋ����U���:��!��T7��ioO+M+�L��K�*s��^�bF\���I�y��TF_l.��V1f�����e97�O�	�m�[��q^01�V�ڴ/�ɴ5_��M����r�3��iU��F���V��Y�`B�S~�z,���p�&�[��و_�70�I���' �gvi���w�O�5�=�>���u;�Z�䷻ц�U�WY��ؗO*����M�>}��e�9�����x�+���
a�d*��G��ƌW��L���O�F��X�
�R������]�>j�Ew�������.�*i	a%��bq��;�0TᩋS(놀)=���iSx�J��v)�4�K���f�<p6-w,u�Eq{V���5D�O�r�k�x��%Z����Ù��ž=��v<o���M��©C��{�#{�b���`/�⍰/��Y� �YIo`(*�K���`��;)~$ϥ,�2��vذf��L[s�ǹ��Q��ڀ�\������>��3����p����?���B�H�F��)�M��7 �rwD}'n} 6�����o��fx!┕�E�n��mj_�*�W<Z�\-����D|�¡��e�j���\�.��>�Ȇ���%���ev�LL<W���b�1|�}�zux�,���c!ۤ����(MͲ�Db�W�OZ?@y�����y����35�նx6A���l��SO3�V�+��!2�a��_C�U@d,'Qy}�l^z~�	�ݫ�`�ѳ *5��eL"[=�����5I��C<I-�ħc�Y��z��SY<��[��!�;��[�?�K�ў���k����ص(ܠ&^��a�D�}�.�)xs&Ct칅ʄl���"֙�'�Ѿ�FJعdAz�Z���V�����<G�Ή2!���0�ｲ����&/Bƾ�\�b�/����6�dC�����_���lk7���>�m�ak�G{tJ��Fwn_s�bܼ.�`b�S�;���q~2���G.2a9>�&�x#����&ƣ�Sȁl4��z2�_麏j	⯎WCI�9�._��I��r =L��En�f�p,;��H	h�����>�zBP���K0PK'��P�Ưt�����^&��h
�S3����S[�Rj/�]��8��F؏7�p�r�����4�IV�Gޅ^������v�r�^��|g~���������NS�G{#��О��)�h���y�v�C��ê:��}��[h�5���G��y�=`�x�J�pv�ژp�N�s�`>S.�l���\�n�nS���Z�Utza2&�7W�}^<g�|����XL��*�-�}9��ȀhX`��y,}d��;����/��]3g�������'S�y�g������>�<u!|�������<����
���qБ�@e$�/n�B.w��~А��u^^^�w}j�[b!����$E�޶�sO�f墩o;n�]��l9��K�J�k)7��B)��� ]�EUӦ����5���>(,�EO8x(,Y�,z]5�x����e{�0�|j��>�'�T��(9缨�R�����~��/��f��Ҽ�Mg-Me�S�l��k�;p#@m�����ZR�R8!�n������>���}x�>�R�1�c+�^�Q�=3q�{���C�H��kR��g�� tK@�L���f����:V+�4��U������D�m��r	k�3��W	���ʎm��-�B���ʴ��|x�|�-�e��7ϑ�.�#.~j7xmo���k�Iw���Е⚇ ����yyƹ��ڭ*O�}Y/J��l��gI�.���/�"���q��i"�Үsg���q�N���V!�f6Ưm&��؉^$�օ7�MRf��$$�@���m���M�O-��Q���r�y��)]F�ׅe���,���
mF�#�7������T_7����I�Vq���Y�fUQ���$3z�!��[]EJ����0&�a�`4�El�*פF�iϚp��1�|V.��,�Z�~��⛴C������P�7��G�������ϣ�u�Ā�F+%)�Z[N~���>DOG`�OƜr�0j��ߓ��'�LNg�����K�g�={�73���� )��[���5>'1��="�> a������_^����D�a��I�BXQ�	U]�P%�Nm祤���$0�Q� �t�%�a�Bz��N4�����ܿ�tK�T^� ��q��Y{��>���g���l�[B؄pvK��7�����o~��E�Y��K�>�6ƣ�|@������O8�H��2��ѽ�:�&�W` ~��O@R�WP��W�o
/�-��`������������vƍ��4��cӻ�'���:�;�0W�g��~��ܾ�U����&���b��+�e�n����[�_���]�2B��W���uX-�uz(���!��I�Zlf����u_'�4�e�ٚ�6�b�%�������t׊c�
��1#� �P$�5�j
��L�e�U��7c�QiUOAj�w��3��x�\-/�f|{M,ǧy�*)�_"�܌��P�e���O�%��.ɶ.���<�T�4B���c#�Aމ����R�&B�p�n����W�_.v�_L��k���R�t�����<��8����(�u���捖��<׎�\y�9)������ʷ� B�Q3�����|�_��8>t�A </.�u���|&�5����*G7&��-��h��Za��J�\@v&��m��6�"F��weNH���Ρ~��4��e_�&���w�������}~�3��=#���ކ'o�z;�R�b'�~p�d�~�&���L�F�[��E�g��M;>��4ɴ�Tng�O��ܛC��n�i�[u١ ە��Px͆�H��k���6���^0��~�O3ӏ��|"Q/�t�� ���,V��%�y�,6�z2p^5���I���5�#O�4���������%g#$Ez�3[������f��m�7�nPj���=���jb��w��Tr�I�ݽ�P����,��ۨ,���C�E|���H��D��kF��[�EB�|�v"�Q�+�6*�-z|�?��O)��2��Yg��Cv�~?>&��Q>)�Խ��N�rӶ�7d>�j��H�f�y�T���ix�ZQ��>Uw������UW&(ǜ��(4��x��nqo�܀Oh�
�@0����Ne���?05)�pҞI^��;y�|t��<�N��Om�.���Dd�9�]���
�}�5�繱?�7&��bBP!AF�Q뻵�ܘ�B>�A"�m�)v�ͨ�-��:X�Z��=���H�QhVo�Ĳ�W/$9�LQA+���	��JeI�N��׏<1�8���l�˞H���#a+�s�i�EI_�/�a_wxl�^4zxz�!ܐx^@�ߥ�U����T*�%�:�{S%8U����	)s���e�������~�� 9������F����Є����jw�FP�)�,�O4�<q�z��.��#��������o����Q�=�P�7;PI��<��uqK˨���Ø&񜉄��с��� ͦb?\)k[o�U�1�y�OI�i6f�|����1����@�mLD�y@������f!ԭ9w	�,�}�B��j����=[���/:97
c��(\������ī�i����3#���୯�?�����]5ᡆ�WV�kP[$pdy"����N����v==Cր�]�٭QMpiL����ha���-�,ZzUE6����0K{N~�F�S\�"n����S���t�%�����A��,[L@Ԗ�ov�-�p"2�S��H�>7y��������QJ.�O��8�ꋇ��6�(�&���;���j��RP��zO2DFB_�w���8ɳa�X�Y�n*唤�c��.����S=�7����^�T��Do�k�����"�S�Ś>#h���Zק>���8�A4]EvWx���Hr0�>A��bᄫ���N���uo���a<��{�?�_(�L��T�;*]��I��/���J�M�JO6x��e���11<���"q�'�}4����ͻ�;�M���$q�8�6������Z��R�L��#�hኩ�GyZ%����w��3���_�w����Ǩ��_K��y+ �Ә���~��z��7�U��5 ���G�M���U�D_��~�Gak{Ä	&�Z:<��	A�R���'�?�I�7ij�(�|��)�D�6˸Dw,�ʹ�I��6߃܍�f�M�Ԯ_���}C���8],Z5r�^'�̒����$��	�e�-b1���������H1���υAc�l�BW	5��v��z��*�2�F/���ư��H[�����9t'�/�8���u��.1��Y\FH�;��Ct��g�l�D�ϴE��;y�<k#ˠU�������};ɰ)Pܷ+#3��8��zvQ��oT�$q3�{��Ω�C��g�(8�0f陌d-Xfj� H͸5�W˭���v\�}����a��O� l��6m@��O��/�"�6�_K��w���ơ�v�{[̕R��d�X��ݏ�$��VT�jS�Ϧ�Xɨ�+Kg��������,�>���lc��]�~�Dnf^�9g�@(e1t���-�{���#Y�����3��3vƧ�.���9�'��Z�:�M�H%��(�vJu���ʯ�,��_��]bU
��׍������uk�$z��c� ���S����g�4�;c��Gow(�	�j�@峺ؓ&�2Y���U���m��;����Zkc��Ԅ6F��Ww%����]:ݼEo�mJ���h�=�/�֨�ʻ�~w�㰞�ڣ����Bw ��C��Ǧ���y��	�z`��V��w���(u-�Boy���E�i�̓��s{�;�Ñw��Y����mh(uQ�������e�P޲��ğb�C�i[�]���K�2ӄ I���Q� ^� ,_���QU^����S��B�^���3��^M�ˎ��Ro���2�������d�����ZmU��բ5�Z���ڵkV�Z	� FUQ�R����N"�S�V+Hb�"����_�����r���{�s��s�+Dq�<�]��&=���ˤͻ+&O�u�fߎ��t��<~Z�l2J�<��Ws���_j/$!��G���ޏ�$;�z2�C)�>%�C��O6�Ylwwl�����E���z�N�1V�[E̞�iYi�]`�IИh��f�������/)��%�=뺨r��(�=��ؾm�_ڨc>@etz�y*<B�&A$�=�h;�P{G)�d]�����3\}Z�P�}4��)U �^��+G/{���c�[�6-���c����k�����霼���\FZE(�⏍�Y�QZ[�. �H�k<�W�͸�]IS�!"W�R��uq�����9:�P$�e~��|9)Ǐ4��\C�"6�vI�u��|���p=[���p	(CN����"�v�Q�T�T)�����|�#����F> ʙB
\���tfI����ޟ;�T~�z�)�������lݏeA �/�ڵ�Il��p�RP�[��N~n�U��=u|c�+��M���*��`+���%3�U��`���!��3и����'�%����<m�X��L��YZ�\ ���ʇ��5���9A�9���#���`�Ѹ=��E���@v�KЈO�H(i[j���=�8�3w�h��R�����t�H2����gh���GN�d�y>݀cD\��߬�������M~�Ï��	�e3�	MQ#� �I�2�<�(��1 �n�rUsW��^�4�/�rh�2�v�$"^I��,�Q���މ��؎]�I5���O��D��w�����9�$d�̎Ӱ�DX`>���u��XŖ�˲�
�]~�d� {�t�N������n�����v?�`���N{㟿2]��[�u����n�C�E8�NA�p��јO��kևujq�����w�H�b4ؾ2Ρ:8�n�p�۬2����A��ߪ����,���~���;�f]�{{��؅Q��ѠK_>۰����U^`����6z4����/�<��r�Ń���ScSk�G�Mv�ɣp���KW�~�_ȿHzx��,
�JH�A�@����5�S��$\�rUW�J��X����[%�e���p������".@��}0mh�q��'�WNo�el�r6�Ut)�l�|7�Q�Qy>U��:U�P;�����Y�_U)�$v��*���+��� �@�� b}"�Z�T6�?z�;0w�LS [��?U�f���X	�y������q%�"�_�����jQ��W	m�kk�P'�:��=��eg[������5��%���]~˽��QF0��[���gE+�?�΅9B��C��3|�J�-�J{r�=1�b/ǜF��K2'zl��g�[�����zU�������x��NX	���O�;Q����/��F�U����{|��j�X8�kq�P3��bq���RY�h��i�Y��;H�;�)�f��j�ɒ</��=�Ĳ%�j|��$<p�p�� �o?��T�~'�Þ2^��l��@�@f_����Lץx���l
Ʋ���7��+���1=��]<��TX��q��ĵ�7�߷/uc*�[27�8��{�;���S�B\
d_�_�\�<��=mXk�1=7FV��즒O���L�2��[y.p��=ގN�ܕͿP 7�M���
�Vlie�D�2�W,�V�m� ��TrBŦ��N���S�'ܲ/@�z{B����-��П�+�H;�c�eG�����bf�%T�����t~zwӰѢ���Nf��wㄗ��v����|V�x��[�a@CXIOT��~�K;���;��ˤ��4.r	�+:Z![}I�����']�&�}7�k}�I�3�K���B9����]����+v�
^�K���,�M�jR��/���
��/��4b�����D��Ѵ��~���?�K�$Ī����A�V=��cb�ۧ���\l!pd����L��48��~X�"�>��a%���n�+�c*x�r�>������*���߅>�c�8�6k93ih��V�e{r�^�W�Ґ�*m��[�?Mr�����i�K���K}</��1z�}��}뼬���];�u$����W K�ru3�������b�cs݊�)7kP��*�e� ����!d��0��M�����+�wD�B��E����R�:�a��n�a���<��)Fլ����!Ƕ�R�zL���ɀN�@w���d-��1Á�uM6\o�,Lվ ß;=�����I~��˻n���K>3��G%�z&w��߼���Op�nO>�8}%��+j��W���t�ZSo����+����"�#�o������_�Oʼ�T�����sv/�
��0�M:���v59;d�R` ,]����}�A0��V6t?g�H��.?
b�^!�z�t'�n�����xt1*�@�l���Բ�����Ti���ۣF�7��%����2ʿu�β#��.zgO|qw*�3	���pX��w�ع�|.��|�{�ԗ|�����]A�L!�
�7%j{(rTh>1t��[�)�t��C� �����g��U�1+hw~�:m�� isb�]��z����������9Vwn_i˯<����4��I�%D���`�&�������S�UgoR ����>�_#>vr/6���\x1�yh4�_��5հ�]��0.�#�����_׉�H���mۗ���6�	̇���&{@��Q�O$]��z�Uh�|�Kt����[֭�j�UO:�-���C�e�d����'��6n���Y9�������+T!�o���h�����)ִ�y��/ar�hT�tFf��'M����.n"Zu����������j�����1%��0n(�KE����[��ш:/���Z�5�Z��B����J	r;�~����V1wZ�?��!����!��3s��z�l^��YA���K|P��:O��j=��Տ,YF�ypr�(6�b;�z��Hw�5�.�|�'hR�Z0$!�ʣ�{�~����~M�N��2WY��ڸN�d�T�Y�GN�Z6���Nu�����ˎ�ɲ��W�T�p#���9=�ڤkH	�p���nu�WRr�QS���w��b��5��@=`�_�DFF��?s��=�4:���F�8�A!�e�߹���o*�
���\�h,�&��q��"&$��Ȩ&�jW����"�r�f"����ME����o�VT7M�6X.�ny5?��/��M��)E)��
���0��?V��}M�>�ۼ6b�v;�8I̙%���[�U�s4Ռ��7Ҕ��F��|�n�UF�]E ��]���鍥1��ӄ���(O�����鲵�����y�G�P�%�r���2�Sӧ��ɝ{ʾc�>(���� l&`�̥3&˗��#t����nH+���ef�"̣�؇%�c�ء�=Q����}i^���~��n�b�ڿ�>ק&�C��biP��ָc����a�ޞ�;&���Xp�I���^t�n��S
Jb(l<OE�^�_m�_&e��5p����Q��\��L���c��gָ��i7u'-�$��Ն�"/�W�6d��!Z�D"��Շ��?��4��f�>��,�f^ �H��T��������٨���w�M��e��x�I�<W��n�h���#�tMm�9�}�5�K3k��6����2c���q�*e/8���h��^�(�|C[V�)W<�����f%QK|�Q2(�^��d.k�ػ�MIf�:�Nn�;T1�O\*�����B���v��,Q[�@�}e�Ax�>�=�t��cV�x��R�D������=�W�������`=� �!�܍8�'�@l�D2�J:���Վ+���G�؞G���R�-�g�R�8�o'��V�Rt��Ͻ��Q�H�UޕCU�P �^�v�$-�;�:��&;��=|�D^�8� -F�����n9�W�(POd��udy��N���l�w�`���/p����̸P�\�8��a������2�W�8������{6�~��(� ��\�L_~ҡd�5|@*�	�*b����ԯޫv�۰�ꮗ������0N�p:HͤWI8�� ڥp�Y�Yn#��i0l�
�l��{�WN�l���.��/sl�{_V'}��3#�+%�NT� ���R���Ŕ�$��%h�V��&��@�4_|��~w3A�K�`0~:�;1�wd��d�9n�1Ujy����W�T����*�_���t���	���%ձ0�9����_��u�݇��ۧV�PW��&7���'���}���7�R�n��N�)���Qd��s�;��?��w0�ܳ9�k�*�QEX�����.X\�'�H��[��č�'�K>l["�z
�����L�E3�=�+:�"��
�N5�Jӣ�̤jS�X��z�fvjE��_t����9�m!�^�\����d���A !CmygO?���v��	����b_RY@�&@��mng5��^�ۺ� 	��=�#F^�̚!J"lo�yp�Қ^�� �n�9:/���췦#0��}�_C(l49�7z4�7k���SGG 7�Df�I)���A����M�����"�;S��S�O���Q֖л�l:�����PL
�}|��DUs?�����uy�OeD/��kOf�ˬ�r-����F�6ۘ1]&�z���e<��{Օ&������ܪ�[�+5K�}>�c*@�I\�Ito���<K����^��_p-.�~�"m�t���Ö�a�s5u��j�6R#�u� �5��:ӳFWA^��~slZ�{'%��x�D4�����4o�׏�7�ґ,�Yd�̥� �|?˪omؑ�x�+u>�%}`4�����6*�E=�~�F����r���r{>�O�ɸ��p�/S�M
ݰ��"�V�&���e�h�XH��$�CJp�3��@�	�ec����_���`�'�a��9�'��~ߩ �(���.w�W��+�\�
�a����N��mU�xד��U�`|�2���&�u	�G?,���Wԅ'4lz���4.��V!�������UA
נ���U�f�BzL�4����������=E��޳]R2�!T�mk(,�Y�y� ��4_�������u@D!�4�"~,T�x���@�a�R�<I �����kZQB=��LG�T@�dڼ��M����y�
�UNT~�@r��˥�W�z��嗣`HrK_~�!�<�UpZm�]���0�(�5_��dD0j��f��qeO�Wq�S�-cZ�������2S=J[H5I�wg�{����݇�t4��_��'��F�C����q���{��!��78.����QlJ��I���O�Q>7��3I-8��6�+\�0X�ީ� 7�����.�⥺�N����Թ��� ��F�g���S[xq��;��3]��`����8_��� ��Ȧ�
�kΡk�K^�|�TNQ#i��]f�7��hh��Y��;�>��X�sC��7�~��:����㡼wt�.w�G=6���δ����̶�'v|q<�������)4�)�1&sU>��V6��;��z�;���ut�`fSBF]+��ⴀ��>,ό�)�r|-q[��ӗ���
d�Z/��5X����*���1ZΠV��f��5�R�*�f�MS*�˱չضQ2��@~��=�[��nv��܆�b��n��<�/���9Gq0�+1�n�X��aAh,�ڄ?C��v�)��N4{�e��?�Q�[��+��n��D�v����k�?k~ࠎ��2�=��A�w@Ew ������<��J��o�ןQ�]�7dg-^o�t}]&���������+R�󩕖
�yk�y����4=!<��ia�F�1���n�i]��a� ���7L�)�Y�b�V��n5�D���w74O�7�y�m�D��ˇu��/���?Ny(�����V�m��Q]�U�i��߹Q�?���|)i�-G�1�"�*�žSux���Ygab�[��]�	��@����c)\F��u�'z�Rq~O���4��Z��r����t2]�dI���f�'�����Y�_Rc��qߤ��,�w�1Ήk;k�3�"���J]�WOM�\\����FNߛxk3��;f�ϊ��Y����D��Ԕ���Z��PklOw��[��c��P�ά4�+�F�=�R���F[@�����\[�?k1AD���4عh#a�|�K!K>4��5ZT>.�\l���8�a?�`H6�NA�1�����P�����	Hsn����i�L.�W��9���	i$O�5C,i�'=Uf��ަ��p�x��\GW��l�q8����u����/B;�Ӭ�Y��	�6�0ЀY	�H���������1��e,�KNs��lw���X`r��ՅH�6鈆�n�Uf�A}��$7@���O\:z��+<0H�+]��J�h��U�"�ɶ�� �����9G�yF������90U��!���<I���\z@>������ ��;cZxN���,2o5aJN�p�yp5s}ǉ:���MA��:�C�eb\�
~�&h(%-��e-�"R
il���ղ� |a���|�G�tw�<�1����@�r�}�$�Oԃ�[̰��Wi63! �-�6�<����#��:�%��a5r.�9����R�hn4^O޺8E;��R�%�Q2_�ҧ�����_$�$(Gq�p�'C�ni�wO�2Ms]�ΈK2}�o'�_�����@�k�G~�W>��c�s�7�K���� d;���w�s4쫵v�b�b�4�,C����0����P}�*@f\��vUO����^�Mَ�hpy���[vwm�ӫ�X+$��'9n��a�c���u���D6D;o�~�"Ky5�;�#���n�D1��|q���C�?�N˦�6������I*՝��7{��������:Q2�^;���SB֪H��(ݞ���|(��y6aa:�����`sO\
����K�� ��o�Xz�Y{��O�or3����|}��Z!�����?Gz4�V �V��c�O.�ȥVcll\�шa�j�7'������|<�W�Ƅ���O�J��L��;���>x����4Oo���*�Wt�Ҏ��?Kڢ���D�&rS����iņ�:��H��	i�O�)U8��\�6����������[�Z��tڜ[J"��vjE5����iMf���XJ�{�����TT����l(���b\�"4^f�a<�n�S�òXA�6W�����u(����=(7Q�z�̋�<C�dU~)�/�e}�_'ц�=cxE��3�&IPh�R�_Yi�}��Ӥ@����+Ѹ-��E�DtrV�"�bA�(c�M
��iu�oP��Y�zE�#�I�?ɧ臺���EYM��ǏP�kS^%w[E'���h͖t���2�>���Q�F�χ�r��I�'�J	z�(���ׇS=(�m֗�IPw˺�ݘ�O�e�!ɫ Al�I���v��N�s�`0�<�@�u�e��1��}�gyr�w@:��Q��3pe���^{�Z�9���������-���P;��pL����NƎj���wN!9��w�#(lɌu>o�>,L�G�����_H&�����������R�߮�1ߨ
I���f���D}=��n�V&�#��c��n�9�"K�(����b� $�`z�b���կVf9�tr����;ƒ����LM����GP.U�=7�$Z�WWv�F�т��L�d~�hn��7�l��%��w,���u�%�����'����lX!�#_s���nn�EB�mxngHlu+ڔKu�\,yN7��BH7�E��S��4���<Wʲ[+l(����.i���gڭ�� ��&�}��Գ�Sudb��ͽ8[�r" H]5�h�=�$ lXߑ�N����'ms����¶O p�| c���h5~Rv� V-G_�9J���/��Tђ�6wo�u�vn�3���(� ����k���ad����}6��*.�-��-���?�/Q�1��(�Ŵ�=�طH��,�1�~k�����J�Y� F�M��L[a��+-|�+g	��X������k%��5��Յۮ��{�)~?6�����Yk��9?�B����{4h�q�Ğ���������`B�rO�(Їn�@Η�d'��x����b�D����*0j�yy��ԣ���[S�k(�ڪ�_�
R�r�蕣q=~Z��r-�ͣ�rZ�����8C,��׾�����Tk��
��w�|�	!��T����Y�(�c�fH��ʕ�8r����K��5{U��(�m��w�3B L�pkm���妶�Q�ۮ$��i=�n6��CP����:4�F�U�����CCm�ʨ6���;m!�6c�=��v�b�-���_ݟ7d���'M'�6�U��ԙ$��f#j3�:7�H�7�v�2��=��?ޤ{N/j���xk���0K��������,d@��sbh��F>�����n����ʢK�\������77�{B�J�/����_�%�����Aa �ғ|�S�$��E��vH�
�.Ǟ୅#27'E���ބ�����27�)Z���&�@��d��`8�e8�'��x�5z�n�JX`��S�b�-���VXt 3r�5�"���p�"&2�~��E�d�<�^~�9��kv��f�23�m2\�:�%�~୅�� ��$���qO�}�jK6!�.0�(ό4��Mr(��A� ������&��`���`�ds;!*��eM[�5�,8�7�_j�Z;g��ܜ��f���"���@s��<|�����%;�0-�k�mY�P�4.Px�+��1(��FyE[���ԉ7�f��ѫ �_짱���sn;q�/k���y�	�#�h�z���uIQ��D�]�ji/�"Ѹ�xT{�[f%2d�6+�Z%zs�퍑ai�HI��*��2Y��}�n�^T��A�#nRm.��0yV� ���X��p�X?���:Y�*�8�/$�;}i[�$��}i�O��G��.q̀E?!��v������X�q�%���/<!�����yAĢז���=Fy��ڏ9 @��F9�jF��'�(���ԁ����{\5^t���E�刄�opk��Yz��;GEir�m�I	�<M�K��7P���1�T}�{��%��p�䭻Cw�;�?���劸vw��'���X��ۿ,��1�"�o�ǋ��l=��r�,�?�Mǉ_��Exĝ�+K���; N%kf�{���[E��t�b|���B��2���	BA)lza ��w`�����<�����X������v8��i��A���;�4��/3�
l��Lz36|#C:*�xIJ�,$�����c�H/A(x<�`��\j���b���󚜱,�6i?Z���Wq^��c�I�5E�̐�E�Y�U��Wvz�b'	{<��y��UKO;�%��]iH���slR�N���jY}�
��[Qhqz���p��E"�����CRkKw��\C�)K`�2��n����/S=����x���Hi0,�����N�����/�<�P�ke� �2���^K�-2n�	��SLg���sWfJ ��G���CA�+�x�A�0��pqu�U��^�P"��f��j��LK�r�'2��1���F����5� k��Ý
a4�5u�$�Z���'Ĺ|��^4�a��!S���I������ꅗ�xV�kz仝H	�8�7E��g�/WV�ퟒ��ў�̗���"@Tm/C>�-c��~H�;��
=��"q��so��P�-�+}L�r� W*��A�����g�{M�A8|`�b]���A��R�,=�|��6w�����_�.A#Xؠ�_T����YHQlD���j�h|�ty����x�mZ�D�W���'��S��C>O��&��"�#��҃۞$5��&�?��l`A5�g�7pm)�ό���6y���]�fN�#T�1p�%3�(,9����zp���Ox���>gRxX��x��06�T����s���w�s-�UF��a0�y���&�vbD�u\�?��`�#uB�iCQ��8.%I\�jS�}E�����z;[ž��%�w-��xa;k�!\�TJ`��$3NbJVN�WZ� <B ]`/����AI���>�^x矾-�z�T�?5�{�<>;��k x���e�����AĨ��*)�s^C��10mP����������%�U�_�ݽ��x�N�_�Ұ_1��G���`�����@���O�I��&��͊��+� �,�VR_y���
2��R���h�j�.c�a�b���7l?��ʗ5��R~;��]�wz^���G��L~Bv�f{g	e����w�����*���2E|��S�dR�18��(��=��n���L6BQf�R�TJ�>�`�M�i����|��!	�P���/�0�B\C�B+-jӌ#�G�`��r9�J]�p�ڞ����[-'M=�"���#̸��U=!x����9�ap�x�������J9�@=��b�+fd����#"�z��̙����2�gD�5f�\�}צv��X�����U;UF���.�07��Wί,���<[]'4���yT\$y�r�G1���h!a�ݝ�?�>���7ގ��1?D��Xj�QS�I��/혚��i�����8�|��L>���-��t�Q�r-��}��qXCQ�ˋ( O�Z5nb��狠��;��O�X�f������tS�y��V���"�������pH�~Wm� ~.�c(��- �ȯHa:�����f��fÆ�J,֭�ԯ<�I�eε��sۼ*�e�k&��d�ں�B��'d�Y����"!+dy\疃6#u��
��5���L��#�Z���A�L��+����v�,�8�]�3�,z-��|]�OF�i(B�u)b��tu}��O7�u��؇� ֬�#��]o� 3�%��;�@̄ol4/.���G5���(7��4mc��HW�FI�8K��=���_#͞���E�]׎!�)��,ZJTZKT��Ϻ�>���Ce*~�fQ�2m��/u2m���aԉ�}w�H������AR�>��M���� �iL�*�iWS��>Ų�{��|
r�������������Du �7[Ļ�Ŀ7"@��,�|�i�9��u���� 
7p]�̫0��B.i�z��[��ޱ���Yկ����0��D�>?����]��*��#�p:x�WUS}��|V!��N��8�l\�q���&�$i���c������-��}�"��P�_��g+D���Vw���^Lj�s��,FM�_�F�<����'��7H��M}j|�K3�����DI�[���eї��oc�;=��#B��yj�1�hW �<�4�c)`	�Ӹ﬽���ܖS��ӷ/=�_�*A���th�"/���_)kn@]���Ρ�j�� ޢv������{<��+��9�??P�=8���8�~y����VG���n�^ش]����7���qw�6|'�f���H	�7v�fl�m����1��+�ƴ��%�\(G�d[@�_�7]$I���Iй��$�*�?7��?)d�K��������(&&���+���q���r�`9�M��0�geHԿ��H���98�(q�ةX���Nۛ��p�c-m�	�aE�m����%L��7��j���g�J�H?�,;�1�DѻU~}׏��f�RQb.� ���|���u��o�n�����3�a�"OO���j7����%����c�ҧ����-p�今^|�N�������2���r�4�3��{��׎<<��=��o:bŞ�׊�*�~��p�)�K�~�It�W�D��;�l{�!��=��i3��Y�p���E(�	�U�Ӈ$FM�ۮ�F�q<�`	-`9��u��{"��a��m<l!����;+)�:�QIDCL�#�D뷳O���UŞ�W�n<7rO8�c�
�}eߟ���1(��ښ{�i�����.�_���p��%-Ѷ���s��Ie�D:Ŏ����++�y�9]��W� SQ��~M"I�>��Ŀ�8�Z�I�AW����>��ܦ;�)TW1XE�Hl�X{vtd56إlo4�V���/Gܞ��6�&9��yӴ�g>��r�+�b.h�$��t�/�ݥ}i�
F��9�?�G�##-}���5C�E�Îvb�t-�N���/џ�|��ʑ�:�)RL�1xzkT��ĝơ%0']H~��v ����_�ؿr͂D�U1��D�S?�`�t�9��t�cK�N a������ �N�"�Q^�3����|�g�ԇh�}n�y�ˑ1V������ٜ�d�q��V,.C�lt�4@�������;b��oSi?�8��\��Άx��-_@>5K���U���f��v�����MW�D�� ����Ӎ�hz�x>'+�%Jm�su*~h.aG����2������_����0�=s�>8!9^|D� �V�6����l|�9c��+_�}�a���Tͫ����&��֑���ˌާ��w�Mz���j!r���"�3]�[>&�?^�ʧ��hن�pY�ͯË�=5`��$���K(��!�WH���9�OT�t��ь�*O"�f�`7��;�;�T�#N����T� ^�{j�?���%�hX<��;�%{���A��:�Tmk ߴw��^��e� >�?��&;g��� ���U
\��P�C�!�:��c����5�P�8��cڲ����h�Ӈ�`+��y���]W";��n�����Ԙ�F�����J�PY�
��|vvg���b"/N�ӧ�B�k�����2	ߨ7O����>�N�7��W�tnQ#���p��:��C��Q��Ϣ�Nw�C��X�'�ֵ�\d�Y�{�$�w���}*c���_m�N̓�"0~��1�sX�Q�^$f��L���\��dk��Q�<������$gd����޳���I�]}�=��S���f���k;��5����"c([2���y��"ޘe[Ti�n ǚ<�ä�����ݟ-u�Z'����ٝ�Χ���*ߖ��,T����Ut��w�v�9�-�w��z^�2-��g3�;�c>�ߛ[$�-��Κ.�tۮ0^��^=O2L�Ů۹Л���A�d.:i����[@�����L=�8��Y����1 �Z�X�8�M���F�����E�rRa$�k��r�;/@�C�&���>,W[���i�l��e�=��?�b��(��Ұn6��-5B"��\0���e�z�L, ���A���|8��y|�:�G�E�Kn^x�U�(��5�d�Z��C���ߋ������6�1����������.W�0�d2[��<�E`���Hn�y`~����yBvw'��P
&mwP^�3T2d�w.���Y��f��zE�E�r��yf#	��.�A|�SG�\������n=�C'�m�ç��+��>��25�����'v��������z"�i2���b.X83`�����v�nKFd>�9�X�%^�Q2� �ᷗǯ�
�{-f� dԯ�X�sKv�G^&�6�����2!�U!�3(��A��Y���g!!O�΂b��qeqK��?��1�2?�-ɢM��1kKc���r����8Il��N�A��_��<�w�L��Z�΍)��M��VߤEw�#x�ou��[b���#���h��?����76/`�g.�Qo�k��"���������g:Gbko��}Њ�y��3v�6�g�5�iwC�ycu��ĵ�ya�_N	�%�nX��U��Ix�Ѥ���c�K��HLA�1m�4���Dl=��i�Z��S��yq���[xa!��h�&~�����&07���g�;�eL�7$AFt����w�Tp�6�S����x�7`W,hk��P�P6d�eg�c�wƜX����{�������j��#�g�.�N*��y�#�_�r8�� Ҳkq������y~��jcWu������B��[�R����wty�`���!K\�
��`UNo���{�,А"'�o�]/_C���
����lR�U}d?�;�?���941�G(\���4|�������n�B���g��y;�Lrٌek��e7�Jts'�9ρ�a��>K 
ʙ���L�M�m���Wz����~yO�� ���31f� .��yg���	��HO��s�Y	�U��x�_E���7Q*���ݪ�66��{Hd]����_PI�*y�%L�r'���8.S��AYa��䣩޾�7��� C��"���M�����I�濸����3�v�C5��(g�Q�����4��gȕ�����������`&��VZ��r��'P��ښN>c	e���Ƶ�188K�����=�(Z� c����3eA���g���w&�|�50���Y� %h.14��F���~?�TM�x��{�ݳ�&��v���@ؐic2��Co��4-@k�y2m�77�IJ�hm�0c�Z綖�xB �xB(�;<��6ٚ\���
�K�B��fq�N̩���"��f�ij��;n!��
�y�d��W�ɸ�&����$c�)~�5�\lS��9��~��k�;#Ա��!p�,�ߗ?��}wBy5�`nā���
���"�V4:��E�kZЉ$����H���ѭC������ɹ;�Te�4/C��;ML�T]�����q�1f�'�omP�=�%X\Y�n��C��cV�!�Y���8qG���@:�,�,)4�\i�2�~��0|�~z�B�3�=maX��^�R؏1�I�����1,�-�Y`�e�;�-K��6��,�4у�̸_��ְ\H�����73�wj�b6�t.Qx�v��1���|{�K�m5�q4p�~HH��歋�0D�'�z0�����s�]h�Ȓ���E�� ��:(�ܧ4��]�,���J�)�d����<�AQ�j|�0���VJ�=duX�����I�}xI(x���`?8+,�s��*�?#�q��G�:�dwԻc:R a�K6���zy�D���9;����^0�3���,�����W�������{u� ��/n��.3aO�\�"R�R������*�����;jj��q�����z�'���~�Zn9Yg�`by���H�ױ���H��^�1����q���3�tyt���ܤpz�$��GI���殧;b��y�^5>�h�+P#b<cW�?h�?ք0~ 7�i!?��s��h+_fNw��H�4�r�j���qAD�/�O][W����F�����+~�tYp�9�xp��׶H�|=M����tQ����JMAF\[�K�\����%�(2�Q=��jm�8�e	��T�Q�έr�7�w�4�,#��c�J>4�*�'M
_����h��+�j|^}3E����­Ք�2j���Qk�W�9RJvz�y1�v*�	�`��{�#����s�Z��d�Ə�l�����-�²�q��ۭ>�$K�����&/s~��ϸ-�T7��a�"��rU��G�o�����_#H��1�/6}�vA��w�/ߞ9��ví�n|�%v�Dp�OO�XͲf�s�f�@�@�x�n�Y ��3Άo.I�q�%?s��U�=V��пw��5��V�,�]�q��VK�I�0t� �N��TԼj#�z��ۛg��$
h�4
 .>��V��glt��K`EMj��'��W{� �%��x�� ��R��r��13Jv�+�z�fe"���G>qy�?�T���4���X/�.+��ױl��*���h@�_�=������x]�R�P���cTs1�F�ɲ�k�z.@�B���`9:3���
#��u�[c�l!k�}��ZJ�6����!pC�c����7��EQCdX��lj[6�K������lY<��9'���fV>�i���o�)G��D�5�C;�o�����G��>^$�i�����Ûy��?mB��%�7��eh�|�Go�TI,��׫óc 0�f��������Y������=�&3�YF��D,dQ�W����n�U{W`<����CT>��R��)&/�ۤ-�t�h��]V�g㊍0���vg�x���H�I��W�_�aH(`?}+�g�ӥ�{qj�<EE�D��Z�e��goٺ[ş�a&Ӕ��,e�۞>�;�Q+/�Ν�U�G��ܲ5#�����M��e ��������n*mgؠ�T39�%�C� ���> u��N���N���x��Bp�q/4�ú{�����P|�M��b����yr�����v>r�j���^�t��*Y,�u�d$�a(A�Z�X9�s�<Xt8F�������<���(,pH�k�z<���L=�e1z�HVa�$'(�Y�N]�5��@4������ˤI�rX�:�w$.72$�-4�h|�s�Tk�N=�wOL;h��N�&��N�=\\�,���:Y6�j���ɥBY���ٺ� �׿}\�Wi��%Ϩi�i�*ü��'�ú�k�ǌ��mT�B�/�I�1�ύ5���=�7Pw�v��'���֮�w�Yp��8�3K���9V�Km�S7q�A-�+c���)R�����dٵ��g��Vg�8��q/@Փ�ZE��2Τm��ٔ��X}�kL�a_��i,���o��B�md?ѣl%�j	�� C~o@N��P�Nj�k��gn��������a7�[p>�\ �d��X��`u�,�����f���J��O�6��s5��s#��h����:���x����7��.�0>
����z���]���D��u/�]D��䓲��v�c� �����>g�'.������_מ�:���}�'z�ω���$�M�����T�d�=�'j�q'�:�?���|Y��,�*;l�}M�V1�@���`�e��2�+�"+L[OO�����~��8b�� �U��������J�:B��B�!�J9�"1�!1g��9���C�P9��36�D�q�4��|�m�3~���|���}_�u=�}?���:���r.��h�H���u�?([��:�i|皚_��̙�5Jo�,V]�O�Ԟ���G5P����,����q�V�����������=!��N~��L�O�ǖh8J��n��)��_O�~ù3�!JГ�wy�v��ST�mͳ*�S�̀�:��3*F�G��E�D�)�Dw���N��]�|�����̯w,fqQ��mw��
�Z&��sw������>G������n���^����*C��b0?��S�x(K�tZ*y(�X�ɍ�'�vKN�t=�N����|ju�4�v�J�׼�]��Y��_2�)>}�u�칦��̪Cq^Ý�5]����~&� �nz궤��Դ0�p#��ZѮ�6\�OOĞxv��Z�q�z��%��K��t�28Xt�W�pJ��锳簿�����R�/�Tl�:��s��|�n�~�[�-����[�ŝD��~0������l���w�; B��j�g-iA\>[�z�H����|G �5��q��^6�ƛq��q�)$2��5�r+KG��c�+*Ed�2=��fI^����~��%8�RR�/!��xb;���0���V5~p|�^��,���89	�����]�p�Oy�lפ7����@���8 ��cf^N��oYI\���4��tkޡ�w/�
گ��S�>}��Yġ�j�����K�g��/�gx�uD>0G���Jͷ�WF�2*��"M���B����v�L,���bs�)��?F�ڭ�kf����yH�����L7���C���R_�yg����?���TJ��&i��Z�|D�|��E���:��Hv�¤��0�v_��|�N�^ԩKTQ���%OK�H�x��$���[SUx"�zZ�ܿ�N
竒�u���0��| ��9t#�����2D��YMl\�"&#\��/v�ԕ�3w>�x��.����ԍD����.����w3R[�,i�CjW� ��[yT��jD�,[�H����;d�EPc�L7�ז0�
�Vdl�s �K3�.�dձDX���X?�H�]�N�,t�Cd�[�����"���W�;P��/��(��.�Q՘�ؖ ����*������w�*�^���}��hޅ��>���G���w�C����]4���+kz	��R�pvn�9��XH��~�\zwSC��pT�ş8S;$�V��zc�@t������?8���{�4�v2c�[.V�aI0��\h��~l�DDخ�T�%1��ދ�&�Ş�v3j�JJ�R�<v�;�׏�)7؁\�1O\sa��T������_�:�U(@��<+�,j����sȌ��/L+]�sxO]T`
���P�:�����;�7(�p���X�fI�Ox੠��fs�CTpz�j8uE�]��(��)�9�P�rlzИ*�ܪ4
TИ�}�˨������*$A>�@eˮӡ��ڝ��_�?���ԥ#V,�ވCLZ�$'�#�r��u��1�DJ���T��m�e�8_8��;粞{�0&����{�m�Gӭ�ouVv�OR�����2YUN
�Q��0Y�Ip�B9���I�D�>�>�S_y��xܿ��$HqӚF��!��2��W,5m�G��,hWk��`�+K����f���)�p�y]����QZx;�����w)��)�}Bs�5 ��|�2��V���< �����"_έ�����ⷔ�ďE�=��>}5��%;͗�����K{����/��Z�����z'
���]jǠ���T������O��t_*;]Ӌs�+��Y����N
��!@u�%*p�{��	(?dh
+�G���i�I���'6�ey��,�/���/�����Pp4wƾ�8-�����
I��S����i_�KQD[Y���V�������'�L���;��dq�㵋M~yXiz�0v_���|���a�[);,�Q�9�7ȣx�Uf�ԛ.�3>�W-�U�w�<.܁�*�Q~�?���#+U��� bm}����h'4Ya��es�5*1�!"�ϗ�&&��x��������;�dg�%��!l����.6�����<k����!�^y=����u�Z��Ɨ�����[�]z�?����v^:Up����{��$�5���?�Yǲ�:6<Z�#M���!��o�_іbz��9����d��.�x��kZE:��9"�A�r>��[�2�E/D��Fe�}�st"�Ъ�x������f�/E������a
��)첀=���#�T���c��h��f���j���!A>��� �EP�`k� q�6|8%�wc�t��w���;��Т�Kj#��ճ�7�j��1-��8�jm
Ms����%Rx�����ݼm��{�����o[;���/R��	��+3�}�^����eR�]��tZ���Հ� W���~� ]�F�c������X�������SO�"��Se����C�^	7��W�Ao�_x����N��d��<����p����(!Z$"[��q_J6�/��[P�<q)|����[)���>�&+��C��~)�`���Oz��HC#/��	�s�;�Y�q��3�q���#��d�ߣ����u� ?�=��.��2T���"eq?��@��U8�S�q	�xT��`�ZƖK�YO�Q=G�a�^�[O����=J:�tZ&N��{}|)H$Be�0x��Y���5�$��+��P4�ks� ���2i��n�������@Ϣ����I�}����b�X�B�`>_>�4�3�[��\�q��j �GG���:�󟈔bL��$�~��]��7L�Z߻d��y�j��UR�J>��ּ���4������4b{*��EB�E����&rR���9����u��w��Υ�U
�u��^k*�*U�t��:��C�d�%w��ݫ-�N5��O)�����\��W���2�݌!9U
#}�nM�W�#~���j~�ųKѐ.�nr2j�h�A�F�0��&���w2���o����x������3
�]~(�0/:+1��l�?)L�I��'�h��渆����0�)��#�KT�uh��^�;d{b�Y��$�dg1/�ϰ]�[�xU��NV �|Jk=Uч�q}�a@����$cKh%�Mt�[��駁��<����T��CM�x#ޟH�U�n���A�G=a�9���+�l�<Z�ٹ��4D��{J�*N0`��'��мٴ)^�Ϣ)���;��%gl�We���Q+�
w&�w|i�'���A!)��XZ��A�E��k����� �RaN����J�4�9JV�Mú��)D������i;�|����g8֯�u���9�{L7[@(2[D�%�T�SbL%���=$�h�N�c�8��6��8����E��&mɯ�E+(�m�,;f},�{��:��LuȄI]���6<�9��B��E�C�{�6����á;�)�C��0����;[�5��a�ȯ�//�Z�)��5S��t��K����GB_C�YS9:��;�mcB�b�tڽz�*��@M����%�8� w����C�cQW*�3�^�.����ap:l��������K�`���ü��҇�o�SWF������8�f�l9Sqs��M���1Q�3(���G��UV��!�	�j0�������{`ܽ�"���#;�pnb����PV��\+T%�N��w�az�Q-Iwz?��m(s���<�O�j�D����}��y�N8TE��	���)˗�G��JJ�3-��	�[�:'G�t.�]��j�楤����}�N��݌��ej�cq�(n8�K����ۥݲ�w�֍��O�����N,�R�F�!6,u�C���f�V���w���v���i[���8����,d�3f�RM>u%��uDPo
��l�6
�|Ta�����:�7,wk7�Q'�T�jg�.�"[al�T�_���d/斘�����7��#��A�e�lu�!�+��Ot^<��C����GJ�����4\���*�hξ��|ŝ����WP���*z�L)�1KXeH!��~|������qu/M���c��ſ,�e���v�+����\ K�'94h����-�Op��dȈ��Y��ۣ? 4.�]��k������6���g-P�9�a�����4vtF��5Ĉ�H�/k�(��*�ΰ����׽��)�G]i}M$�a��Ҽ�"Ĭ
~{���K�ym����CJ�;/�ܨlÍ���x5߳6+C���7h�P�?�6��"�B2����YP��[!�9����'�#x��ͻx
>��(�[I��9Z��R�(��)w�?����-c}�#�~	�Ǘ`�ϵ��P�8P$5<w��>�{���'Z�P�e7of�xE+c�f�9��?���F ��>��>�<-Z�Q�Q���K?*
[_��u�!B�xɩ�Q�
��)�� ���1��O�f��ͺ�휗����gPg�H?;i?OqӁO�^_~�2�r7�O��Y�Ȑ� A�o��ȭ%�r���a����H\�?�;��U��][࿗�	{�����5D��`�u���������$$.���5��� �s��J����i�����噍���i��^�-.{M�LX�a�m�Gy�(��W6`��.N;��aQn.��-�D���{Y2o���D�\��j�a�)�k�w�fO����ػۢ�.v�,�ީ�Yi�������Vu��YFâ�?��5.��S���^��_5��F�g�6[!���u�ܬ�4��v:M�J�}5��4�T]x�~�#s���vl��awH83k ���[��J.�y������x�5+��4�AR�I�v�m���\��SNJ!��0���C�~-j"���F6��ID���5E|(�z�E?J�SN��p�B.34�������o�FwL�R��Z�i��g66Մ7⛺��hH\����=;Z�x��MI� m��<?���i&���gֈ��i[���� �Gk�,-l�V\!����ͪ���;��{0�+���1��t[��<T+��{.��>!�T���u�9� Eh>Ye�7ཀ�ڡ�8@5ir��
vjg4�����S'��S�J ?���$!J6�=z��~�PGe��?���5��ZV�;�k@�"��:=Kׁ��-�^�L���9��*�۽��z���������:����f��HB^�oтO�)m�m�!$J\�]�f�#Z�̨��2��t�Ԧ��Py�۴�ڈ�*���ԕ��J%(@lv8S�&��
j�`PS����Z����a��.�>�0�� L�w�VŻ���o����d�Qd��k �Y���<�K�a-H�΍^	m2�(`oNxQ�^Ӳ���N�"�^g\��IQ���$��/�]�8��4���B�Qn����o1����Pf�E�>�X#��)���n.�>>g>5��G�%j8�5+_�ӟ�L����u������i����6vX5,���鮶V�9$��N�Yi엽_MUm�5��A� �1��Sݣ�n|Ѭ����w�jA�+���#qx�9�C���!]�C������8�8ST�:���BSC�N��[:1Vj�#�`��w��<��k^�c����2�: %(^�l�C�U8�2��	x=v�T�7�g���KlV�K�juN=��g :[�"��nOa	s��7�?-u����Y��g*���ΰ1��I���L���1Qe(�c��w�%h�"e��ʦr|ù��*�A:1����lv�'|��2�	
���l~V�=?+�#�g��"b^sg'���M16�[����a؞�*�Tb�LD�-��(3lm5C	Y�ۛ�_�.���mQ��"���Ӣn�.�>
+��������\̴t'��D�=��G�-�?��������*�:t��+aX���N�N���H����ۮM"D����%�a����C��U��=Yݼ����'�[Y~�F�3}U�^��E�w$jҕն���U?J���i�<>�������1tY-���l` u�4q�7v]�ޏwHs�nV�\� y:
U#R��M��`�W|�wkMg;���K�rn���6ˤ�M����>P����ǧ���Uu`����v�w����|���\W��c�n(���F?�p�^AHB3<��wzV��ޟV��˦�&�\Q��`ҳ:��l�NT&�6��M#R�@��KI{+2��+�qvL��Т�ֶ�fa0MG� ����9U�W������A�'
eq?J�lVH����`�����SOy��pZ˅���cט�B�x�Chk��`pp�hqR '���ǎ��YH�q���v��r�L���T�C��֢���לӉ4%����/��	B[+'�K�dx�/��g���S-s��F��3���_�/>��15�d��t,�O]�h�wG��&	��	)/��E2��R(��Ru%��s�dgԿ�?|$[��g�278����8�z��Qi�_kܤq��,���#wz�	X�J-�p���!P�ӷ�3	q�PDY�_� ��+Na��.�K�m�)�?��u�=�0W��к���s����k@-������YZ٫n�Ӳ�rj�ۑty�B�ma�X�W�XA���}۹B�>�4���F�	u��*�x"|��)�G�wS��.P�]����ԕ�������ym;)>�3�[���$>R�31*џ|;׻���CYĳ��H�H��>#y%�C��=���mP^ �ҫ�K�.n������_5�z
�Z�F[��c��"�Q�_c��)?�F;Wn(���<�./�g�YfIDߒ'��7x=�SO
">^]j�)n�����e۸}�3�%ܙ$�����Hz�1�K���T<P�� ��B�T�d��L/5�d��e���a.���Ċy�o�T��S(���#��Ƅ�O���!�~��A��c�}�"D�z��@�Y ��l`2@�|��I�j�Ә��zͬ�H��
���4�u&2���/(��nW&�YZJ����q�1�m9�~��>����	��5��(%�R�ysRǲ9wvv�`��;��ц��5�,�HD�Lx�n�B	/���!x�þ7�۽�|c0��UxJ3�.i�O5e���:XܾM�fa�<S�ƴ�2�l�������7!��/���%����o���g���p|d�S�u��c�%�gb�Qp/u�~�\��y�M�g�o"�F)��.ۨ��8�3zp�MoV�JRĳ�eѹ�A�*3����`�� 3�~Ŗ����C|����t�Nv�i�tV+ix)ᵵ�2CV��e��օ�né���u]G~��o��u�Yǒ3�fF�8������=���:���������4���_D�K�	�Tl:r��ĺ}RԻ�oC��h����3������p�%�,�L0����E�D�0���-�HX��pN I`6���*�{�y���w����3QUƔ��S�p�`+�O��m��Y�'��p)^|�G��p_**��d0r���P��N�2��ɡ�S``�ela�G�n���#���R��`����@z��;ӛO=7�1��~����r���>!��&����W�f5'İ
	�q��VE_T�{� ��4���S�A�����;ęp��c"������K��Fe�=�+�� �$����^�v�W�`�>������潊���%K�02�Tu�|�p�Qu�|*�c�3�& F���Ža��m`��`��L�I�qS���`m�iy�*�g�оU��| SP�.*��%�ӳ{9{��1�;��s�j��{�V&�Z+���?k�������A���m��	s)	H
��"j�*QIȿ��;��#�[�Y�4��{�ѧ�W$R@x+We��i4$sn��viD&��v��E~�/�y�$2�~~����|�R�A�_���� |�*���eg�՚��n�,��| ��6*m%�MR���
��$�%q����d�Q(_��⠗�׉Z��۩$&���z+x��N�}���+5rU���u�w�_~�����/Th�*n�9���'�Y���i$w�>�����΃�o�J=����E@��4�wi�?�7�)Z�M�eq�� ��	�!���x`�ax�j�EG��u .�oڒ�˪\�yv�F���N� 	�[`~����E�Қ���1��Y@v�d1�����%�/i�k��?�{�T��kK�mv3֙���F�����7J� s��l���;HGj�7�K��������tʈ�sO�D;�窙8Q�����?�e��D�
�͐7�k:Z�0���|��-G��������@f�~3zA)�O�4a�;Ƕ��!�\�UW.��ej�����9�YǊs|�9��;'U�M������1X	�M/L�]߰�[���o��>������4�)��3��~�O��������HB�5M���,`���bF��H��5����;���IW����=��;:#�>��Q��I��<g��[oP��a�֤4c$�q/��ZS�%-Oe�Z�ƿ�8}��g�t}E�a9,@����M���?�H�Getǎ�{�q��@�ُ{��f����m�wM�6����'� uȚ��"Р����i���w3�7%R͒�[��+��O:7��q�'>#��=��:�d_,4y��J�
�6_�R�I²��T�l��pAʗd�S��.+�}=�)6��7�Y�0h����>��1�&<n�B��qw�iK
<z�&`�v�񔳧�#1lȳ�0yZ\�l�;sI)��.�2BS狽X$r��u��B��a|C����/�����y�[�**ym�����E3�L����h�i�|{�|0��F)Ü��r�P� O��;[�M�흲�i.���*N�qA�L��MHN���|���0n�p��k2+�=��RR�p��v���&s�
FyIq�$�i�Oj�PJ>��Ny�����_�v�2��ۚ��3�>��o 	!�;���*mֽU���
Q�Va���E\[sF�˨�����ub%g�.�����i)<�g2;k��A�������R'����*�m�l	���'PR�jND;<�&�f���󴻧���ʷ��)���Y���񌏹z���٠����#K�mȝvg%�j3MAr�+TW]�CE�B\:�N�}ՀLq��پ#O�{d��k�܏
Pvm�\�f���nn�]ôB�.��g�YƤ"�����K^22�KR���e�8��a�_�w�`N]*�x��j�����D���w7�{`��ʼ�yO��������!���z2����F� ��}�E�Zː���t���Ӱ=�i�n.��2`Y]
r,�6��I����ˠ�d�ѪtuH�.�å����X����;r��d�T�7�wV�{�ӑӻw3����7L��O[�a�'�^��\�s���k��Z>y���mɊ��P�8�+ܷP��� ��6��l���`30`d�5��ߓ�� �#������� ќ�1p��D�_���Nj�\|:��Yz��k_�~���1)���6�������'ꤑU�)�3(�aD��q�g�:X�`�_��u,�-l�� ��iM-�<g:�|�WRp���Eˈ)3�v�`��\l�I'9EM��yM��[^Q;�ha��F<h�G.$U�G���.���8_�ž+��Snj��]=�V����>G|=G��N�k�_��nuT�;k�_j]z��dy�V)^u*Tu�۰�����,_7�a��N#��<عf<�r��� ?�=�Я��_�V�bV�:�u�ir����ä���E�u��� ��Z��?��@ΨP3��0h'@xd�d����l�U������������{ ��ߓ;�s;%�꼢5
}MN�?��=����P[ּ�`tG��/!����}%w��$�N����DO�2ËgD�3z@_[�4���y���jw�Lu�x�ܠ��0�[�8G�$�i�|���=r��爰f��h���vs�hD���.�xWo�Z��#��A���j��{��t�W���U�
�W}!krc6Z��3�ji7���&�V'Fķ[:
8;t���(���x*�:p�J:��V%Y���Q�y�yJ�"���R[f)��U����ј\g1v9r�k��TNQC�hH �v@t�l\�� F6��������I��;n%�n|tT���8�aZc|׎G��Vw�9���c�:Sb�u�KPA�<���d_�f�%�*�a5�����j��k<��������b4���_�΂l��أ�$­�u���3W��5G켊��ރ7�u�/��Q5!1 K˶kj��q�s�G�_���]�����3�e�Pg�A�'T��0��W�
R�W@x_��d�W�*J.T�P��{f`4�2e&����'Y� "��������՟�����t�s�C��������0�Hi_��(��{(A��2�V^Mȿ{��Z��!��޷����A�����g6]�CAJp;5�w��������<Eԃi�b��z� �Jr.jec٥��q�KDbקB����n:"��_������LZ'���v�w����z)�bd{�)�5���N�jg���_p�n��A���x�r<��RE�x��$���z��=��yQMk�����w���@NCi㎮��[:�Os��
�������2�`꫄QF�	=����IC�����s'���j�� |2�ɺ؛�$"D%�E}�ll.����¼0�w�<���6XO��(�-rDQ�=h�s�-v�W_�c�T9�jQT�5�l����O�2�B!v}���Xk��Զ��c�q���_9�+%Y�\t�9P�˪�m�lTI��&�qGL���j���6��¦tDP����ڽ�?��<L:�I�Է�j��oBu���@ ע���?��`�7���k�91@�3Q�Q��y���7�ئ�����+��#�D��4��ƺS�x�A/�@��+c�3���K�F�&��-���O|�(�Ձ�Ҡ��V��"�o1�T$o�jM���E����7�T��Q�c��#���w +T�?`�[���y�C�Z�����Sz��^R҉��?l��	�/I1A?7��Qt��i5��U����%`��㻌��V���q�΄/¦�}}V����{��;�C��J$�������(�e��"e����q�V��d����D��J!�HO�N�'Ա,�̺,ٵ�f14op����*�!�pcF���ŃkyO��UQy��ͮ�F��.��BK��Dl<���>j�cd9+gW5m�"��fl�wK��=��m����Y�ʶ"�
L��\S��I_��rh-�/�b�Fm�S��/.��Wld�{˹�i�~�	��V���=ۺ�X?�Æ����:�L�!3�wj�����*�BK�֬�hRs����e(i���W]Ew@\��������v�|��nZqS�985����1���[�K\(Qĩ�����)�֗�W�X��=��7��m�ˏ�Nq��t�i��k��0eƺ3�&��5��Z���Mf	e#(^�3�H�Z'yk������3��|��bDo�EE��6Ç>=������&��*h ��/�V�`1>ۀرk+�נh4jT�> v�)�b����[�[s���Y!����ogk���ߖ��`�}�z�-~y߫�Ϡ�U��)~��֗4�}��_lYZ�vo��k_3��	^��Ăٳ�N�w�r�t�o"}�-o�d}Ŧ$0�9�0�IMx�9a���䙡�Z��!P� y�+d��4rS$��it�h�Z��7 �,w�Bh��º��w�-�'ڕ��1��:�@�������"���[�5�����9��Z���8��8~ߘ`E�"WV�Sy�����_9�c`W���'����7�S� {�*2��N3�\���֬�SNR܅�������Py���G³<����|e���3!�]��C�
�u�@}_~V��ʯ����KVV|�{sGɈ�?ø7��K���0r��n�Uc��!�1q9GU��35�ӡ��%��#/��>�:}��ْ�.�%7��F:B�ʻi �Mn0Fy#�����ɳ:�sM{�0���������c1��]���GBb�ƨ�[�ϻm1䱔[1�����	<�8�~���on+�E�MU3.����zڮ�8n�3�N5�>n�1�N�Ɓ2#H	����������Cp����i�붥�V�]T���m\*�/����;K��k�u�LV�o��ԜMU'�D�݇5����L�iM��xp� o{Y2jqK�D��X�p���&��(�����?���"�X�,K� QvB��B̖�Y���3j˅+�B�'�TP�+�B�Z�O�C"�L�H�>�` :�U���{�TX��o�H�3_}	�|�nE1���Y�JU���_�`~��w��2{
c7V�`v<��ּ�J����l�(9]�o:1�0��\q��v�_Y�������d޻��J=����s��QW�d�j�k��6�V�e�s�F"��z��/'�ɝ����ŕ�&ↂ.�0֏}���ܴz�r���3�8^�����=�����H�=B�/��@n�9ޘ>�!�e�ޏBG��S'x`Uj�=,��AZ��%E�W:.߫4�et�V���3���)��xW�J%�r��M�P��Z YV��Y-��y�S��	�&.��p�?M�Q��P|i�B�T�/tf�k��>�[.7XG�1y�9�����}���i=��#+u���Z:ߕm/�xZ�D=X��4�v6��i�NU�e���` �b��G��T��ӊ��{W�XQ|^�p:���O�ҹ�-�e�~sҪ�鯸����銱)�Wc.�����X�G$��(�ιCqs��I�<Įj^jd���b�x���wC+�'A������(`����um�o��h�iSՑ�cO�PYt��SdM��>�*:��E��O�f1�s��1�7�^���l�dU���,�\.��G��d3p�f�jڌ�x*[`uJ�S�v��]PM]����L?a������F毠�e�JGU��X����Y����z�mB��zKsӐ�ܸ���JN��!���Q	��'4�[w3��[���e��޽��'�[�_Yj���Xf��7�F���R�(p�q��I���z�����
�v7�i]_7Ae��4�!|f	L�����1Q�}��Y�I�#?O� ���q��׫G��)���i87�0��$W�_;#��R�
z��]�\� �}���ZP�4�������nf��XV�w��)����F>kX��s=�,�9�(�o:{�ӗx����}����"���e�ڇ���C�Όu�S�^r���+O� �~�c��0b1�v@���*�I��7�.6�)c,�S��gR���E��/$D҄ޕi��ێ����3L�߼�wz���E���&jT�f��z���k���KH-6J����W#�S��)(o�$[̚7X
oL|,�s5�Y\O��ܳ�
M�\���b�ύ�a߃�#E=��!���=�)2[����^/9���S���\�c��UF��4�B�'������@u������t&g]rH�I?첤/dG�THm��c'�fԧ�FA���Yd'��-�8��J�2�h�$��h� �#c�Ym#�"B���K=���Ry�"��s�+��p��/�p���b鍄�k�,.��׬����q�g �w)�ї��!Tp�9�t�T���%���^[3'�Wg[�?pAˤ�-���V:Y�b�_�9�lZ��3-�u�M�l"�a��ֽ"��LG�+���͌��?��C��#*��Q��'���w(�P�vܑ���%�U�Z���]M�{�e��[���8�9�7n�����yrW��;���A~���oB�0`A�I��a#��3e�;8Ů�|�t�m�}�	P��>��4����
��J���]�V�R��حѬ+8� n�2�lv��%��oY��y_uY�b�'�;*�"k{E���A�G���������m?/9~�`��J}1�͎$Yv�r(̞�Ң�����f�Y������߉�<C7�@�Q�Xi��,�y9�n��S��p۰���,��f��t*CFS�xK{P�l�#f�>1�2|�鬂�|�A%�)ǂM�S��b�� ��ڂ�
�|�ģ�!���茄�3F�����Ґ#+?���F�u�1Rd�Z;�������;i�Sc�S�.�7�M�r�����g)������O�M�l�oƂB�[�'G�2L;�U0k��5��`��L-m��#X/�2����n�q�����s � �Yh��0�֧8��M���%��`@[+ڽ���j)�K)�g"�2�TܛQ'�Q�8�vz�SR�QdMM���Hu��;۪.K3�����{J%���	��9/���.��ԅ�P�����0�J̲�Kؕ)Dx���萑�Ƙ8�E�'�.��{�H�(����k�x�x�g�����;�s��
ͥ�]��t�f[#�:�]"����6"3��b?"�λ��� 2�)��m��+�F~>K�F�3v0o2�]R�����L�B�ЉɁ�����&
����ܭ���i
����]5\�R���9�0�����KfH��Ս@����u�vP�!	NPU����-�\Z��G� ��:�J���q��
�){r�Q����{p��&�N|�%������m���������;CP		5�gM�U|�O)���<2���4�V<ߟ��W��+�F�t��ޛ�+W�1�!��irNܢ<2�_��+����4�����Q�z�6��d�#��(�S��`2[<D���/��>��|5"9'�M�3������,���f�כuG����:�W�z���Cj�����kb�ɰ����w��۹z��{��ٌ�k�՘�D2�^��"���\[����eL�>���rl�	F�f<kD�m�I������ߞ�oZV�'�f�y��s@�T�mW���@ J�_d��q��i&����sh<�f �u�t�cK�S��i������|z	�� �;簃as�����\R�ztì��Y�t[$G0��.y���YUd+If߉��U�^Jѹ�-�����0���l^�JX�@\�Ǝ�烴��ͳB���a��F���Y��4@��].߼�e2�rdja���Q�3���kr�O?ra�W�9!�V��������\0К�ш�p��d�HGP���JRO|fi��\��4d���b�&2��:�F�	>����U�l�lf�Ȧ߮:�Ca'&7L3]��2�\��E��YQ���NW� zr]4����5 K
Rp�N�/��@�v/��q̸�.�����Z�Gc�<W���?��eJ_�/��ܰ^�ǰM����{:x[�����~�N��X�\	
��ݔ�:�!j�ƕ�^Z9|��1l �� &G�*�6Dt�$��p��@Y��-*0�犲�HSg�&���7~������	��/���!��s��PuHu��ϙ�й��B�+���|�!Í��C��T۲l�z~���f Mcz�<} �ݿ�+��>�#�+��q&,�)������R�R�4�9�ݽ�jV"�{'̆����m7�'����){�O�.7�;�-�J�܆��y/�+���L�aE1f%O�[7�d������!9e�O����/�E���W��F�ީFT�`O]��^�S�]�TA�*+��N#hD��]��"�!�e�9�.�l�Fy��n,_��!������əOi�W���M�u[Q\���K��n]ۚͰ�s��S�gEev�#������졚���Y��BW>L���o���9\У�-�>A�Z9�=h�ͪa%�����Lg����F앥�0ٳ�^���9]�5�~�TV�x�4`�!>�se5�0�|-�nσ�����2-gX��%H�dܖ�TەZl�tY�-��D��v���қz œ��`�/
 ��J+(�I��Gx2)5�4�8~��n�!�����5�"����<���}cFWܧ:�1:N~����=cqfo����0� ��z�S1+q�Y�H�ל�{\�i5'��;Af���������I��&�n�V$SRh���)�tV�qtr3�j]�tuN�*vyy�Zf��� ��.;X�Q~��E��5~������yp�J��J������c���2�z&�E$�7G0��[j �g�#��N�vҾ�ϊg�t%V��oZI]I�UK�Y4oL���N���I8\<~1����?�"3%�˦l�)f��?���D����ȄO�/z���KD	�6� kf��8o/�`�0~�$m���V�׷�Hm��Ծ�Z�����׏:�,�/k��������y�v��%.���	j���c��XhE��o��I���+�����M�?,۲g֙�w�e�Y`S[J����?�N��|):Y>�����|S��m"�!��7g�V��m U件�����?���LGP&��STۙ�ڵq�\F�k�>��?��"Zt��ѶE,\�~�*�u�h��'k�!�p6��sݒtX��޴��(9�8M�WB<�5���d��s�Mkr���Sm�/�f���nv��8��Cp6��,�N�����Kk�Bs�W�F�L��"il���1C@b��ŵ��8
� g�����i��� �ٍU��)����bb�H���Xuxn��H��>�w٣lo9r�� Qz��sl��PX$�`�MMӊqu��Z�3)5�К����= �I�H����-F%@+��7�pp����O�n�}�h"���{�<B$���<x�z=�u�1�/��呩���thu�W�8A0;��~�>�e�х^��j�����X�y|7c��e��@�K��F飯������J$��x�}�[o�������E,�AQQ�nP)��&!#�:d�ҝ#6%��5Bb�6r�����}���8��s��y��޻��L�po��#�M��"��#_BR��_u�kϫ�Ϸ7J�(ǽu4�^�y_�.�2|Oe�ǵ��/��E�W�`͇hlW�Ȉ�M��~XJ����1Wb*��qR�}�\��@\���\����Z퍆��nj�ԉڥ+U��Nu�c���Ch����!极�8�bƘ�����8 ��fζɃ�����ʋ���Ƀ�G�ubU+�G�8r�H���QS�����h�{k�k�O�?�?ZX��H%�����|Z��H�k�	�d)dF���SI��2$����!	� +�ke�����V�7|���	>ȍ}BL���%��o�{�6q:C���A����5��<H��c��rȜ`v����琯�̠��9�~y)���?��q4h�ˆ�I�/ӽ�J��z�Ǭ��7�4^6`Yf�n����(�[s��<�k��Ik��!쐶ͣ*u|�N�ڝ)2�r�"�N�����;W��tl?�;�6۩�SⅬK�vNC���=Q0�J�q�K-6�q�`:��W�����~�@��sJ$n��话�9`��4�C`c�J�QC�6գdo8�%���D᯻����[�3�J���Ux���G/�̚�8��In!J�D��s�y:E�?��>�I�_����v��tx�z�S���lu�Y��S@�4��Z�%�B����:�����mt�ʧ"l�X�����N��,39�S��L��� �%���=�@�+W�)&��rD�ڸ�9}ϦR������?R�H��u� �i>x;�)�'MB�zB�E�..�.���;ƚK���[�SG?ɼe�46թ��� y�G�ߖ�˳N�ћ���<�~ƉC\4k�1�Q%���! ���^��$����ɆL0�
*M"#�8����gG�-�:d�j�����������Ⱥ�����M_7���냷:R����5w>7J��%3	[�.fL�?Ѳ�I?�YJӈ�
ήb���S��[�5l���2�}<f0� �ͯ����B�Yr���p�]�S�74�٫BB�E�Yū�M]=a8#`�ekv�|�&�'d��9�P�1�BN�n����@�V�ѩΓ����V�i$Ef���;7�w�_��W������ T	b
�1�ݚ�|��	�J��eUi��Bi����B��N�|�(���->���ŕ_�+��c�w��fE�+�S,�'xLڮ\�����r�/S��n�|t��im'���;d��R?K9��N��W�-	ׁS�6�P�n�y/�ʗ��Zc�Y�=1 �Dt�Ovs"U�̃����6�궗��	�,�\&�r�o퇯 �uF�9��H��pM��)8�j3�ԇ��]��z�Ss;��X4J�HM�sQ�S�bcC� FՉ��-�R��ᨄ%��!�T�S�?�>�Qmb���F�5+�Ӟ�T��<
�c��B��\�jH�|4�k���o��館?;�ψ��0["7O�y"7��/�@3�7Ȧ�rb8U/�.�{y�z϶lENI�R��g��~Q���v(B���Y�m��m���,�D
r\∯����'�z.����;}�5�lQ��L�����s����!j����\�9�t�\	3�ie����������j����5�5Ե��F���Yc���d��*�t;Ƣ�Y]�?���*n:�����p����%�)��'!F���U��p�/3%F�o������.��c�N`gZX�nR�lfvnU$pYD0/�V\??�;���S��p+ؾpaJ�j9@�>jes���6�A�d��Юu�iHG����OD�T#��[bCg4F�&͘�U�G�2�5�L��-�"��*��m���Ut�틫�����Ix�se�SD�*�N1�8�i�:��R�]�Q�3� 1\Nb�bc+{�WX1�"g_�~&]?<ܚΔT��B!FS��*.�y<t�.�~ޟФSj���Cs���p�祝�QApNJf1 ��Xm!%#Ο&R������8M��kdDF�qT|��f���ŋ�����\�@@������h��*Y�9�G�8ŷ&�y� �+'n����L�J/�X~y{5�Q����"wD�u���tJ��I�pg� pD*�!�G�{d��d��Lв���"rI�����wg�K-� ��o���f$� 9NDo4�p���%������H�G���_�/"Rv�-HY��v�÷P�aX�Uv$��&�@�>��79�_5��B#3����Ő�/}�FQ���"�e��><�T�e�v�|�r��L�J�C��(ֿ���(��~�����,j���Ҫd? 7�w�0�:l�R��WrO�̢jw2�;�U��\���G2�z�&C_Ԗ;�d�d�q�a���w�a{P*�~�t��:=�	~ �o���zTN��~��w9�@v���Y&Tυ�ߚ����Z����~"Z)��\�	B�6����r{T���O�Җ~)9p"��@@z�$��U��@oURH���~��N������^?��y�F��Χ�'��=���*{���/k@�s�h�{3u�E.R\�����}Y��n����0A2"�p�f�w��R��[Y�*��r�s*�^Q������hO�K��J!x�r�@pc?S!f�^-�4dD�+�GDD���K��(~�:p�W_�#H�s�0ǡs�i�g�؁��o[��+�u��C�h��:���\&�[����kY�ҿ�18*����[bp+�+����vq�|�:���8b�)����M	�DQ���A˒�s��J�j���˄�w�����;#�Uդ�ճ�G�}�aY��C��H8��9���и�_M9~is5p��@OAE(�+����rMZ�CZ�����g��?ǯ�|���rCM��^WPA`���7�`�!��{.��,I����L�L�L^J~�L\_Q�MnMʙ�������ĺ��Wz�򉇔�#ǝ��,c���o�Cv�s_������k{�MK��P�>�����h�h�	G�:�+9�~5l�#_���}�~H+n��7i`V�mm�ep#گ�L�(	H��J���ɟ[pt-u���� �!qY�z���lU��]܋w6u}��e�>>��������l�$��ex���?�o)WO�S�<��HF��t�۱�$�旡��m�R��׍F�Z���~�x�7�?�@&%��r4���V��iur\���PF��u�x�P�����{�F'������JI�3�G`:�w�f3=�@�E��%M�j��UՌ��������9� 3����haTNڏF��9�<�RS�3������%^w���/���Ì��x���X}��ʬBS�*,�(,����̔�$�
�7���ϴ�n�V3��|�G�\)ܓ%l�h���O��D�9�?���Q��8J���-@<���7`�7�b`��`ݰ���F?4-Tn�g����(}4����� ����7�ʂ9�{\��<������	y���m\�ۥ1�F\��W������z�2+\MPe�����--�f�U�X����J�W��,���U���w~.B����~_���V�;o̾��d����xC��3/����r���4�h�k-O5��&��5���h�I7��J���n�����!��mkv["���^��|j�"�GC �w��Y�u���I����T��C9��l;�k��{K�<�[>���|��R3~�Z��=�j)�c���_���G����2Q������?���MF&���'iH�m҇k��݄�c.϶���-��/�k�-���v�\y&�y�� ��~�1ۚ��
ƟB����>��� �!o#DH�-=��>|�V��#��8��i���G��o8�O)��J�v��{��R�[�%�y�:/gWX� {.��p,���Y��z�4u�ca"���]C�Vwed���Le�#U�Y�G.u1o��|���1���ˠD�� J�*�?�eM�_��	�o�U=��,A�:�c�O���l)�����<E��HW����\�O`.,r�Y����ϵ �C'35a%��/��I$���/����꟮����n	���u�Nc�,���"ot|#6��&�7�W��W�s�âT����DH�}$vM^&X���P���)h��IO�o�l���4�ܰ�&BP\��uw�u(؁��LknBZ���Hqd����Jx#|�8�;�KIB�HX�wܜh�{!�,�	���ԣ�v�x����U&�(���t<H.C|^�	�������^S��tޟ������F-b�'��m��N����Ph$�K'�̿0��1�/HS3]�t$U�/�]��|
��7�e��ل�®�T��,��U�ڳ0�G�N�92��'�M�' 0��Lk�T�4�]��j���&�߼�W���B��o�k���.��!��Z�#���Р���/�Hp��m�����'/�}E~����t�ooBʈ����3�&���X�Uv~�8�h��T�t��e%���؀�����A��	�٪]�y95��g&W��U�j���0��@��şjTe��cìG���o�7)Q-�ؗL2?��}�=�PxF�&2ٲ�q
u9��m2�^��+2����k�ը�����^�P�������^�otޱ�� ��|:�]�4f�$ nrg�3F�)�*
�b^Ec��s�Yf+�
�Lε�����T�8w���+�P=���	����K6`U��׉Y�-��7k��=�����~nq�z1�K�����4�N�c��o�3�JC2_��ϔ����"FF�ƶ-E%����ְ:�����Δ��= c�1۲�8vJ⛥ii0>v���&�7��7����;�e���O��v�a�r+�B��\��Si�������R�������:YB9 @F�B� ���%y3���C��Nx<�x�Op�~ �9��{o2��R�kf�V��B�۵� ��,�8E`v4r���f����qX��)���Q�%Wa�����ŚF�pRR�X4@�t�ԅ�7�Dn9-�E8�n*g���v���Vw-������V�̢�̋;��4��"x���aY�6��L>���t���[En>�oPv{v��Qnv̠�q���,�\vC��^d��ZtJ&ǝ�w��]xgC���ٷ��?6*�vs����j��6���q������:�5��F��D�Y�0��ʭ�`B7횄���-�G���d����]����p���,a��8�����/4�!��2��Z�����!w�$�O�����M�)�4]��{� ����ɔʉM������'z\@�t��M��=�],���h��Gr�s%ݜLvu<"Z�(^c�3[��i^f��px���U惀�O��+`8ʗul,�y7�6� "�C�r����cN#�b(ZJ���$����[�l���;7��v!��/��y�n��ն�K.1_���Qʃy�Rw�����R�J�\�����O:��iI��[(@Ë���0��ĂNk=M��Ѵ�Y<���Ľ��9m��b>��L�{���U�!��)����$�������T�J(�u`y��Xm�(���v�6f}N���4?@�Z�=j��B?��ضB�����A��X��v��+���}?��H�"�P�#sI�/rS���F9Ъ�}#��LhM�hs�)>���f^~�(�T#[��#�}C�=��~&|_�:>Zjkp����H�/|l�}�U:K�bd��9Qu?�0��5r�;�P�H��"�USR���}���
���<�LE!�79�#��15��`\dq3�����"T�%��4�����I���<���J�Y�^}��#����0�%Y���Pf��@�2��GtA&f��M69-�}���}h��P�+e5���6�e�Y�#�lj�J�RS�e�d(�Vd��ϢH�d�8[6zp��w4&���1�_��?n��_?�4�9"ZA���B�������p��F��-��UR��(�̦�0��ڪ��y�F9�+w���= ���yy��I:�֬4��dqR���!gwu����6ã� x����l��2x}8��ܷJ��m��[����"W5��F<r�#��0i��FN�l��+G��7V�m��va�)¯�T�N;�fz�-�_�VK���ʵ��V�r+�F1�GC �b�	�4���D���Pt.aC���b�Ǡ� 9d��È�n�_��Z�������6�=*9;��	��o�2Ί ��i�9Id]S�6��\T?���ea��Zh�e�m��9�W-��t�L���o4����B]f�B���eQ�[�M2"�'�R�Rqgל���%�����j%򵴎�6Wov� Nx��q�"�f�:�v�ʭ:�u�Xi�K����a�C5�):��T��O������]-)F�"9I�'���2�b�;ƄL����ߡ�^��I��V;��5�BEf��%;.����TNT�n{Q;V ������@�e�#M����N��(;b���eU��7�49wr��#XAs����nٓ󺎗���R����pKAR�Y�i��[�K�K�! �����Čs	A��������p��r�\pS�~�����j�����N��X��ȪN�����ڳ)�_�
A�c� VE��fY=��iE�O�59�C^�0?��'�S�r�6o�d�?�G:�H�)5i�W�����[^&�89����x]�/[0�<�S̒�߸-+OU��\^wh����Z�{�}8y�����y�K�]���m��:�J�URB"Ap�^]l7�3ߗ/��l��P���3'\�������7��\۬�v�~���2��g��`c9̷�]i�J�>k�&�Se���+�*=��KN�8��hZ3.�6��&�n�]��b��J���z�c��/��N����?F��C�ٺ���1�|y�_ܜ�|64}
����r���>(�E���	+��o�V�v�Dqo���28����?��{�у�\�׹TM�Γ��}z��>V�i�aX~�$��w����Ss�^��L�߭u����!-���߆iDvj�W�M�W�ǁ2�S����Ž_�I���
®�5�O~z��_9X� �O�n4�կ� X�\� �EnoU��K���3���m ɴ���xǁ��=��:�ʶ�2 '���S��!y��,��N�a�maU�1JO5�f�Pؙ�p�\�-�ֆ��mH���kͱ�>C����yռz��V�z{�sd�{��49�iL��? �Ku �i�|��9���r����|���@$W4)<�ݴ;f6�:�����|��e�=;�ȥ���[��E#.��lo�{H��WO!�[eJ���-�e:2"ͬu<5��Ǜ���Y�\��>i?~?���po�n���Ї��C>�%�_���h��{�󝍮�Kb���/� JAs����G@��0!�k���Jnf۸����{o���ع!l��V�{���}4���H����*N����΀L)0���c�7/�<��2��(eR���UWb��O�h��{3�a��[+�l����6�N�5cShX�d2؎���ZQM58���]�}�D~���%����S��ɛ­�pe;�W��9��6�������_ɒ�0I�K���V�h\T:j �E6o�i 9=I|�.0h.ۺ�^c��`tf#�bBI�x=��������a�P�y��lM�s<����E���{&r\��=��*��9�N����N�y�o��ZVd[3�[[m�:��p����N/(�c�Z��p	�d�|U��:�:"�I~�J��Ǩ��3����/=F��JV^�>M�����IPq^���6�5C0q����&t����T�_�����5�1�O`���kwz_�2Ɖ�_�F��Jn���L�����M�L�s��݊�#XcAo��h�j��/0�(A|�_�j^�:{Lʚd�z�r�,�(}��bo~���ね�Ge�o��r�{4����k-�jqs4���T8j�g�;�=im[��t��}��d���v�p����zu����8ҰMҢ���Hz�߷�%眳��Q���/�<n/��Ҁ9	�M_��}˯>C����M��t���W��<�^���Pu&(��7��p#;�{�唦^R~/g-�l��^� ȯ�N��927g=���F�N�ӳ��R���[@o��ª���K��B��:*;��u��<2��1VG�(��Ŭ_�5,C��T���~6Ee2�����p8����ٺT��^.������K;`$j9!h�ѐ%������\@���P�,"��VW���۸�B�th�}��H' �K�;����N��:o�'��?w<X}�t_�a��]����u_�P����*bL�E��2�Z\�N?Z�8����/Ff+����
$�O�"����Z�IE��zi�P�z�z�6��O0��'��/H�k[<�x��Ŗ)�1	G`���^��qd&0��72I(���X���h 0�6	'�|����F�oB8~VDJ[�#�p��6z�3�h���O��O J1��'h�*��@f�x�u;��@�I�|[�C\?�/Cձ"Ԥ�Hͫ/7����k��"FK�n��W�J�C=
�3gTTj,fNM*������8Ko����gW^<g�Nݹaxj�"-�j���
O�x�5^��|o
'h�G��^4ى��L%t�_���%"��hSȑ�ϔ��������T`���.U���0�"I~�Hܵd�z����1l&��j���W�[��{��-I5.b�l.����j�֯>V~"���3�8�ȏ�✥}լ.�3aP-ˈS�|��y���T�Lo2���t��@ܼp�a��2+�1�L���З������0}>��(�M�3ɩJ�����A��78~�A._0*�t9�#*`�S����N�/V���#��d-W`7,^��2���}�c~>C���T�}{���>7`���� ����=�s��BI*QNa��l3/��jN���@Ff7�ٷ銭�w���_F3��D!IE�E�.��>a�g��) �e�2���[���R�wӽ��>�fY���<g��z���߼V�Ni!*l�6�t,AƪeͲSc�C��~��f���պ�����6*<�6�'ɨZ�r���Ő�]@�Y֎	g�Q숰{ �V*,V�3x���`#Z���wyN��m��>P�[@#��Zŭ�[��R�f�+L�;�Ti�:2|��� M��/�|�!U�g�M��_�-�\����I������i�?1u�ʢ>͍l �r⨾־��%�S�^[���_4G����Zz�y�;��ka���3}����Ȭbh$hQ�Yq��L��ei B�sK9������E�=�V{��o>-�
� ���F�l_v�o���ž�m�A�c�k�\�%�.c.�m�X"�� �>��A%��H�	�;sb7�^`y�I�jyZg��2���(xΝ����Y�p\H@9��=٧L�xϗٞ�3�_V̩��ه���%���|z\1Y��s�<��x��g��_��}�}���t� ������ߔl�671��P�� �����v��xO���D�5��r�;Ǆ~!rc�8߻=!��U���H8��̝����ͱ�Ά���te�7�F,�,������}���o�V�]��s�-��;pc�n)ŬH��*�����xX@�wn߸��*��=`���%��C)b���32�x��}�����y�{���<\�2-Y@�R�`����i�V��5ĉ��=��ޓ�Ϥ�SF��l{\��G����o0�*�����Vƚ��&f�R��t��P��1��D��������;�(�+�+n�)aYf$����wn�l�tރz*��(��	����_]a�a��H�9��-{l�Ȕ�'�:�>T~� a٪H�.������&w���12%x���m�����ÔA�,ȨZ���&b��_Dr�=���MD�� ޫ�+ºp�����0�m��ul*��ꚹhhPP�Il��EN>���a�Vg>��쪌�?��������I��5�A}��f�Pv��m�i�uwܡB_��I�C9�5`�*ﯡ)�m���ŀ��Ï�������x�N���KL������%\z��qF#���N=S�6��z����s��r��d,�H,m8s���I|z���$��|���޹]��q�+A�����5�i�:x:2"F����P�l5�I�ǵ@^���З\0ۜ�p�,}J٩�qM�K�
P`ԃ߲4%]�Ox���繉��%N����ҏtm��<��+��[ps{�ȷ,� I�Gx��3(%�%`��
=�c��4# �!�e�������6_c!�=�y�Se�$r�k�'oO"���
�+Q&D�^Q����xM�7�Ĵc����ODc�a���D�������b�H���;�8�!���@�H�6�]?do��g� ʌ_���pih�$`����:!=���A~�o�	)��QET�7�v���<��E��U ��V��_���{؍M��5-̅c�ܑ:�� qώɠ87`棙�WD؅�Ua�U���R8F%��w՛��q%\����++j��]��
l�R��N��ӗ<�W���]TsK� ���?ʎ��=�X�l�&U�]/�MjH�'�
�"&F9@�p�����8°)�h�P��J~Q�L^�7����6o�/�r\-a��(0D���� l���۞���ݕ�wk�H6�!��3�=����D�V���c��p���ᕈ��G�L�����ŃrmJ:�>��/��N��X{9W�.4]O���2S��t��6<��t��qNF͞[Q#��-���ޕsD��D��U�Z�d4W��_s�W]�N�|��)� |�8���u[Y=
���S(&���Ig\��F9�:��G�SՂ�Q�(�K���5=��k����z_�E_�����&�#��C��XT1[��/c�*n�������7J{I��n�ulP�,��F,��OJ��݆;��[��x/y���E�J�_)�{���+ �al�=ʱ�O��(i�_�����S�bi�q�Y��[������g�We�Wn�������`��.
����`�P�M�h�o�,�'��w�Wl��NS�� �]�|dp?]�����H���;�k�$���i��D9�yĚ������/����c��5Ҧ���F�C$�k�zѧ��#�5Sݪa;-��TK�WW�BmNt��e`�?����}����#e��5�p/Xsh���O��V�[���s���Pcp�7��8��A���J��R�9�#���0�ۣ��s=��b�,��UTZ����@6|"_ ��'6$�mv�8��e�i�w5K��*B�f;�]��Y���@��[{�d�	B�V�%ڠ�U����m���^o-TNl���	@����p�V!̘W��5�i��d�?��A���}F)?2�bJ�:��[�2!\X�Nr��劉�n�`VO�*��/�U=Q,�C�J-č4����0|�OH�v{M��jh򆇎3�]�����ӻŇ��x0�pW!q�u|[w�a=X���+vS[9�Wž�xcjF���	�������а�Z�y�nEe�Mۙ���฾�O	q�ps��x�I�i�#�v^����M��U�E|��j�x�Q�����1���MI^K;;����z���4�Cr��މ��:��<qx��|�^(�Z�,;h�jĀ:u2���s8M��"s&L$r?KZ��:�Zak�ZQ�<~���s#S����'�"d��ޅ\î�;�!�롂��0Rf�x�Bf��_�c��D�vMFM����ťQ_����m*�7@9G��=��[
++:�v$�~�)�D�~�zim-�����M�Կ�yH�d���6���2S���uC"��5���*vξ=��G�N���&��T�\~��mI%���''gǭ�o�:ȳ"�ȷa�~���Ο-,�ޚ��pJG7��3���|Eo��6��g�<���2�M\^}�mx���<���<��ہ#0"W��v���{�Բ�V?��X#z?����Q<�*�C�^�}��͆(U:�k"�;Q��8g�>���Bo5<ΖL|3)j�r8���k���L�Sp��u���4�U?���. ���$�p�'��\��M_o�[G�ס~�F�!�8�o����{AX��b�|0�)�+PLq̘�ۄ� ��W�JC���P�.Nw��cÕ�[)R������#j3;��|�jHǪ��#}��_����_���p��� g���|�n_��q����X#1�U������;���u3$		��&u��.x�G���uQ���Q�M�j����D[X�����K�l��(�;�F�&)ɫCU�i���˫�6��j)Ш7��$Ie-fQ�<&��;�6n��佪�zM�Z��?4h�fB�{��z%f�Y���~�F[$���R^g�<>����|���-?�t�2�J���mJ����h�K&��J�|�0��b��7�y��k�`}1�f��N�6\��!,Ck��ŭ�H�t�T��<���=m���:;�>Q�D~9�]�0&+���3������;�ڷ��փ޲�İc�G�)�WA�����+c3��p��2�GnoJu/�>�s
x�ђ��iwἰRV��D���p�p���D�/�\��:�&y}�y�c �1�c��%s�uثХj� �E�E\2k��]qܓ;�TU��/������;��i��E�6�/�-y��ɵn�B��wy��?��� ,�He�ٝw\�ϩ���z�g9X�&���\��uKUYb�ǯ|v��1�57�o�;2r���M��t��ޑ���K�nN,n���~Jva�ټ'~��C���(J�H`�L�}�tL�:��!�k|I�Oj�j-a���`Õ9����4^��3|3&��j���0='�ѥ-�y��(��ZH
���4��?=�g�ũ�/�.a���5.�@,I�"q��((#^W݃��y�/�4�@|0��(t�m����{f��e�%6``؀k��u�R3�N5`x��\|d�8�]�C"�K�u��؉T���ݎ��{aϘ6`r��W��$�F�Ϋ����'i0K=��A8e�^J�H""V��1��2�/R H�Q�YWO<>Z�d7`��_�
�yƃʗ�DV~
-W+9r�C�0=��[����tf�>j���q:A�]r��{���������3�����Ȓ0���j<~�v=O�z�3{��x�����{�`I���M�Zu�+"7_�����>9��~�`s�d���_�������죝�D�qII�]
�?Q�n��,��KG����.[����?�i��oT�:�+��-w؟��"�ȡ�{?�]������v}��zDҡ������~t�'g�P�k{m���#'M���k���4$
��å�>)���q2`g�/	��o!�.���Ve��0���Ua�`�	�Q�IC��s��)�UĐx��"y�Q�(O3!h���ȿ%Oh×�?�����T8�����'�-�$������9��V'Hr��������[�ј�j���� jj�#V������<)ZP��m3��9���8����qi�)��1�����s���w�X�͆�[α|���N��>0�+����m^���cՐ�"rg�;��6�'�~�P<�����O�.Ь�Cӹ�"��^f�>J6����;�É!'o��~OdaU�@n�����(GXq��Me��&x|9��Xw��N�~���?�G.�,�z�et����*��sP��tk�W�xǠ���s��ږ�8�ZE�&�s-�3�up�Y�?��63�p�ٞA{K_�_�@�w�lNMi���=y|�]��=q���W���{�E|/������j\�+�͏�l��׍j�&;�/�)�ڪ��'��,z>H,V����Ik�����-��OWp=�36%T"�[V�h*�l��8�D�R{��ÜM�@mTc|�c�D��{8�w���t3G�
�f�A}��?�<\���$��������]��i�P�c�$��_��O����j8٪1�^|o���)� U���^��7.R��>4������f�X�������T�-��Z�'�&1��;���ɘSN�x�W]���>��;��z�a�_6.8���>�:���a����d��OW�6=��3��
e�D�K]��������98 m@hb �x��Ѻ�u3l�ְk�/# % ��U������Ӓj�Ǽ�4"w��@�N�����XuU��a���F�:�#�au#���Ou��K<Y�?���5�|H5ݰo��N}wK�U��L����B�t��Ɂ����j�����p�P��A���P)���'eB�[����O>5���QI��>���5�o��x_+C�pB[y��/��Oϰ�52�,�7E㼞��%�����^��;iݕ�(�+�H�w�T���K6m����UTlyM'�p	�+$3ݘQ�}���\���ږn.��y�ʈ���g�w�f�N: 9p%�f�3�,>�~���y�1�Ș��D4�'�ߴ����_��-�`�8���p����:�H��gI	��GO��H%
 Qw������n|�ӹ׊���L��Wr'���<�J"�d/`1�+a{�]/���B�)b���>#�k#�*Š36O���8T�n����e�����έ�(�W�S��5�mR��7t��x�� ���J�v��m҃�u�8U���wIGG�!��g�_Rx"�Oc�\X!�BE�f������F'��˩ec�@���a�ZL`����,���;��c�R9Y6j�ʾ޷����mR�������2�����RGL~�:������)ͤ��\5E��p!fR�I%�sNAv���Á�c�|#>��y��K%@T�!�\��>p?�\3���f���[,��������=�r�dn7�R��R(�O��EOl|X��ez|��Фwt��Q��ɽ@��8_l�u?�Bp�?+g����"7G  ���޹+4B�9��N�J0�j��W<�t"5�Zճ?F)ޏ�z��{���~����A)����J������b��\̈́	�4>�Ne�����	��|p�k��{'8ݵJ;^���j�:~�ȃ�23پ� �>����Z���-~>=Y܆����H;�����V[Y磌�iu����IIo>���=~E��(M���"���[�j$TkD�:lݠ��2��5s��X����苯(dz�OSYl��S�xV&��n�������;Ɣ5qh���<�nXײ��e}�pƉ�埔�c,Xv���ԗ~�%���)A)��U]�;)�5��σ�9e�[�T;�V��,
�A�nqi��CW^� �`vy���U���kw=�e=�m��G�lִ�B��n]�[G������{�aV�FM'���r�WWQ(���_m�����lPk����!���+����,����<��Uc�L`�1�����[��u�q"���_�ƈ��>�!鋆�+S}�=�"n��H��F��1�[��t�?p�Aٞ��Q���s��9�v�aR�6`.NY��Z�S^��U�8���hLby����d��bjQ�O>���45H��]O1(�mаZ!E�:t�18\��ؚ/��Qے�P�KEF�e{��}y�?�ȹ�su:7�>~�7�%���K�W��L��Ν��9>�8{gYe��ǔ�ؼ���W�۪!4�^�Eu�1�P�a�T�2�N7'���D{�S�J%߱�����P��6����\�(�+ݍ�S��7,�-�L�{�@Y��i��nk,��b�j&V�����[�V�{���|���[�����5w���=�
�` �h�(M����Q;Fu9�$!�҇�f)/�T�@�o��doǲ�8� XO4߇`H,l�a#}ױq�"e[�4�^"��b��]��a��M����)�T��iT�dK��?�;���8��};|HD=Y
HM�1=�7���f�b#%���i
�";�)+"�p�%� �gt�|2���Pdh^��ԁ��q�x�����,o�cm��S�XPc��F�}�~��/S�wҘ2��:�#�Mz���`�(�������,�q�������|����%Z�9��)��vq�K�����\/O����O}�_���M	$*���[����������?<���6�bŘ�A�eo�1"�+��Ēj��#��[�GQE�ͺ=�-@��o����~���;�LO�J�V����)wL�r�K`0�,rR�7s�ȳ;y�@G#!�l&��?�_B�1	-����-�q;�,��P��)�ii)E�-ڱT �p�O��o�U�Y�G��j�!��ڥ�;���Mzz�-��)�����*����|F�@g�����������RqR��ޤ����*���1�pE����9�� h��!x�G���K�p���}�|8�ۋ#䐦��G{����Y&�a<C�U�|�ð��b@��'�<�8�鲈e�v�VI��)��?�}�ks��m��bU���z�=Wm�Cj��u�5"�}�'�y�%��*	�'��p"O���}S�u?��Dƞ��d�3�H)%��B�Y)-�~�߻�/����W������_d���o\wptX�7�r���q73܂�h�};2�$eK|	��UuY��.�y���:������,�iqWxg�I��+V�����m�#1�x'���7�#�(�
j"q��V��нx÷�P��
��i���ix	�70:���'2�{�2h�&1�c�[�0�E`N&�6ְ�?j�앉��hxǈw�J$£���c'�m�>0iTgQ��%�Z�z7��T=:I?�����{uO�X�0za9��:�凿%��p�Ja>�#�I����8��n�6"n�����	vl���K5�*5ty/�-yrA�ܪ�Tc�[�#ñ�5��q��q��N��3��P �Y�F��+�z�Κg����3ˣ����K+&����S�s��ḣ��2�V%�IV|e� �l�s�ܻ�06y,�[��U0����Ыe��yE���Q�nJ�!��30x��u��.�����ީ��_�Z|���P�QQ��� � �R"�-�4J(J!�0tI*%%H���0�ЍHI�C��}~�^_���s���=j�5(��.������(\c5^SF&&w�*��"�/#�6�o����(��f�^�Չ�00v�lОE�}��a����������S���L��5zX��Г�^=�F�|l��+�#j�����$!b:2gџ;��P+�1�4{�%�mkrk�WF�iT�N�*��Nb�ٶs]�s�����cBX��_�}�xv��9�W8��Z\|��Ml8h��qϭ��{�l�팪2w�#�&�|񿞺�z؅�2�:|�?= >�D	uĠ:�8|t���7Ζ��Z2�ٶ���W�3 �۴V,HN�bw�����Z�P���	u;:�l�я/�7��!�h�a'u�'^#m��Gr����=Wj�.��s$3���L���eb����\���Se�h��Y�cO�1tl&�Yqr��^he���s!b�A /�N�)��e�5�>mk��$a�P}�ֲ��/drO�"T:�"����<c]4�?K99#ј�z�)c��hi,�ơ��-JN���R����q����(�1�8}�;Ъ3�O��\	Z#��1d�	e�s�ݪL��mݬ�m��^�	�#�,��1���+ ��!�5\n>곑��S�34i�.}�%�����콱w'8%W$łe�v�&t���7�3\��5�}aL�Ò�@I�!?�Yt(N�p޺,Wq�?���a�{Il�Q�]L�����>-���f�T�/;��u$3�)����~�k�=��pV�7Z9	�d�u���s�#[>!���P[�m=�r��F����T�S��ӶMW_ϙ��I��a|q��o�'�̹ٵ�I��4Q�;cJ��7k��u�B$�M*yV���U��U#�P�ϧ���L��.��pIi��C:��[~��9 ڇ��[���,��V�s����}��l��r�v����;�F�L�Ui���9L�Ϲ5#� ��8���~�����y�Sѿ$V߅��	�l�Mg��{`/š�A�rX�㮳��tx_�Z���R��'�~��l�S���TCk�_�)v����sĬ���E1��M��u��}������A�� ?����[Φ��Vͣ�oF��^����{�,5/;���x´f����O����o�X��*�O��g"QL�������gK����1<�ױ����s��I#�r���NOڈ�4��*�;1���@������l�%�{cm�4�<�<�}F�~}�� t�qQ�B���&&u5
1Û�X���ف���Q��PW��B��T�����#>��(�P["^:���1+�G�4�F�������&P�zQ/�p�=����M��;3���Vûi��:/�;���v����A�h��VKC�%�9J�C�V�����+sg��c;�/��#��{�A�Śih�]��-��o\C�����KN��'��F���?�����2�ly9\�������w�'���3�$o�f;@˭Em\>�]V=�﹵����A�;�b㓸m��ڲ�\d׆�S(��l^�yfo��7n	�8� ���
`ڗ��R����[Ӏ��*��ο	y(�ld�������N�Փ�/����{�>�8��^|8}$=�v�'�"�Mj�@��b,�EL�nI�Pi����x��On*fM~���(���Z����K�qv7��~ǹ;��gn|krU,�<�/�[�5o��;�O��}M"�Q���nw�a">���l��t�x�>�bC��G��Z�U�\��s�����k�����͜?��~�!��i��g>��K�r���:F&^�[B�2�7��54
�	�i����J	8�݆���d���*i'j$ĵeZO�Zj~	�{z6���a�	n�w���u��$��l����iJm���j�
��J�!ވ��i�I.�W�xw��`�{h��?4��v���YFz�M�W�F#�<�&�[�;,S�h�q���]�,s}��4����ߩ~M������'��7l~I{�3�
7ȭ�|�y'�7>a�n�fw���z�L8utB;c��C�$y��5����_����Ts�ZzcY�4{��L{�֘x�&Y�y&h�y���SO���GxV��MXp�B_޻^���C��r}.A&�#��|��Ŝ����rň#T����1��vP�By��$�O揠_�)��������M�_�?����1Y�Y��k����?r^����wOk�^���L�l񷩕r��9v_���`�&��a��`�e�x1#�Pt��ʽa�����8��.�x�����)�G�֣Tԡ-�� $듕Au|�� $^~��ȓ$����?������|/�Zb��(�-��"��9�&�	��'�c�_�h�	�f?�$)j@�pWV(B��F���
�Ю���x��n+GTRx6�5Ο2���3��~����}8T��2�u� "��}�}*A�A��,�}����g6#?��ha�{A�6�a��`5D��Zcy�?�M�f8}��4�ƴ�!a�EУ�2�,��s}�
Z#�`_��s`���w� �N��נs�vAZ~78_WE
�ˇ���_LF���A��cd_"��d���i���ﯳs��A�ɬˤ��=��#m�-vi�掎ͬ��a�ۭ��;����ļ_Cz���������V��7<���E��>����x_�ul�S���LR�K�ɶ!ݼ��㦲������̄��SÖ6>��9���T���[�gd��x�8�&�{��1<۹.y���RB6��c��$���y�p{�c�� B���S����a��UZ"�UdhەK{(yO��%�T/�^�b��v��{4����՞����+�t}^��
��K��oqlS7+7��"+b#*G.Xb�N����ݗ0�:(ט�P����{���6o���>lY�j�5iP��[�	���7��jܛu9kk�P#����z2"�l���������P���Q	yt:�����z-���	{T�-R���?�}��������'�YW���In,�`�z�����l~����������a6m/�����K�."�~�0.코d*�7�{�!ҷ8sL3���BD�&q42WR����
s��{�Y�~��ȲD),O���on��=vXeb���kI��|��e���D��ew�+���#�87"iz��l��\��K��SM��Dl��y�xySMT�uE�4�.�Ӭ�{Գi�ګ��Ɨ�Y��z^���j���y��� ���bs�0�"'-�S��3��ƨ�,��z���s������(�������Wҹ���5){O{����e��-�<���b�,��#���:�����.`y�����!�Ћ3U��z���(�Ь1ص�h%#`��d֍:�x�T�Q�T�����X�����[�I��B��.�f"͂g�FnL�D�m^D��wQ����+�d��-�hک�� �NK|�I~��p��:}W�$�nL �lY�.�i�lBL�<��a������Y��H�P����׾H��7I�塥��>홰��,z�W�hv�-����q-���8��g�9G��<�Jnu��s�t0�>S�"���f�R����3��8^���g��^���`e��p�#�L�Z�p�	��h��O�EW���^K9�R%�YUb�"�j���i�k})���x�2�>6Λ}y�� f]�y���	j��H��\��[�ְ��3�O��IδDc_��D��⾠�q����α ���\�����?"�a|B�Cl���Nv#�磣���k
��ѽq`����ƃ ���H��2ׇwpg(���_;������~K�nوt[}|+U	~r�b��SgfW[%��k�,�X0��gS�)����s�p�m�7�ĎBB"�z̭&��o,�x��pr��8���V��b�:R�N7>~5QjPv�p�j4d'�����F��&�뵦R��jBa4w�O����_R|�t��@P	M�0��>}]�E�up���м+k�3F�x@�>�:��w�*c��kQ��^�HX���rf�_D.D����c�t�%�c_I��!	:�Kd��R0̹+���\n�D�H�3�/�y9��%�軍�nw���l<�=��K����9R��G�s'o�M�zv��܅P��>�� ��a��_;9��[�5�����P����͞��Z
�M5`3��C ␻�͡�-5lK�ȋ�����ʼV���ȬT�/�q	m�0g~��g�z��&��=�E0�;G�^TM�y��!j�����+��u�f�n� �5M�F�N�.t-IC�̌�5ń)w��4o8�J�%$BiY�&��U�L6�N
�Xu2[�oB$�&GF������|[��a�/Q:��=� 
�`^G����0;���#]O9I
��Zԗ���P�?�U��7����w���0&''Q�v����\�0�v�H�a���wL\&�m(�K�5��ڹg��q��)��6���e%�B{���c2�[::���R�2�)8�f�>�a�_j���c��ٛ��l�[	1�?�,'�^�:�'�;��nR���ެo`���U�2���;z�]����=و[��R�P���m����(u��2���^�K�!D�6���Ez�����K�� A���QW���Nu�{�d��c�a�1}T���1��n�ʸ�E�D��l��w@�����0^T��/>�+�تƍ�aj7�r.!o��ۣ n���#�4��[�&b���gё�'��w�ܴ"�2�qk����	FH��wS \XRoo���ۍ��kq�'�>�e��G�o<�T ��,����vYa滋>�ׯy����h�&
@���$�����t=�a��JSB-��,�y�~@�_�ەD��|Az��x�e�nP#!�x���ԍ��O�ufA�Ɩ��p�*	�&畜6�N��i�Kj+���X�4���]�/>��o�M�xw���c痩&hX�����D�N7�l�G~f���2RFդ\�������:�ZY"
[KNҭ���§)o���"��M�/���@�Q0q��*��j�@x#�:F���B���X�t�H���_�W7-��HDF�10@� � �^%�=���'w%�D��\E�H=�`S��Y��~u1�;ܳ��t�	g��/E,n\�'
�^�6�Ab��`9V��&z���T]���v�Z.�g��G�|��q���Ty�:�i��*�-��f�G	����z��]|��8�
�w�M~چ��ۢ�S��ax~o�s ��#�)1
%��W��yu���vF�"k���b��F&��i������VmV����&��Q*�γ?g\�����y"���iˍ�l 鰰��<I #1� F�\�r7[:��+=5��%�E�)>������M�ZK�>��v��W�̼b�`jc�X�Q2�iߋQE��S�H�߾�a�3������z���՗f�_]g-Q�n �7f�ū�� ��M��DT� � <;��i&�
\��}ԭX7A3_��G��?ۀ+¹$�EHQk�%��L�kT��nB��9`A��c��'��7��Qؿhc����!�r�t
�8��Īy�� ��@8��<~�����/捒�j�#��6f��@�G�Y�%��4l0a�%�E@=+M����s#gI�B�[I�w�&�)�+�������[9�G!�-YU:_ŚwdP��C��T�
����y��'�z�>�Dě=���3S������C+���N0X+�Re��5yM8�d����+�4]]���z�f=0���x��̽���ϊ�~c�ӷt1o8��3�J�7�`iz]6K�C(��RjB�u��\@kߩp�<�"A�$��p�_VSBlX;E����a���o���� ��8�e;����ݕ��a��s'�B"�]�f�F��a��ܝZ�g�r���]�2"�.�RK�ɘ���&� r﷢�$\n\���p׷|KN����c#���%FY|���g|��@����#S]X���H�9븪��a�"��	�3�1��4��ɀ��z{��޷%Z���4���b:�PEϵ���aAy�X�w}K<$��A������R�;;sVXd�9�����>����8J]@�#9�-�^�Hr4|>���s�-�G�.>؊Dܳ����̱�z4��=P�Ǭ���q8s�Z��@�^���	j�F��~8d�4v��T���(ʯ��')�҂�~O�� 0���Yhw��/�Y�o�M��޴�Ąs�&X�ljF͎;�jvm�h�Gr�*:�o����E!�Q�ِn}:���%��O;wW��%�Q�
iי�c�&�s`Ȯ�n�����̫�&Ő��f�cii�A]e �v���nQj/_�6�2b���'�a�Sצ<�H��Q<C���;O:���p�mh���v���T���|M�����N쫞�}޸F�!��� D0�Y���7�ﭫgVU��ܥ�4��"j���,hj2sc�"���1����eQ�{�����Mi&���{��b��(kl� �zP	�d� �k�Y3�q�	�o,��N`�E
���1gy�2�?�!]��V� V�L�s�61�� z��80����0���:��7�D�cs{;��{{�,���� _~�Y+���?�����
�X{���w4��3��3��;}���Gh'��U1��@�-@ӗS�a��Z�^ޙ*7���u
����s������gt�uS[-}�����6��9	�^(Z�Qj�y��n�b�jfW>���p8Y��u�����L��ϵ���{��:���g	=��  ���=&�r��m����g�ǳ9#��$���}.�q�����8�d��ŸŬ�u����D�{��%����wHnH�������k��뵁��L{�����7�"�z���+��pu�C�dc�趄����£�$��A�!�I�~x�MӔ�ǉ�YK�Or���޹U��O�-k���:�ce�Q`���>`�
#��s�9g���,i���`x��簴�+��. �|�z�ǣ�O� ���� &���ݷZ3��	�>.$u �tgz���dg�m���sf���{�-��4��7�I�j�/�\��LUᛴ��ظ)���%�|:sMl�.�b==�����Tra"DڇL7���ۣ���bll|�gk8��r-`g��=��]e�:�����u�����iO�	���qjg}4Q{Y�̨tN�"}ǼT|Ǎ*�6��a�*
7�6�0j��E��d�q���c5�ќ��ȝt�����(�ܶ��	�!A�Iv��v�a9c/���(������n�(�&���b<2B\��^���=Ҍ��k������x� o����i @���$�� ��k ݤǮh�=8(����(�MN*��	��a�Y5��j�0uk��e��o(&�/rl�ȗ�x��/��Z�y'�g�.Rwdb!!�+�C!�γ�N�oH����1_�� p��/9~�Y��j��8N�����.�W�@c4ǻ+�N�m���`iCxǔ�n�{Ev�ۓ����� A����,�P-���x����Q�9�~�����\J=&a/����7ٺͦ�԰ %ſ�V@���Ҷr�l(_�M䨆R�=�~Ni���=��>�mYʚ8�s������2 dl5�N�4��/�r��)�P}c��C�����3�h�(����5��������4�x���pϿB����GJZ�j����%���/z�g�)z�Zs=SIy�	��[��s9e����2�Ł6P�+�ɦ�G:�|����{�s�_.:������?���=ʤ�P{�r\���h�Y��nre�������2,7��a�A#��K���xH�����Qg�݄�^a�#�Z|��֌5E�����A;F�H��wD�z+#�5B^�Χ�
���c��]��1��~����9�:e�CV�L[~�խF�aj�g��ck& ;Q��n�ӑի�Q�>�մ���2�O"�+��sX�<ｘjr��>��Jׄ�UX������\V���ˀ�]`���*����e�9H�0����?"��SHq,�ɧY��E>8_��z�'��]|����-]��K�H�h�'�0������<I�r���wԤ�glp�|w�pZ���ȧ��C��ݰ*Yi�n��<�i���E5S��L[?�Q����i;#�ϟ?];��d���𷷷�<��3����)��$��a��Ȧ��]-ф���U}Ҁ
[ۿ5�S9rp����z0�Y�Ko�!��ԬS{U�y����$�3"+Z�os�N`�A�$�ҷq�|w����L���Y��^踽AZk����\Tdd�ǆ6���W�X��w@q�/5s��Or�ij�&[UbU���N�SƖBW	m@7�|�Sl�)�����ᛊˤ�}���Y2�[�YrM�$kq�� }����l�x <F���>a�w�����; **���OR
��<F��z'�]��R�e��V��G�
Tb�r><���ZI���'22�*-9-R���k*㻴���hBm��I]��� Z��|z�<�@Xȹ�'�.
�/�jG�c���,Z��D�ƼW�-�H�.�wjYx�m8t5�Wx��b��f�@{mwAY^S� ��:�ah�^���i�ݢ��r>�Pi4 �)�c�khT"�\�q�����hGO�v��Kǅ`|����H��hn=�"��/	���"t�fڱ%�Q��|�9~̳ܵ�� ��8BxO/�b����[*d]��ŜkQ�񰴞�!4��ss�ewj4u��u���h��{Vwe�$�9�E�X���>�9���{�U�hC'�R�����q�����6������{â��}�.�P1a�ȳⰳV�x��Y�H�;���|L3�����y?�W h�'������nf�uML����Ff��p{����P����ř<��FV�C��ca'�&(����p�ɬ�s��7�ϑ�8�!�ok�LoKP򽿪q\Oz�C�:���t�@��?]Ƹn~|s�˻��i�Ա���.`I�z���	���]G\�|�8q�����B,r������Gu��B��15�dt�K�|@��Y޸�P�d�c���,�����VRڿM�a'�y��n go���>���(3}��A�-M��#� �k�!S��U��r)��R�\���ISi���%���Y��@(FY�rV\���1�$�ت��(��y��霢�����v5�#2��~��M�B�~�q���4�F�,��� �9�����'~�x'8�Q��:��sV���TJS��v�p�sUd;����޼R	؝N!�Z��G��*ρ57��u���Kž���C"�3m*�Wh-�H=������\J�Y署�"��3a�x�I�h8h�7Α%��p3����[��t � 9f1�ٔ!�g�vvܨ;3(©��f.�+M��~3غ���1񖸻{��j��|�%��NoG���M�b�c��%�?�9a�A;�PXaC��
��.�p�_�
B��M�Y�Q�1�-����AGIEK����r� l���&^����B`��05���.g8T��l����j�ȉa�?10��@~�q�x���C��5�Q���O�ݦ.IA�IȽ���|.����0ʷ����h��U��������	���gѮgי�Y���KB�W��[��&�]4Z��4����(�B��^��w�!XR��������p��n7y3��m`������IZ�OШM}XPc^Q�GHB2��]�i�^�3$fz�"�˟PK��a��[��e��ȕ�kԁqQ{'���`�Uy����h~\���G�!U�UV�$轴 P�{�T�>�ٟ#:a>��F��:,{�f.�|��l�a�L�g��z�F~0b���얆�8{h���q��L$F��22�������2G7~��,��:-E�vJ<:�s�C�>b���j��j����+������z��m��T!9��Ea`��7�yZ���DU~����o�Ht�������]�������"w-x���̺��ʶ[�� �ӌ5�\0���	��/!����_&"�q}(0�,5���_���	�q����H�����3���XX���ĺ�Ԏ�ʄ��S֔�;��A�3���>!��djEF��/���@�1�#�o�dZ�k��]g��p�[wh�ZJ�] l���^�P�E�9L�H�Ѻ�ސW�P���[3�^�s�������c�|���-���1���0��'蘮ʝ[׻b�>zm� h>�V^��a�J�^���:�s��[�įu�,�'e��f�a���9ˆ��q]�,i�M�@�8R!wn����l�ov�;��z��TX��A�
F$���3��T			� � ��c��1���j��T���ü�K������up���CJ~/)�V���(��/��)$����}PV��S��s�>a/���g�ȅp*��oj k!���/��w���j_�n+��=7ί��%m[L @�����k�v?�aK�=�����N�ؠ�����v+~�
�3kk��ʾxFiR\�љ����~�}:?#&xC4���%��
J49M���xƂ��U5��:�0��K�>�f�j���5P#Ǎ���!�<!�mt��C�̇z�U��K#7^^Y�Z3���\<<�&�gF��bmr|U��?k�=0 ��&ۋjXr���Guu�*���q�??Ҙ����wl���e#��*RL���C����0���h.6�0�����@4���[�h�02�g��"�X]g�Q ���l̘:q�&B έQ�_����/ӂߏ��j�	 +d��lw��
�߯��9�7���n��u��k�?:>Q��7�0'��:�u��$y*P����n����C����g��a�<!��4�a`�2ԮDW-�'���~���t�|��;@�Y �ִa[�����Yom:˘)+
F�S�90��e[���F��b�e�6d���@>�G�e�bW��;��4��`��a���̯� �0'�l9��/ĹJ<��fYf�w�!u��μ��
n��`�~��l[����ՌG�!-?`�Q�>?�;.:�$�+98��]���vQ�3��T�z߷.����N��OTSْ�'�mj�?��9[F����C/����!	g�����ub(l�70 !�����g�����cD���m1.)�cM�������JJ�.�Q,Z��li�#�Q2���ђ�>ƭE̮z�{����VG�f�����V��x�l����Ą.}�!��-����VsX�}4�W�w���5A��c���f��hGƇ��}5 {�<�yC�̀�9=�!�`:`��sKj51�8��l�~�h�=Z��xX� Cͮ�i� ���n�4x2��"��-nd�Y.F�S���e{���?j�\�B�c�E,Lt��X�0R�J�����.�!=�|�R�`���9��Ġ�1W�+e�"�\��ȏ+|ځU�����)%w6�i"��������{l�z����}Ԧ�$K'��qx������̣�cz��(&?�����g�֘���Y/����rI���g�f��Rj(".�z��%�s� 2*
P:/��@��=3����(@@�l%'|	\�n�@P�Ls�nK�z�yۭd�i����v��t�[|�橛x��n�v�wX� 	�TKu��4���v�..}��}n@VȒ��/z�&���Uv��Ӗ�EZ�`]L�t�]�P�>����Մ���w�H�4�$�!���Q��j��c�ȵ��R�9�B�2�����%*
*v�%*O�=M���b7��k�}�2�3d (���n�3��m���v�b`a����my{�d&-Dؑ�>3��91�!��Î^���?%1��ALgko߹���d��km-��Ty���N5�D��4>?KQ)-]�\�~��_el�~MϺ�1�� x�vBO0xem Y���!�:<.��X*�c~K8LW�4y�T����:+�;Z��Amو�MiRI��߆�k*yټ;��e�0�1R.|Y����[�p������Q�YU{�'��6�Oϔ���1r�����NGz-wF�l�;�:o��� ~�MQ����7����?ޔ�n���X�/ފ��NS��b f#;;{s{[QM�
���`���C:~Y�r��>�&힟&4B�Wq�Mu�-�˭��n|j
��R��!���h&%�k���~`+�e��n��]ޓ,�٘ʸ~J�!&�h��|{	򿻸�<ۀ�o�՜w�.#ro� ���rFF�M�{��7��y���vd~��|�����"����:�"⟹v��	Jt�����B\	��07_:���P���ca f��g~��'�G6��kj����<�����v����j��$v��s�I���@U뮯#�?:��CF�#S%�טO��������q�c�L�Mo,��V͏�V$���za��/9��
4�6�/z?w�Ċ�v���h�Y�2�O������,U55A99����";HB9�ϭ����2`�l�
�����Mc��%���y�w�okk��D��(9Z��Z*=##N(ţEv���?`JPv���'�f��-HʧO���sXo��]�z F ����T�уl2��Bw�3Z�����I=s�H�Є�����"��J������Q?�d���G�!�U�Ѫ��"���B��&9M__I
 �(= }��-�)�{����.ˉjL�&���{�(}��	H��&O���!VR\TQ��bi��g������R�^7߳�1|rX���uf���gxQ�8�-y�8���.�xF& #sX��z�Zp��t3R���n���ˆ�:*<0�h�@�{�V�\ ~���SB���&b�?�W��3�贐���Eǝ��M���n���9�1`�m���qt�n�3��'+]��y\�	<%��7?���z����*��@ش�Y��{��*"�15�o/���X����q=8�x�탨�ܖ��kd,?�1V;�Lw�P�X�V��%�}'DQ��v3��E���A�P '+k�f�@.�w�bo�m	����t�!��-�9�iq8tu�	L��8v������*�׃%Ա�v�^�w.>��k	>�PJj*
}Ξ!u������S��ӡ�m��^�13w+�(�
LJ4�>�	���������f�\>l�szv����//ޛUl"6
- �[�*v�U�i��z;���j}[z9��yʇ����d?�)dlL�z	G>����qſ�:��WZZ �8�iUE::I`Y��	Ø��R�A�旅��υj%���{^�@�7θ�w��:�8��#��oO�r6!�~?o��/���U7%,0��ծ@��ݓ����Ɗ����kh!����<-����`L-��
\d5}0<b"������NQcx+��� ��.��s�	��v�-�^�������R��}�z�ñ��Hb�gX�ueea�z��3ҁ�:�)��p�ߟ�k17x��#��l�M�3NW�d.�!�K��Ӈ�󀠛=�q�镯�����J���n}M�r�曱��:�h=�L��8K���`ߌM./�� �m{�\�,�c<��be�y�r�C��)&�Y�����ʼ��6����O��+6� �w���t6��Nϖ\V@�zѵ�R���p�
���= ]`�DH���6���Ug��t�-�*G�2����l	���|�[�m�7��y`�]�fl�=9��/�'����e�/aiD�eDǝ��M����<J�5�O���+����Q�d=���� �r�t�L��H�ï�ľgVY�|�c��D̥�l"��!��/ pn
��-HU��gԳ�~������8U"Q 2�׏��Fo���i����� ƭkcu��7��B� 2�+��g�QFei�����T�j�%�����4E���c�t�RV�������Ys��ÿ13�8���p��;�	�W���/�S\��R'�C&�����9�3�i�gg�Zb��2�#����2��)�T[[���N�f�/:�Ќ?�� ��b�����*��1�v�(��]����<
(��Su�B���ؿ�����]�����#[��Q+��?/��O�ڒ+tGe�!�y�0���gX��20y7�|hHNE�u��Vr�/2�&���n1I�K���F�g����"w�ܜN[�%r�K��vF���+9���+�����DC����w��=>�,����ʪ�k���q;�[�2^J�*A?|��S�����p��,>A3��o��IJ/C�;��D��ٟ#��@�.p$B�!���l�pש��t8���kM�]��a7y͠�����V''' we�:X�)��Q�n��2�Qds���.٤1f8<T�<�c���`�
]9��J6�##���o�.���lcNT|���&oGϞ0�z6	�]�*q#y[~�C�l�HD���}���DRNߧ���
��|������������
�nE��@�����U\��*��sL>V�q�^Q��B��s����4�غu+)E�x?œe
-�Y"J�}㦦�<���yï�܊bsL�Ē1�H䁜;��'nSؼ\�;���Dp�����{5����Q�����7*�N��Ɋ9�6�ea�m)K���Օt�pN�^�*m���P�0��'ŀ�j�NSJ1��}��1��y��
�a'��u���V8��{^G�^7�����P�ii����8�$�ɵ�9�[��h���s$5�A�"W>�g��?׸p�³خ�pq(���U��\D�I:=:�8N��?�z_&@ajk�]�B�q��|Kjii	H-^C���J`��\��ѿ��1���A���>��6��=&���n�����M{�j���\��A����.g�e3�I���/q���a��aq�7��Րϛ�/�#
���[h^�`9G��;���!	��s�gE�r�\/ (/S�j��5�,�����ߛA�}�$�z1�0))����
�4J�fB,���Y�?��&�d�E��<�ш���\���.y���`j���"�NU4G��
[4�tD<m�A%����QR��3�8���|��3Ab<s�:{������pZH�#�ٻ4�
%x��tȟ���3����o�(n����oPy�����e|H3�]TRwݣ���}WT�UW�����X��G���~����I��KX�)�#�I���{�}e��SF�����E�?��1M��^�1:�3텑���<}��9�/ƅ�yY��}�
<���o7�vE�!�A���5F҉���%N�K<bf��P���N�;0���*�wۘ�^S�.�妙4ʗ�.m��:<rt	��Jg�I���>��,�d������\%i_=��� ���4�y��3�����|���x/���h�-�I� !������S톁-@�GG �z���s��B^��u��z�;WgA�=io'�<	�k��ГAȑ�[�B30�3ꀩ2o��pIaFE�����壩�� !����0u|t'z��,���xM���"�|�)�����=*6�:&f�G��m�_�.g���H�n�m&��&�lV~�!������=%���s*"x��2��ߘ�+<����c���e������Y�rߏރlLDk�ࠋdu�#�F�.�x�vʽ|����A5���M[�4>=N6��@Q�� 韲a%Gg(�C�p�I}r3�q�^L�iǲHMH��m �{|O]��y&/nt����˜,]�'	��8��vj�����cofNf��%s�"��n����.=_usb�{�h����6G/�q�.����RzL��m�Qd糙u0,�(*=@�fZ=�k��v����^�s��>�'��#���d�Tj��<]��:����N3S��uŔ�/ßLv~[z�e�Y�T��^v����Է>�<�<���U������;���Q�{}�� q�!=i�jUp���������hh/�WG�|]_��`�J̚�C�o���ҒxQ��3��V`��C1P컑�	e(h��W��}t!K^rX7�U�&Q[*�->W�g�@D�&�{o.�������
�3j'�#��yqjm�g���SW	#:��Ej4���3X�=��w;kb����2�MJ�߭���}#�H}��iY4�bz�7:y�Iʰ��H���ёp���|lb�!4�q�[AnKwO�#A�V�
�<KJYF׋���Օ��@��ä���)����#d٬I��ԨA�jXtv1���L9�(�������O�c(w�6dF�+)�h�����u\7g�^.�)E��y�N�K�V���/<��Ǿ�W��(Qz�����;�(ʻ��8m2I�\(�<�:c~@8�w
r7���o+�_ׯ s�8�ҏg�O�u�4Üמ�z)�CR/����s�	��dk��a]�����+湳�܆�Y���$�h澩��4�ݬ8���nҜ��>=u!,��Bn#�3�s(�~t<4Y5�.^�uv"W(�cֻޅSآ�~���{����X� �eח`n����*\�É$PouP��c��?��n|����@����Q�.b��}���r���|��Q�����0����a��2���M3k��wE0V��G���	�b�lS���b��&���TI .Q9�������J0�Qw��&^�/C���Ĉg��",�� ���2W���`�U�>땻����,���%�����|}d��� ��?}�Je�)<R�R�Xt�0�x�)	��(e�^=��� �p?������-J|L��Q%F���?�'І��������'���E�����*h�s�]ٙ��� f=®�q�8j� =0w�[��ӨB��H�C}�	��љ��~���|%>�<��Q���������k�;���n�HiҤ)H���&�w%4A@�� 
R�&��� ��Ih�BI(A�=����˛�a�F��{�9�\�����ۿ��<K���ht.����"	QN�*��p��)�����՗R�ݽ�$}���/�u�f<�����c*4(��4�6@�`<##E�{08�Ϯ�$r�Y��Uc���;�l�'����%���_��^큳��v]��n���g�Y�>էy�O�lSW��u[i�S�zJ؍l����p�l���g�޻�8s&�[����ZP�U���>�񪕭�#;9[T��d�h��Q�#;���`���>zT�W������������o;d�
aI(��(�6����U#30׏اo)ޛ>��;8zfs��"�nf4[��Eӽ�!�^��M5!讷��.�e�h���6}d����� �+ܷ����%���炣�WXnP���gJZso���}������η�����=�rk�������7�,Jݤ�ކJ/���������b�nBk?�X���o��j���}�{E˭�� �`ŋ|��F�2�u<��ci�-A�t3��4^O�Pؘ�;N�u� fbW]�S�V��8�6��|����+_���wmxO�}�2���>#���Cj�0��F3ڗ�;lV���:{�����\��R��X���3�<�uc�nX�)}V�
P'��՟��C�ZGa�:���瀑ac�sw�p��k+Ò��	5 �`G��T���K�����w�]�6�~��1򼆌\A�f���:��׮���
{c*�3`w�t��EbG�]E>�׉nN>�~ȕT���	�_v�zz�j�>c�*��+��Uv�r���C=�8��mb����6��+�74S8f�M
˻0��o�����O�)����ɤ��9��9�� z�l�����J�a�������}����K��a���x�7����)i������Wb�+��"?�"WR�14�G/y��~�D���	�l�D��O�*�D�������f)��w>��
 ��N�~��nc,������$�\��$�R�
ѷm2 ��h����y�Ω����W2���z��-�/{SQ���V�+~v�bշ�d��\^2U��JR����(���\Q>���T��X3���1p���aER��d���x�8x�=��A��J�R*3�7˻�ք���<_PO�sMX����X8#u1��������P��OA����͡򟋧x�%�ºOw� �Lqɩ|�1/��wT�uG�ֻT<��>�z2K������-��z_�pڔ��I�)?�E�C���'W˰����%�y��m"0 ��hg�N2�6d0�X�uU����<���2`�6<����16�F$#1�l�#�;�lI�h��źS���K��K��Ffg��S�; ��u��`4��N8j�<�i��C^�-�O�X�M�n�OA�2�\��x�a��-��L��L��zqV�xH�x_ ��@��W�^��'j�����g�r�m�bً��eڞg��H�D>��ޝ]9�zB�(y�5_1�I� ��r#�~��O�#ۃ��������T��zߛN;�˳����4�����C��CNO��`Yœ�ĥJ�$B�3[��\{�g��\����zE����6F1`5��4,Ai`�_�+�':���p������e��1����ѷ2���X܂��'���J+j���Ey��{��U6p�B���t���y�~\�\<pށS·��" �w`LޙM_�
���X�CEa�òp�c�[�xk��UP�>��qv�N/;��O;�!�L;%0ڑQMC_���J쏨K���ʹsڻ_)�]�ԥ�N���+�J �*�0�(K����L��#5%���V��L�jn�bއ�[�#��s��Zʾ�ʹ#;h�߿"}~pɪ��PhO�wP��s�I��UOk��.����V�zaQ4�iַ�&�٠�2��Y��7h~K�m��G����W?�g̈\��y��-ғ���؜���/_EMkc9t�Hi.@�7����+(rܬ�`�(�Au��R=�,r��ҤxX[����͞=��7��S�}���4�Ō׾d����ټ�y��� �Q}Z��=#���U������O���oayQy���dۢ�[~�q�=<�{y�0[�S���7B��!ݦ1�IbQ���p�&Q�}�0�9)ЈBa��� g��v6;��0���.ϰU���o��'?�/�?Q�8M۵���b�� 84��P�AIz�tj��f2�y<x'$ȱ���$u������_�3]|����f�ѭN<��xl�|�s�Uty�}?+��Pp�(dS�ЋM����^Rq騏K`�5dag��h�����c[�לa�Ls`�P�-��Ԯ���3r�@8�B���9����a���/�%�<aS�{'����P-�?�)(�L�)���̦��@+����g�	x�����T@n8m�����k���ƢΉ����:��&~�GA�KCd}ξ�i�{%T���e(EN�,z��}���&O߭J�?��O�4b,�������������7��p\�mmgƥ�s;����\�^���0�.`��z�x����_>oA��n`n.�t���y+l�kv�萫?+߼o��q��?�G��ƭ�GA�A��g�r&��?tƋ{��T%����߈)�ٮ�_L٨٠��Wy/�y��}�pPab%L!�Q��/U�n	f�}�5�q䟻��x�+�<�q;l b���`n��v��E�b⻏��t|b"���j�Lup֋>�s�N�Y�nЯ��i�.pL/�r�B6����2��@�c���.��E���,���������w.���z�{�,�Cҁ�FG�mUb%�O;>��kb �O��犹�`��BS�k���k�Q>�޲��9�j� �߶~�Ŕa������ƃ:U9=cɤ@uѤ�/�/k�����BHݵ���#TFs����=��������/�Bq���ӎ����Kh��/#b�����F��ſ��]ئ���}����uf���%�˄�i���n���-�'�(�R���7��NO�e���b��rZ�	��[=~�_�I ���Z�QWx��ٳ�z=��|넘��R�t��4d%gw�"> �ʹ@�9�+"�z�C��7�@�ˉ�*ǀ��WTQ��Z���ѯ��5��zZ2�E7��[�}����-U;��'D�&hd�KL�˳[2q���1��|B��0�|���#�Ώ�2��JG�r[^;�怡���S�ҕ�#}R3�q�	��Z��ª����n���ɍ��d�PV��t����6:��z�d�m=�%���y3��X
��z�P/��51Y���b\||�p��P�$��
�j��7��^^c{�u��u�ן�U��d����yDC�#?B��X�8���!y�L��$�ρ���s�3x�d����?}=Uz�,P�\��#
'���fl�ή[���{��޴T�O5�sr�@y�;!�����s���@O~U��� �8���{���=/�H�RÈ����8���IYe_�aT��cFe��T��ߊ��A��~X�����#�*��).�c��JFl���2O�\m�ؼ1}☦�t�~$+����8m��?/J���1�%�p1�Q�E�Y��~�Hv�L��囓������p������ʃ�[*�5
�Ъ����pO�������Á�K���>����o�
i��覉UO�3ԸH�_[s"�D���wqw�tM/��鷃, o���@ؽ��XZ3�A�U(v�y-�n�pTOg�U�����o����w;���jE@�!��U���#!?o[R���m���W���^
+�*VQ�H*���T�zl�����R�Q'��nE�(�ϩv���>������<�	y��Q���r��pta1�?/K��j/d�]��S����YzF���ě�ra&҅�5����8G
�׮���خ��>k|�;,�u�u3Smm��)�:C��7�fX��Eg�.�4`r�<-9�~�L0�my�z&����K�M	�n��&�#��G�Zp[.`�ڌ��|��2����_�Ug�/:}/d20� �i�P�M��"�$O��(~��
�~|/,$���"l����6Jm���!�X�Y��^ ����]\]��������{�	[卍���*�~�~�2�u�J�ejZ� 6���JPȲ�s�r�]*�3+�J=�q�ڎ�0�K�Yuh'~�F^��}Fɪ8^)
^��o�a�^U��;|`��6�������V����:|;F�v�
�V���z��a�i��P�v���fc�*eea�'�@�ח���O�?�pO�~v/@���K�;~T9	{~^��NLL��Ɩj)���j�h�%=��U��𐰅�9��b�g{��Y�:D2��
9�~a��k	��p�X���g��+��oVɴ�=0��qP.E�ĥ�l�%v+��_Y����������j�=��;����6|������"
��\��o߮�>ZDJ�Vb)���p\)>`����d�r���CӢ������]�t������s��y1�'����Os�ӵ�m%F�!�}⯿2�6a�up���Q�:�Ϊ:M�f�iI�d;��lX%%�-ۄ�F�(��?��{�/J����b$A��Wb��@��E�fHx���eѫ��Z���U��B�ߓXo�e���V,)�d���q�G�����2�fdʚ�"R�HǶ*��x"�%N3*���>  A����}R2�0��~��Ù��s�r񻘬�N��2z5�t�ׄ�'i����N�Ҡ�SWS�>@��φ�_�5�	{"��E��b"�i|�Mu�`�C|����s�W��O�j�	�q��ƭ�ǀ��#�w�)�r�F���)���-���k�X����Ё\�O .&;�]a�^��3f�#x/�7.�<��0x��e���2Z�х��b��.�Q�K���XWOT�9]4�JI�����U�$u�#n`���w`j���y�vx5+��ߴ���(Q�"Rc��ܐ���Ί�=�\z�&�J���6K� �f���1�斣<��W���;�A	�>�p���*qCr��IP�6c�u�fլ����ũP=(��я�{�7�QQdȌ�Tcܕ}��~���85���Fأ����	�f=���$�H�-������n�Z��!�C�����{�|QO]����/�H�����ϾT�_d���-	�=���q@>r��m2�e�Ѹ>�JSx�mKES|'�HM>������)����g���`��-f���:tD�_lCq����1�эzP�@��gkgl#������
ߪ�/���b0�uj�����H�C᫸+Z���o: iJ9���HʓjF��DR���Oڻ��hC�\U�g��$��s�H+�\+��j�I�[���>�]8t�]��_2n��X���,:��-Y,�_�r���1�C���r��{G/+�u�p���O$7�����&%r���;��&�~��/E�\E�F���y��Y�t������lve�z��k��"^�zT�5_��N�xXW�ib��]�H1p���|�s`�O��1�-�Xxs���8܂�Ȍ��O�Zƍ��5�J:"\���ߤMW�.H1Wq*�cp$eV�U�+Eè�T�os��h����eq����O�fm����s��M�2��������d҅u�gjs�T���t���{�����m2�J[�	9*+�s#��F�,���b<L��CQvC�J�k E��le���۠�m��T�<��:ܨڶ�g�a�ߣ����< ���L���D�}z���������#6�S+[ނ�� ��Z��Na�9�����vp�\*[]L�A�6�BD�^���Qўch1��t}����\&���5a�od�9�G�'&T��Î<G�e�@_��&*B��n�
s�z�.��n~�Ӓ?�1F�q����-p74�n���:3�mz�#��[g�?h�b��\�$l�*q����¹�����ء&A��$�iE)u�����k�7Nῆ{�Eu*sf���F�iO!<Dd\�Y�$��P��n!d�u�WkI+rtl�㠄���������Ϳ�39���c��=�þ��\��	�l��]x=���-ʑ��
W�,;��Y|zRx�sy�;6tug,�p����k��~rT�>L�i�� G}��S2��3�C�Z�}��*B^o�糮3�>��/1�x�c��c�C=����$�� >rJ���|��B�y��ؓe���6��6��D�?{>�<��`I�ٙ8?%˟��ė�/rT�i�r�BG����*�q��2N��;[�a�߈V����̓�k+��1Qy��_�	�ȥ# �räʖ$+�2"{�7�bE�*�����k<��f~_�8
;E��v��5�^.H��t&P�i��\�Ou��ؓޔ����Y��lz˺��a��`c���.,��SK{c!R(��뒸.m�����D����s;���I�$2��e�Ӡ�úӘ��V�m�#.Ц�7`� �E�����>"�a�pP��#BPb!	�:}~��"�r4��*�ĉ To�ՙ�h�hrD`��MJ!'����5a�p9����sKTX���>;�ep�FϮ�1mt»#ۊ��5�5�25���m�Q�#W�b ����lo�?�ܶW@5�� �O�٩���|o_�&��^T�2���dU&��r��.|�%<h9��'͂��IV��f���z`�`9��&�l�ÝꙌ�f��&���i#�Ĥ�횓3�v�}&P��u@7����"��(��.����O`n�N�[�u���Į����0�1���!-.oN�D�Iw�s����gҊ7'}h�^�=�V&�F�[�u�~�_�|��@e-3�0�(x��]ce����P9w><����8�Y�����nt�����,b+�Q�8OgeB��������3��aZ+��=C�R�zۻ���b�>A$��c����#�O-�ñ�p�\S��u̅4o	�~mִџ���G%o��'hC��)�p���`X{H@9�k�D��������!�/��[9��(���Ї�z��`޽ۣN*!�磯���0�i^��#��p�(���W�_�U�}�l����u7�+�0����wu �7Y:��C�[' nA��pWݱ�2rpڗdr�o��!��6e#  �Z��z/��{��)�{�j��p�'���~�;�ၮ��;����b7�D����1��=ٞ(�P9�P#�\���J���5��_P�q��ν2%�1��+Po������0�x�	m��z�I*=
����3��7�y�I�|Q����X���ν6�D��)�uI-B�A�fu9s;GnIs�C':X'��@G�z#�E�ŻQ9f�j��&-#��LR�8�y
��2�j��I��#��4% T�nG'az�O}~�@�����GO���-�`��3Vv�磗��'��[��bʑ,e�Q[�A�3V�Nv���}���(�!�_	KоF�q@p��ȼ�S��m�%2LeK�������9������s�m�����M�|��(p�NG9~�[�dI�����4���3���#G@x��1����������4޵���C]�x����Ɠ��!Q!����$J$?VB�]��'D�j��;~'�xa2܇���бpQ:E�#��J;�����ȼuʙ	2��~Z���ݓ��̱��5��cIp�PNп��v29��o;���p�_l;(�LC�b���#� H�Z�ke�=Ѩ� �~ӿ3i��a�p�1�sӭg���=4�O���e�~:��ީE�������W�rX�G��|/�,gi��G^�[���H�3u;4���>�q���	�	�J��|���j�:��e
Yawm_&6�ǂ��u�����kD׹��G�\���`��eF#۲���J1��FG��/��v��.v�	��z��H�_�b��_���T~X��e�����*��&� ��m��[Q�4RG=�ܾ^?/P�l*p^���A�v�J�~�߅��^+|��[h?^'$�SJG(*3�k0�K��_�������󌽆b���XU�`�VL��%"����G�
`s���f�>.,(���sO���҄$ �`�b���S3�Yn!t{�|��dUs7_Ʒ]��Z�R)�r�np6f�&���*�&"31��f� �����#�\C���R�� t�@L[k�:Z�l���:����fΘ�	=O�Xr/�&�vE�����/nG(������
����e�����9�æ�٥���e_9��Kpŷ����w\�*t��_��"��e�[��N�1���h�//�.�O3�!���=�݇x.���儜L�H����[v���.�a�y�����G�'c �j�3G�t���r®7�3R]�P+�m�ܰ�����8�@��Zt���i��o=,O8��҆mZI��Uo����$�����:��|�\.;߀�(�@-��"����Կ�Л���Ϧ��Q:����ޏ�P�C����m�5�I�`ۑy���`հ���w5�Z~ƍBӇ�<j����]	G�Z�cD e���3�eb��=(���F��zj�"���w�&pI
�J-���[�q6oi"��U�`�i��ӱՇ��FB�K���Zܜs�Iћsc���U�`��'D H	�kΎ�$�i��#�$��B�4��=OT�
$��a,���i_���JVxh���'�������=�����IT��\57N��
D@��=�#�Q�UU�v׎�?V�.33�i}��gC�������n��q�?��a�qj���I��#�b�ښ�X�[UT�A�Xd���`����-�~��O��$�Zb|��9(\�p���s�16�����4�{X�g�я����D�%pe��,���w�;�K��H뢁?PBNB�Ph��y�+�޲Ӄ`�-�B��r���M�+c�Sr��N3���EK�!>�}}"�l q �+N�sJ_O釳��Q×��
^�DP���p+.���)k�HHO��!j?�IvUC�K8�t߿
�v�M����#:�}	�?�@q�3��9�[����֙@�!�U�r~>Ȓ%��'��G��FK��出�:�E��g�a�.�m�p(B���z3�U\ѹ*g�0ɛ crT��׈���G�$8O^���T���>9	��pa9�j�<��'�`s\�|���)�Nߓ/GO)e��L)����1A�h�h�S��fbv��5���0'|��ݔ�"U?s5�=L����}r�a�}A���S�v�H{F�Q��ř��O�"$�,[Sx���������]��JK�k����d9�p�h(��fn��A��Ĭ��0��⢜��-f��d]ϒъ�&��@�s� �����U��
�p"
8Ucg$��@�j<�	�&�Ɔwn���Fjp�5ֺ��s*҂�@/�_˃@̏�Ӷ���	���5��8�?w��|�z��.-�:�d7<��Mϙ������C�F��(��ef"��	)�$����e�Bh:�?��c�l�B[F&�
	�mW�2Q�|��[_>��-m�]�)Z�8W��z����yu_�84~:�d��T�� {������4Z�%@�D��x���>P_����J��D�V��c��3�@�W�n�S~T���6	�o�|`�x�/�0�GRo�ձH�q��?\�"n1䝜�_��g�9�;���@�I��� h.C�3�|�!b����&�������m�$B����>k-@��V��n)l�u�����^'*$Z���Z����a*-j�޶�([gM�3-	R ��bB�L�I�lB-<�m_0A~�.�P��!�(���~�gfˏ�7��n��j��?��Nd�'�*&��A'���DpC2���,�/s�a�v<a/�WmNhϗf�*C�0F;���O�`"?��9s��.%)Y�yX��x�5�r�����!A껻�����Lo�j���(	 ��v-�����dL�F�^�rjO}�;&����j{3�z������Qh�=i��*���f|@��$q�]�/�L:^��F�k��i��=���>���U�P�)>���9vi�>���Tbz���R/�`s�Oq0#cnۣ�!鿇�6��OWk�휂C9��*���Rw ��7��6g]Ź�9P*���C��$�_�T����ɒP��ż=��wͷfB��y�����!�/��yd�6�� G8� H�:��lM�~���=a.�4��@C��_�m���N/;��%�w����aa�ax��������q���0�)�"
_�g��G*�&9-8:�]%��-��A��?��n�=����0�8��S� &V��]�TZ8�la�=}���}���X|�$ՑK>��6v���_���3��]V�ҝ�n���F@�7o��;}΃�]��M�-T����?/����T����n�Yo%Z.X�O����Z2gcj���i�A�q;T �J��� ���Z�C�&<ƼkTG�K>��g�>%mO�ʏ���0Ki�2_�^�2t2� D�a&r���ڞ�R���Gf�s�4�H}c��"�6�=ˡ�Bc�j�L�� ��V���3���^���_?����!/O�`��M��,+A�PU���2����ȏK�Y��~�[�/��sU�o�U���K@6k9̟$G���9Z�ԓN�j���.���ٺdDwW�xS�@:�д̍0m�4��/������\�|P�k�C�,����uo�呿�P"-P2��"����$1��G�倦;���*�iH�pzjF �3W���3���7Y�#K������i�lOЀ@Fd������|��]����v/VC)6hY���I<57������mqㄞ({9��tPn���u�������V@��r���=uG2e�_�u ���=��E�*�K���!V���ݽ���]j��^|DC���\����O��+.��t�"���u�?�����mxK�v��!卂�Hh���C�����_K����7�=6^�ݿSU;��� |6�\k�;�Qfx�_Տ*��z��;���Jh�<'�
G��ٕ	.�Klβ\�c����iw���Rr9�ٓ��1��lA�B�6�b��+S�j�B�eS^��/|�X>τ�>�9��+��5��y���l��$J�էy�\Ϩ�9%�
�n�gA������>-�7(��Y�b���W6x�+|��O.J���
�j#^���"��o�L��f0����|��q�"��vK�F4\ѻm�م�ﭤ���:�g*���*�&LpM�M��t������Q+AҲ8�%��lm��Z!��V�b���>����*��&/���T�'���'y�>�ܩ����gg܍rp�W�M��f��hh*�8O)��]�:n'bg��WٲJ5&��±�)s�N��oy���X�p�
E={��6��kȖt������O�F�R��M�hm�_O.�
8��{˦���Y�OG�d�F�vnxa��˧���/����8��={DP�u�eC	�Z�������i��!%��ϪG�(n_T!�V߽H�i���*з�zs�[P6G*T����HH����1`c,F�k�a�F<���!r�]���ӆ=���[����!���@�����h�:p� ��=��3=4ؒ�ɯ���R^��=�}�]���?�|�{矘��|fa��#���cÌV��`�� ��|,PT>���y���r�/�fɲ���0�"v@LH����Q��/�厢ðS����l�K���B���r�� �D�}:�v�a�r�v�L*؅�J�����:m�������h�2p8��p�Ds$˕=�ƌ�!\w�z]d|Ѵ���Y�5��i!!	�e/L���:��g(,E�y뜬�ւM��8`݊��e��3��G��	5�3S��m��礐����-Q��H^h0}�L�_��cC�H�U!(�Pr$��K~���]6��Rn��-2u&\~�$ܾxثU?-�]/؃c�OK���^`4� <�K��(LP�V��;�� �~�ރy����Q�.�N�C0Иh~�����D(�u�Ҍ�U���:�$�}���D��~��Sh����J:ˢX��(���-4s]"K��A�⎃�����m�����b������>����Jr�P;V�$JQnA��wjo�@��tGBWiCM���e΍" 1����i9�Ƥ.����od4_�P���&������>�'De�Q/Կ�8��d�� <�Huc�n0hEFu^Yh�c����!��Vzbp~��1���ُC8O��Ƿd�MV�f����뻻w�k��kȏ��@ �;/ ��lY�_4�$K�I��V>>�k��1�\��ɟGv��q�y���fO�Iq��Kub�l+e��C�P�,��\Cj�˭N��K�����,z���m0�� P8���M�c��ٙ�C��⺡���,6���E�Z�	�z�3�N��3�oU��X��f��v 5��t0��O�a=����EJ�ƨ�[js}��E�ٌ��8b����p���)"��It��L���*ɭT��yw��ن�1_VQ�el�+#���.n�6��L�E�y���H�^���2��#de��CѡRI9HfB��Ԁ���į��E�{Q���P�b_j'�t�y�7z9���$o{�n�e�	��V�rO�I�ݓ5�SůS@j
?u�@���{4�5S�#�-�W	�ک���mIHhU���}C�s o��z�ߍtF���y2�:��/�D��f-�c+�A�m���{�g��H�~�m'/��_���L�����9���JH�R��y�}���5�~ ����(�>ʖ�وݷ1%���� �y���" �1 c��?xY\���&�mk�c�l��2��0��1��*Ztt`�*K�E��[�O64Ft�#{� ÿ,1�5��;T�ǟA���	�j[D��F୭�gZ�^m<(���6��OY�#��&~�z<3��B����+���lWIp��p��CR�ukX���HC�L@F������8���F�n��.ش�!K��kļ��*>!DUW8Z���of���̹;�����(�`�
O��>�Ͻ�WhP������F�<tJ,e�龰]=����$E
L� �����U��aJ��㉖mMS?�o�ً��-�vn��U:߾W�	�.��:QpHk�̘+��#�׸�`=ق�.�L�P���<p2{��Y�S����QlL[�B5螎��t��X�M�ٵ�tѣ��p�S=�i�����?��f��<�Suo��"$7psX����H(��L(�&_k�C�[݊��q�k�Z"��n���_El�\�����-R��~�Z_�ңs���5.�rYL���i���5���o%*����]CfRt`�m�^�\�ㅟ�<���n�R	}ڭxߝ���5����?e
�S����"�%��I���a�d��ѣ�Ͳ�����*��Y�'��/�HJZ$���S��(�F�s��?{K{��
<շ���x��x)�5��һN��E��ٿc�r�=������tY�����ڬd�K���UZ��٨3ӕ5"US���cC��b��U�j����7�*C��_W�4D�￧B��d��6��O�=+�ƶ�.�Yy��H�	)��q[;�>&c��66Iy�w�ꋬ+v`�kj��L��&r��VX�U"/���m�ʜ�9��I��
�U�:2��	+��*G��Lo�a�5��U� !�L�w�(����k/�� "*$a5��z���C��?=m�7����S���H0�����iS
�2\��F$>:��	iU��a�6��ѩg�5Q�p�d�����"����u!���
�N�-O���7L�kS��`hf��}���^�QآNF�j���)/����iw��П�y>�9[)0 � ���?������)�%e
����84����x�a��~���y�CH�8���a�����!�c�߿taD�=�Z��qB��sC�
F����d��E~��?�����|�[���A�{s<YJ�F��v����5�_���D>��-�'@�j��m�����	����?�a���q�!t�<�����I��Wm��,�`����͓����fR�Zz��f�Kt�ɣ���픪6�=��A�b���7�>�o{o ~�����$�t�$�y\D^IC���-3(�\g��m�i[�N�0���2��m .��y�����́�|ڣ8څ�y�ZTIY���`	者��`c,�&,[�#�{줡Η����k?�B4Qh$��"D6ꃩ����|�o�@��V��h�:�y���uO�#��q��RS�$lf�I���㞔�R�YT�����X�y����u�fpy���0��0�$��=�2�>��W
�z�F���*�֍t���&X�,q�Ϛy��	/re�(E������U��6ݭS���╅��W�>����YTgnh~�!]��GR����˹Ļ��vv��Ҝ�����Ø��p/��2��-P"�'^�ί�	f%�6
A�A�<�`Vb��ҀB������,�I���b�����^���U�(��C��8����o�e8��4��2un�ˊpKa��.�5��h���B
���O��\�QL�v�o��Kp��I�M7?HU}b
�_?a.f�u/|�w�b��xr��E��Ժ��EX`Њ����d���~V�(�_[pzKݠ�)��T�`�E��-nO�Y�咦ؖ\�'T�+�1�9����,9!��b����	�C��	R�j~%6��>=g�@KBW j'���P�k�Ï�\%d��ǹuOjP^d�qXM�ڹ~/�b�lY�&�c��sDs�%/������i- �Ì�6�c��G���M�I��Ւ>ߝ|:ٺL�d��Kn���t�"�<{��b�镐��;m�5�z�Ny��iN�iBrS���Qwr7�oT۸VͰ3��:��TO���X!���nݵ�t���F?�9t�蚤��I���4���	�:�Sba�����������)/	���lZ�����e�Ƙ�Y�2�0��R�JqD)�i�;m�=��f���2)A�W�v�����һg�T����M�ͧ�nd`�ϱ�	S\q��IG��I�x��j�Z���z�e��rf��)�-������0k�-������[;3C�������=���I^q����^�lҵ� �!����i2��(dў������4 (H�_a �v��5:BY��e�BX�Z�ZS4��D<)�cx�Vz�x�T��}3m�t狤��]wHj��[i��m����L����6����'�͸��"-Vc��c��(���, �Y�,��p޾4u�v�@	**��i5N=ywK<>�����q����E�hm�c)�e&�����̇)[ˆ(�iZY*��,��)QX�l���Y�O?0�p��	rݕ�{Dx�^�%��G%�?��{����=�����}�_����YXNy��j�A�z�媶�PK   �i;Y=���C; �; /   images/21a1dd99-e68d-47c5-b9b6-5144ca492781.png\zePm�$~��.w� wn	�Np���������C���������nWM]U�c��{z��&\IA
� Y,�U �ϙ��=��=X�	���?�{��+�秴��7���.�,"uf���_9s�-��d���M'�!�������ǽ!���!u^��$@�������������ڹoSNh1Zm�MFqrl�~�v���U�e�Z"�N%5���WmQ���hۡi��[i�.����Y`e���K;��0��i�9��)`w+��nb�����mL���Ǿ��ӥ�pf��	�7h7���(�V$���FH�=+q&d$��ؑ*�uP��w6��Tّ��Έ����]�&�㺝L����ע���n�&�����Y~6�&P퀠�?���?"���P
�x0g��狅���u`��M��2��^M�;���_a��.�����9��D�-�D`����7�Ϡ�~�P��F�;�<1e�٠�e4@uļ�	%�8�"���f�r�	zY1�
���M��)&��@�x����҈��k��*�P}�������)�.�M�~����6�3�4����C{+��Chl��l�.*Ǿ�0�19Q�y5Rҳ��R��0���W*���]+�k;�(`O�����k��X�I>
��]�*���{[e�6�Ü�Z9��I�̬_x���o��N������F1�k\����|��&o�M-D�9��/#m���cū�m�B�����UȩY�L�� ��iL����lZ���� �V�`���~���v���������J+5D�7�;]�ׯ����>�ʞ��Z��w�ɓCiCF���N�/���tC_�=r?Gj ��� ��?GQ:&R�ݗv㞡;x;+/a���r~��?F��r=��{^��;}���3����s�ݝC���q�(BS��d|)b|��.95��]]�d���������>ܱu�& *jE}zP�W��E�G�LkS��b����6έ��ف{$���Ϻ��}d�U���)H��P��#0����⠼Lt��EfJ�7�q��9h<���p�������}9V������ȌS2a~�Oh�>���`�#�늋C\T�v���T���v���#H.�9�����(9g�P
��4y�a\^��>���VV��_�[6�#Ό��+��l��U�J�A�w�>x��'���l�sk_o��Z�E j"��s{f�@Xt�e���
����bt}�`Q*�Mב@�܎}�{�!#���?�����\Ӱ����I�����[F::+�ɱ;��U�I�']���K���íe꽖�՝ui"~��z���q���:��/6I�X�Nq��z���.hB�픰Sfg��b%eR�x�L�N:{>�R;.^&d_���-��Q�q��K)�2�R���Ed"��EM�1]��@�L\�j�zZ�#��n�*���E�q�2
�Tm`Ӗ�g �@?��L��h����K��l>�ڷ��GsԜ��v� � ~���hT���p�7�rX��1'҃���\]p].d�߹�7�7?�J�P��5>�Iwf4~�P��U����k�.}}n>]Ϸ~ڗù)��O\ox`8�Υii��,��6����
�z�%/����|Q������Ԟ����-n�g�Q�Q���&S�A�F�Jp@�ܼ��Չ�.��`��3"B�Ӝ�� ˌ��o3���_���T͔(��� ��D��j��+Z�S�R��TB�I#J�B�'v�Ɨ�@��2|V�0��d�X��i�P���~ ���/�z����;d��"�yu�Bo�\��U����#��bNϰL`���Rg!}7QM
 ��)�t�Gc�Q`A�Ў��ޢ
tA}���x��Ή�3bVصR�RF�S�>2�lx��z\O7us?K�\��F]�~��{R�+0 �P�i�mҜ����AR+�x%Q��b
���d&��6!:� �|%?#4Qԏ%��4M��%o�^V1)�NT烦�����W�Ϟ����c�~�JC���/����Ty�����|�N=��Fj\�����\�����n�BC�[c��IP�q��V��=Ei�]J���=��撖g�޴S߳�c~�[�Wg�a�4=Dz�:`�g�#��_�,��4'�Ɩ��ݢB|�`V��P��.7!��z�?�Gz�#��j��.Ԯ�QQ���X*�z�G�4�ov]�O�B���Se2��������`��i�t[,�F�K�G����OU�cPn9i��!~���7"�ѫy*&��}���F�0Տ��![X;�8�c�<О�d(���Ӭ%+��'�Y���plŻ.���0\���QXq+���@�`v0�N�`X�]��\��I.mj��Js�wB�zQ�h��䑦;�;f�ybo�l�����&=�O����k��xK����",��1��{@�._8T�f;���L9ѝS{]e���/V���������z�$OU�(:jb�;���#���V��nR��pD� z{>�9��f��πtԂ%J�,l:U_&��o�1C��:N��~���jPv�*&#���=��Px)g�0I�b����:�Y����:��`�r�p��p�l�q�zg ��u�߳�;��͑�!ݢ�zM8j��8�'Ĵ#_�7�)��f��"!H^c���2ҵ1� ���D��}߁�y�^V?T���<l��Cd)�e��[c:v<l�!��xP8�u���t�z�O�J���c�Fc�D��;��i��h�N[���p�[�e+�p*m��/�%��ٍ� ��uwď�*qN�8��AV��_��A[�+���׫������$k1v���pҥ1��U�z+��(�Z���7��myP�R�}��pV����,�t\<�4�; �4����ȩ�	���r��;���lV���_�HX��%z]تf��u���҂?�����4ep�x.�-De�Գ��ό,l�������D���(�e�U�TF%��/h� )��C M�A<-����l��������[�E�Պc%��	�UO^�^�m5>�|3 ��ϋ]8����특s�fG�Dc�v�C���@L���{�G�۝y�KD�7i�|]�Q�V���vu�B7�Px��₪g`o���>�93,�5N�6�������soW����l��s�/خ
Һ<Aq��n䐲��!�$��zk�H>��еNӐ�?�L�����D`�`;1�,���,���V� H�)�����:$m�2����Q���~=�cH���k@�L �Q�f���E������dޫi�� ���Ykt���H����,�|˷b��+ݘ����Ik_�������L����\ˉA/6ꍘ�ެ������IQhӥLHg�}2�j�S��ҬLɯ����Sl�y��5��&ԅ"u�(3Q��@�.���ۺ��Q:�3,��"�'�ȨU���[��iZ��D�`K�3S�Q�X
��:��g��n��$�ޭ�u滸�oP���'O&��&6v	/}���8���9)RŖ�
(ڲ��@@A���P,?6+��H؇뢲g����9�P�s��;�v:�]x����C=]�	��a�B�pFL�[$���9`{���=
@=
���̔�QNnb�7�g��[,��bCſ&*���<�N���)�f�,��~u��0��g�Y/�ITm$����<�w�Yw1�=#g��Ꮍ�h��f�a��W�*��,%?v��w�aϐ�ҸL�{
<4i��yV�!�bb\��ܘ��Vwu�₈�l���k���yܯ�R��-[yIǆ��rA#�����N|��@;��t�w�_�I�����AL(v��bQ��ݍ����v���{^0P��9GW$�ހC�#�֋�S�#�ev^�,�o+g8, h�#�9dB�~UE~���oy�O�;ե`��/��3|�ݞ�v���(L )��*�..��Z�g��6��͐УV�;	P���e��b��J��ԩū�t�
�g�ΞlJ���d�EB\����I�:O����ZX��$��>Nka���{�SGD$~�Ut	��C��l8M���(lV�[Z�!D�Nk�V���h#M�@iik�eN&@#�99��y(� ʚM�)��v�[�P��([0�����27B2�r���j8���4�؝�m�+�X�鄇ow�a�Z��v�P�'�؏�㓏O�g��Gr�վ�auvٵ�5tX&_i4��X�3nS���i�ﵚ�_�~��e3.� F�J�l'W���ڛrͧ[R���O��vc�ܪ�Ml��:K�k�`�*���E���䎪zZ��:"ń�o6����(b��emb������������9��9ŀ!D�I��;��<^Ǭ:ɬV�|T\x�@;O��D(F�[F�a�渏����'��J~J���u,9��o����o��g�+�0+�t6N��I�%�iM{G���an��Cr��.��ew`�j��9���PT�/�g�-�</J�@EMрyʗ�JU����M��u��	��zT?p��� �t�s�:�����޷��x�❂#$�7,`T�
MW�@)�ݸ��L�]�����o��0y��� j|Q�)\���g/��B�g�D���oW�͓,!Lm�D�T��q��N|�Ru���xY�ћ�U�E�t��;�����&J�H�A��/a޻^�6����@^�+�&w��n� �ԕ��Ġ^����ڦ3��GF��#m6!X����)�·�����2q��\y��V����;��l��:x��Q!�j&���u�|�mZ,L�Ό���%U���mAY�ɯ W��&K�\�쫣��i�WF��n䌌L�#wk��p���7���B����1��H��8k%�=�՞Re���V���{_��Ǜ�\�.�Z��J�O-t��F�rH�!�M��.�1P��o�8I��b3I�,�I����d�Ez�.�֣m��b�(��أVk0�����凅�Ց�[��|�Bô ��9g�i5�?�]~(V�`p�D��yoj�uy4Y!,/�%�c�os�ݛ�+_���+c�/bo/z�-�(���ߋ��L��:�<���l�Tп=���՛�	��u�Ñ�����ڔ=��;�21�Gֈ����n�Glɥ~B�E/�Ŗ�[hͶ�ե�� �9��h�q�ٸx�n��,7��\��u�w�ikO�Ǿ�*�e����.�f��[/?9a�Ɗ�����h�����N(��ni��1�ԭ���a�'�`.����8����c�6��ۮ���T�)�[��D֍��\S���abe��&��T14���D����h|8�����R�ae�*z��|�Ľ�G�t8[�;�~��~��8��P%�o��M1�?��3�	U]Ǖ��@F"n>����t�2�*���H����k���V�zlw����6��̭փӗ8m����>Fn�@47��v�߆��s-kĔ�jN̖��-T�����d�v� �}���}�Kֺ��-����Ӊ��a��_��k��l����n0\�0zTǼַX��K���L^��� �O����Ga��}1)*�GЮ��%$4������ꒊ�����D)YU&����ѵX��Ctt�]�Ճ�< f�d&��<N`���!~�܋�����n(�����\|^�S?�{���F2����O��������y�Q�!!�7��Y�N�G��(��{N'j<�+D�h�AN��O�iW�G��{�X�v6�����8ͺ��S'Q�{��s�W	�K�� -���2��*��<W޲�Wc�"���ti5�]7�%���d����;}��0T���\4.9��ieC���u�s��w��=�i�lZ�A���{4|8[}C�������5��"y�9����Uc�M�P��M9�R��};б�j�YR�l*�DO���6��"�r׀dRb)�7��j�-��Q�����Į��#V]"S@q�t(�� y���%�^=^I�bf��v�.�U�6 `�@�ɏc�Z��s՚O��f�p�r���&��:1h�:n&H�)�K(�]��Qu���G�w�#��7z����	5;�@*C�"���
={�"i���Ó
c�����SV5��V���d$���$	�?�+������S�1p��,D�#�p\Ŝ����i�D�B�H�_��9d�Q��7�֯~	z��ݍ��J����<�)�����m	1e|M?�ۢ�`���#r~��OY
�ht ֲ�r���#1 �<��0K���Ni9��'h�C#A��DLh�I޹�c�hB�
}�dy���GxTO/T"�t�X����a�����X4��~>����䕦dT�Ed|�|�y�V��z���l�cQ�r���x쁀oATHGo���m$|�Fu9��RLX�Y5�R|��<���vD�g-DtxF4��A �<�>����l�R����;c��hc|�y[�5"c6��o�����tc2U��9�3�ј��	J����������ۗxy�oh�LB��C�A
I�HR>�f+��;�/��!A�?�#����X����(��)���Ϳl�OO8굯*�0��=�g�1f/[`�=@A� �.|���|+E��� ��wϩ�81Q��g����H~�����~P:�#��'8�Q��i�����p�ݽ`Zkx�6�t�	���C�l���lS���q��[��簓s�Ȝ�����\W��C����s�[���}�-r2��"H&E���|� �߃d�U%�</_�]�ؾ���r��0��G��:��NrfL��2o@�k�G�s���ր��s�,E�X��:F~@C*#��p�A\V;��+��^�f��u�6��z�gtj��dD�,~��Pˊ#���r�3���i[�0����Ck�C�6�~B��c����e�B�2���ߟ����*�M���
>N$YTև����\��x�TZ,QSX�!�t��b K��T��?����~�w>�
GR& �W�+�=�{x����A�'��Z���!r�����+���Q9� �ڴ�t����ii6�wd�.<�T*0���� �SԐ�e�޲�d���A��8���GsN�Q�Gq�ގ����p���Kt�P�n���%�xSF�*�Tfv�W�a��F>�ͺ���x����w�]s�G��{T���8�ď>K��S���ݹ�i畴,���#��G�}��	�¬˟O�D
�URWi�7g{�Ӻ� �u�D޸j��g�Gd����Wҫ�5Mx�tI)P{-J�Y՞�=�^a�����b�6$9W���:<j��Y���>ѱ�n/5z��6V��l������\��Dq �m�yc*�����Y.f9���-<�$m�-5I�ӁxҰ��)�":XN�C2��B,�g�����B�&*�\������62Gy#���Eɶ�(��?R6`�
y=ٯ>")w�q��AѸƘ�vT�6�j|��&��\���v��U��g0���l�O��ņ�ߙ��fsՀp�|�Ģ>^4XEe�ho{(��[�LT����H�=^���
�hcNi3�%��wU&�x*[�-Ƽhuy�Iߩ�i(n���~���2�5O��|�5
*��&H6���Y3E������t2a�i����^�T�GL�s��Z���w���|�I��C��uM����ے��h�
�C����(D��dS0/wl���?�KS8�`a����_*u�R�	����j�;��_b�n'��Ź��S�t�IO�P�Y�QM���/oH����E�:��>:���
��B�b�w��ZI[|�F^?�������"їjg����3���p�n�r$D��2K:���)�� ��޸��>��
��=��Ƅ�'*�?&����p5���\�� ���6����3D����bA����6��j�˙$�9t6�΄�`^�1�[ӿY~O�Xq�x���z��L#� Ć��X����K�f��ET����r1����~Nw~�Yjqc�yӽq�Ohk
w��;�%:��	����@��������X� ��%�}4b��,,u�m�!����py����~��ؑ\.����~��4����꒶�`ms�"JZ]���7�F7���T�w���&�l��ke:Y���*db����2yLt������1쮚�/�ٽ�������;��k�/�0k���)P�m�li�'��F}�YG�aɠ��2�u�B"�~�ylMǱN�e ��pz�ܥ�n*� B��z9��m+5{Q��1�	2d�K�]ϫ��!����-�m&%�����^٦5���S�	f�o@��?pF[5�
�y)G�æ�"����J����ſ����vR�pE�up��\	y״v_N�5��Gqѕ������~G�s��DF�9�n�"�|�l ������A���֜�l�R�of7��#_zZ��������3>=CU���_�_���Z����69�==���_��2AB�R�!����G^���G��M��
�N3�L��D��=??7`��+��bS���/�������;z5K����y9�.�,s�D{�njCX�lTȈˉΙ���nw��̍���v2��?ڡϒ�
� �����̬��r��p" y�q(��Ukx�x�?�I+�!��Bj�)9+n�_Ff7y�@��$�DA���a�?����g���_��Ŀ��D:��?�Q|��í���DS~9�FS���$�޶8���Y��US.��w�D�Ε&�l��%��n�X�7DrT2���O_��hs��5�QcО��vI�%���2��x�Q�V���R����;��T�����]/���
�M&.���zޣ[t&�w�V�V$3��z䙐�������"���.�J=_g';J.�>72�4>&-N�����Fl�֭ҙX
z���[���^�.��o�6+y� ���F`R�+���Ej_'8�Ot,���{���������9��^��E�k��q��[h`|�,l�Y�����.��{!.�_0���_�� ���qL�J��|��~�m��CӴ��������I��p��|�nRĹ�����V�A�5������܃6�F���q�_�h�]�����\-�3{��`Ik�;�7�~�a���8��$��|t�SV6E/������Z��%o�K�3�(�� B�a��r��Tj��?��Wa,s@����v�����%ޣ���ώ�D��fT�i:�q�4l�����LjO��噢S$�aT^��Q�LTeR����Cf�pT�>�E
�f]�ld��N���l���Ė���'�I�v)�`��a>�Gǉ��,��-�m)ebh%��֒X�X�^�g��ܟ��;��i�#�#_�4�V�D�H_&�Q�+O4��:c���9�P�ߡ��$���b�OcI4,*2���L'%�n���^���v��/ĵ����Hz�ˮ�h6��Kj�c�k�d���y�����Kr�$+�ˀ�F�%������s�'���V~jN(�)V��-�W�Z��Ȭ֨&6�k77�~�ʗ�Q)&��۱G�;�OWB�#u�Z]5	4�_n���:��jw_��)��ˌ��Ұh:���=���pLW�^YK����~[lq�fE�74��i�1���:�3��&t@��\�?j� �(_t�3忱"��j�����q奨�"y?񩇷�w-�T&����_��*���1Dk�{OOO�RHg"�D��-=��k�"W1��¶�� nO+�K=�2@V\Q��R��g�_ߤQ�������&�޹�Қn��wo߻Q叜J69��ߋ�)S�R� 
$*�J��]���QIu�:l��}���YĶ!d����B>�
����$�kQY�bJ�L��O��غk�}*��hEa�7)��^������U�Eؗ8$8�S��IS'����&tW��Y�]�F�Q�h_c��d�De�����Z���*mñ*L[t&��p���̊n�Q�+��n~f������Y�;V��r��9#�1޸���s��X�ѕ*���t
���H�HTc�	��%g��(��?�ds�M��<1ٚȀ�/��{R,�Q^��P#�I��������*��S�#�����bC��f&t�1d�����50�;���3dA6�<��wz!-�נ(<`�ݎb�cu?���� �$ѫJ����I�������Xyo���ԯ�	��v9�[aO��=�8��kG��4`}�Z�Q#�!�d����n���H�f�2c@W�uj:��Q�z��F��9UL��&�u`��bւ�Z�Tqח('Md�g�����mV]R\�H�����ٓ��X��<	
��ߔ�E\3��w�L��؆4�]y����J8�N���_g�^�wc��5C=�^�� ����9X�0���|�4�.�d±�*�d�R�'�W��-���7��,�ݱ���l��A�Z��y	���Re7������9 ��].o�?�*��}���u6�[�H($'��U �o?�IS���'���լD�1	5D.�m��j'p�+z`�6 ������zwP���D��\�)gzd���ԛ$i��x�ZAռH%����|�.��%���/:���UO/%g������J�EH��,��SS�݂P�%T#��c��ߩ<�֗�S�L���:���lnl��:���J�VqN��MV�"�Ga	.m�t#�5���御������xR��I7�+��{X)DrVr�d��j��g
T+4��h���n��38nFJ�EN6l�(��ӥ�/m���ƺ�4H�ظP,��|��K3�W��ߩ"�_M�\��sb��i}�30�R���@����&qcÅO�a���Q����O����}YC(X	D�v~���9�(�ؽ���-/�F��������/u�ݓk�;�#6�����I����͌2�u���;��I�*x�ܖh�S�d���<]��o��M���u_�(�K�"���fNà#l���u��6�nhP��!��n�@lJ}Iڼ���X�f_��@\�����¤ 6I���6U�o��l$+ݟO*��Qqn�U@+]�{;b5k�/��Ԧ���'�a:@�/��F�J���yn�\D�M.�l�g��C�g,z��:�i�u9c��D|2F8lv"̬t�HI��I�G�&"<���I��O���3��%>BX��N I�u2V�oG"���/^�:���z	�H2E4 f[+�.�f��]0�vq��Y�a��>w���~����Nm�zy������7~ROb��\Ob���F1�I��?�'�*���"C�8��vtC�#`&��*}2\�Dݏ�C�m2.���f�ٰP�ʶ�B��1R�r�isi������48ܜ.<�k�w�ң�\���0���$΍2'���mQR�x87T(��Sn�� ������ڿ`h�ϲ=���+��g:ʢ�Y�V9�Q�bAs�]�x+�qi5e�E��gBs��ܥ�v����������$K�\8F����ƃ�k�Np����ˮ>I�Ү�Xw��?D��� ��G4๱X����p�"�S�Z�G~z�ll���!{/�p�n��S$-�n,Sl���E�<+(fV\�����j֕D�UՒ��4y���:
�ZT��=s]�b:U^<�GC����?���dy�\2GP�����I���y��Z��A����mq7���,#O���5�ᨓ��@��̚vD�&_G�Ê�� n�<,$H���T��뭇�����U��ꉜ�3m���O��BΧzEC��&���!O��J�����c��#s3I����2��l�!��u����!y��	�}�}����)�-?񀌛!� 9)����;^ک���@b�B��h)s�N�y�ʨF%}��wG�?�Ժ[�,q��E�j���9��M���R����MTv�|�ޛa+��s���	��pa����c;U`El�b�!h!������%�ziB���͇��b��R�nf��x��ĥ�$j�>X�k��/Y�޲��J &��O�~4d5Rǵ�م�9���o�b٭̵�,͝PL�Wze� ַ�m������c݃�9�dӿ����f�o)�re�����.�Н�Iy��	qqy;��x��M����=.�~2��藡�i��Ir!9	ޢ�����]�_�<�>M'ٯˍK�3@:�}`�(�H�8���~�u�zB�:���pB�2�P�h�3'�|A.�n���|!�f��l̠�|��@�r�y��!�my�6�5r@�ޘ$>ܲT�����Ge�I�X"F�����)�n7��b�2�)��'��}uI���c�[��X�MgF�P#��S�=�ep~�I.xT-�9r(C�kꚆ`X 6�#�;*�b����`?uֽ�aG�Q��6(��q�o��y!� `T��� ���];��Çulk���f�5�'Wڌvѐ��6��`�8�m�1;@���y>�'h��FQ�|O���)G���W���m��֋D�=ᓯ(Ё�,��3��]'$�Tq���q�;�ݓ�~{o5<�k�Ik�1n����kai��]E��32������G:�ݲme؏�?�'���⏆J���?��l]u��]��eN���\c4H�+�^�ج�L)��C?AOu<]�J����cչ?�S4{���b�e��;c�,�U��v�יK.�j��jk�N�Rg4m���Q���Zb�
�*�\�����+f�	B�����K����!�?r(^e����
�����)yY �����-�(���"�N��b��?���(2+�xK���� �.[e3�'v �Bsâ~0��eI�@�3�&�j��Ci���lM�nL8�0�VD�&��I�������F�AAY�΋���c��v�nS8�-�o���[���b���߆��z&o�O��<c�^6���l����Re�=�0ba<�1��r��|ڏ	�,N��^	��q�j��2��
�J7��W��B�_�j��=?377��K�׷��axi�M���t(�2�ǟ�p)?_��w�	�*/����|��0b������E�ꯂ1���oq�o�;p��$�P賩n5��m��sm@�|�^��,L=��૤�"�м�(�%rG9"C��	�H��)�m�)�~�ĉ�50���
��`W��ks}U"P�K��2츾
d Ê*�^����?op��j���<k�;Z�Y�Nщ�g��.C�r�������o�sB%��_0�]T���8��8�w����VmH��@>u�����c4���,�:U�?��� =�b/�o����hq���Wqx
tZ_?B���hl���$�~��K���[��E��bo<�\�ow@:���g�g���}�
�w�	���g9i0�]�%V޵�|���|@��*�5j|v���6��"�Կn\M��*������lC��gΔ����}���%Vk>�r�])�Y �LL������*IHq�?3�մ*ڋ��3��wδ& "Uo��3�rZ����P-8�|3�|u�R�GRŢ��%f��Gn\��S�	:��{��_Za�����s���~�0��VA�Si�T�q�"�F���)8��!�4>��7� `��,�Za��UNݾS��U7F6=Qw	�В��q����)�6�@�5�,�T��m�ȭ/�͗[�b�w�aN�u)G�c'�H�������h�j���#��i�m�j_>�k���Z�`���
�������e���	i@�%���-�����[��WoŴ�>ӯ����Bc���Ж�׸(���ғ ���t��l����8�(�}�D��&#��Z��K�r��Q(R�M̂5�S�p�zמ3�>W ���Ǽ1'ݢ����t���s���"ʜ�(w����0t|| ��p�zn�Mw>�j�Ԍt`v`�3���"-���A�9����)S8?�VwG$n^:�Y�.0RYt�+���z=J	�v�`Q�H�l֓�k>2���l^-�t�'&�E*��E!�y�pBu����͜�xet,ۭ�	���˥@���$H��20��&K6�bqÇ�~�/�|��3�lI`tv�-6X��ǝ�.��N�ɂ�RB�%�2�!an��iL��,
���#�J��h �q�P�й#��(�|��vF" SF���\�%&YR��N\�Z�R��V�j7�R[����P.m��O�d�s�����4���hP]��<�׺�
��4#ޡLj�ntF�8.��F�쌭�@9�60ԉd�'��`��
I&΄O���@��ޝ���K�9G�~���{C����	n&dc�����g��h���egHU��O�_����u����6��Z����">:��W�[�\�O8H�FՒ�������=}R� �z��Ӹ/D�Ɩ��,���E��EZ�G��.?_vw1I�!~�Z���
M�$ �i�S{�#Y��ε�#99�'�w�C�M�AKGH�!�r��($L��^��<�h� �qε~2+6K/�����V��f.���^qgOUB�3^h�1�ǭ��;p�7D���h|�c�OG_��2�4_��@$o{�GD3T��1�<�/#���э��-Ã�L̞�h�Q_B0�p��d$�1��p����.JMQ�/���4=�c&�U�H5J�e�N|�6�Tc+m�x�,�~�ي�p܏�a������Y��>��H�3ήHz���}��0�p|,��@%���5L3��#w����RN��B�<
�V���]Cռ���0�FԔ;>�+��H;��P��B�v�ͧ3v�g�����bO.H��6=��F��Q t�F�<���,1{��^�F�kǂf8������Jb���ۡ�O�A�^;���f)>��
V�~��Z��]��]Z6�wf!DP�Y6�*�E$�r����"��R���>���S��hX�,ʣ$�SsŞ�W���ƾ�zF#?�Ծ��C�X��~�5�z%�d9��M��W����� ͟a�����I{�ZjG����� Q����c���.xrp��t|��(�}���*��\7�*��[�z3��-Se�~aT�r/լ�1�&If������"�����*�3/p��}|&/F!a����Rn�ԓW�8�>�K"�K=����N��i�m��4"�J-��q&��¾c`�>kDA>H-�h��>RFPD�^JV,LK׵��w�Q9^i.c�\�JޖE�})hp9Oiez��-�P�+}m>��\>��2W؝�V��3 �=�~������yE�E<�]�h�.�d�~]Yà(�G��+_�O�ք�_��>z���ejQ���͛=,F��<�͸lv�.�o��;�1g$)�b�����B
��u��\�'�>J�u���X�~��c9~���SǕ�Q�/�z��Q���r �C�,�/��P�ŏ�o�#��{

�}�5T�84�u��]7+s$,��_z1{�������0���H�l%���D���%t���}�]Yޜ���d|\~m�e_����t�g�A������12�`�u��{���,��������OҌU��8��a�u�ݻjH�3����Ǽ2*��dd��:J�;�D3N+�+�ߎ��mҰ�!�����ק&���8�b�;?�������~(I�DA�D�����7`]�R�RH�DM[�t�$�%$���iv�v��=�@����7�Z�4���_
�>8m+�6�0�&HX�,��Z��{�a���S^��[R�f��T��W��-�~�o�������;���P�frLe�h1T�/�י3�]�Zh���Ō���bFMn;������TG�6Q�HDҹ�=� �m[�<�t���͐�5,+�vz��G����Ot,Z*Y��_�$��+T<Y_E��,�~���-����=����kc\�+���^$ b� &h�ZWE>���Dń�RVR�]_��c�+q*�h����h���=�&>7�B&��1u��z�N.�@�Zs�?�@�~5��?�I@��
q�ieS��!�$Vp!��Ԃ��ki���3��`�����WJ+/�8������b�� V9�a���jakk�sb��j������ӡ�b,W����	Y�DkZ
�R��������}�: �m{?�� �4/<��P�S��r�f���,�����>�t&�kMZ�~��S>0U�u��P�ˮ��%O1&CZ�+�M@!��|���/u���o����v��I*�5x��:_�E$t;�.-E34g"q'��I��#R�z����m� ���+�O�P$ʻ	5$PɆJW��p$X9���/ 4@˿%˘�˔�嬡�Ԯ�=l=���Åe	iD�	f��KaѿRQ����_(�R&�*��I� �]H�b}��r?c:6c�i��.!K�,�� M	&�20P�I(8����e�J�/�'�O��>-FvAB����DO�H!��y�Oe��L��s�v��`~DC�)9W� ��X���vW�z}��!�3!�T'"�&E��D�>s!�/�{%=c�I����.+l�J���d�_-j�w�!��1�lKXZH�nPl55��	����n-�KI{���Dt��{�@%א$�Y��m"��P��]\@|�w����L����PDt���*"�2"� s��W�
�	����^��X담M�6Ó�^�=�p��^�^���k���c��x�2��P.���*���h���^4��9�I��>`�~��؇�c�6�Á�>x�����>
G�߅��RR��i�֖�Z$HOش�C5�7vw�����]����3��V[v�T�����3�h����ʕ/��oE��@ǐœ&ZJ�F?q�m)3�A�g�Pª���G������#]gr�0#Ť������H>��h3����ysa�YgCi3�L��5?c�$�r��d�	`(��,�;����?���FrR8�BJs5�۔Cd<!�C7H�|��m�.CV�h��&Lھ�;���(g�)�y�2�E�-k�[H�z{�o����H�����HJ!ݿ{dU|��Tf(�-� �ԁ-�$��u�ݿ^^#��"�r��A���?
�K�M,�Վ�@9Y*�F��(�έ���r+�-�Hq��2���Ǻ֎�kK�Q{A֬Z���-pj��w��p�]{�:V��~��l�t�/����"��r�Ћ���o�U�J�J"��^ ���Ɨׁ��.
�5��[����Qd�z�����>�w���ի^�sbN��������<2n�U����I�[��(+��W�W\z^Uh�p�]�r�(v\�k�=��g���W��t�Z�\"�q�ҷ���߶���o���?�z��av�4�?��(pl}&#���1h{>DJ}>�~K;D`yw�t���ȓ��S���C� �la���My��2�W�Q��Ip�&������᜶a!�����aŋ]��+^�gM���vs����M$��ѐ�@B�hR�R��t^�.%�L�J<ꇰuo/����u���7/��Yv�h�ap�D@�k֬�_���_w	kͅ�2��Vⳗ����� C���;��_̳Z��W��{�qٹ���ӻ����j��!���ŕ��?���3���2%8���5�ɢj{��i-�(���g�F{���ݰ�g�l:��!�.��P���et5	)���倂M�v��u+߸����J��ո��:kV�u+�2j��v<�ݴ, �x��2�_>otL���w����9�hB�#�x���}Wǿ�J�=��~�%�[��:o8Ķ,[�+�Ö%/=��@PE4�B���T�� ~��b��׍�{�&c	O}o�-����U?�A{HT��G�~�wË���I�0"q��jO�E�LD��N�4%16����_���B��?��K"�6՗h=�@�r�R�Y���piU���B�	V"הǞY/��,_���b��ނ�th���K�Ng����w)Ը��8�"-x����A�X�y�)؆s�9���&q �dWd99�45QNDS[''h���8��L�.<+_�/�Y�\p\���C��p��`��
c�}	S��6�iJ�)�z���x�x~-�D�x;#���׀ ���K�>��6��.�����Q�P�����A���MJ[��C�x�"J2N����wA�f�}�1����0�!�#�ݽ�������4s�(�BM�����<P��h��{/E&�s,��L���D䟙�g�T��>M��v�J�窟e��1"ё�a��I�J��P�a)�۔�6u-�`�̖n�����[oq�WY�udU,]!J,V�gͺօ����"�r�ɰ��ZQ�w�(Ʈ	�s��x������C�_;z�|�b�n)חz�M���y|�݌B� ��8���BJ5Zqn�$�d@J���؟�ރ�a���Zו���1�z?\{�k�3��+�g�s�7��`��Ȧ���������ᡧ��'�}��
˗-�����iSy�7I h窴�r�~BF�	ܱ{��n�X�2��g�D(3ѵ�R�y��|'�B��Et�5�@z���b1��e��U+�%�+��sk7�9g-��g�gv�κ�.�QY>XrpNh�sh+�ru���ĕ�X�v��j�5�P�$|Y��(�(�$J�O���Id�l*�M�����o��*e�!+R�qe���p������;�����m�~e��d�imi�\s+��1xK5=V/����N] o��
����o:g1G�]gby��_'o,���f�;k:�ݹr�7X`���	<mU)>gi⨞Ы'��h��cGʪ�.U��	]Mt�A+�7NDBb��T�SuH\�.������%&d���,�*9.um�|Se]6�,K�JW�o3��JP	a5S[��Z�<I����nE�j|��7-�����nG�2�^�|ڎ�.
,�V��6�
h�@���7m��s�ܠ�cNDd�/n�o�*2�:Y�"���ܓtkx(�g&4�(wq�ldQ��sp��6l�g_���쳦4A��),�8�m�%2J��B��}�`��=��{��g�� ��l,�2���;�&)��5�褭�~�Ԁ�wZ$�<��b�(Y0"*O�^"����"������Y�IBN��	�uN�9�:�s�l.���
~���ܔ�lߡð��Aظy��N��_dkk!�`xNl�F�����X� b=�x�k�@g4�:D�����0c�L��9�d��C)ʖ�y!ϗV��b!���H<� R�������x9�Z�
Z�L��/���|��h�:�1�/��g�Q�.��w`o_ �<���K��*�*~�/Ddb���5�V�bڦN�0���{�D�~l�b�^XolS�6��u�k���%��6�EN�ɏ�(�z���X+ii�{��Q����V��G�j�;�z� X�����q`W�3\��EI�����,>����y��8�U�(�RT5�*+��B^he��`�1��s����I\x|&�4rQI���~�1)	I�׆F{����Ш�X�_X9"�>��]*�������ϲd<f�ws98���}}�q���y1��\�H���p��� �s�h��M.����)7�����Ϫ"�ƺ�� I,�|�ˉ��/t��xC=�����FG���+(�&�ū'��w@��$�<�qWB��w�R�w�a��m���-F~���S��	:�2
y.�N]Ӧe��%���`���J�a�����
����,=�~��aW�l�
pBYvWЁ���=���/�YsN�䯹�2sRi�g[Z����_V���u��0���ݙ��(���\~�[����nD�s��dK�z&��`&m�{p`n�1��1s0WP�Z>�5�bz���1�֛���<���T�<�1�댮|��$�Fn�F��Y�J��z�HK6F�-Ϸ "�_G���S�e@�ql�L����?-z釦�hk���F9�[���;Pj��K����n(ҝ��v��>H��� ��A�8UE<%z�&!	�A�0j4F�cY��)K1����ie����!�����|>�?;��d\h��-��~
���dT mRS��r���'�-UQ��fG�28�e�bj����Cѡ��PZ��-cN����덫�Ct�L�kV�0��zX�5'<ڎ0���:����-c�:�?�e�ޠX�8��{�G�2��N�s�- �e�)��d�/��m�Ⱥ#�x��2�|N�Hf`��-R�Vd&�b�<�
�2���X�b�4��l��DD�+��O6T��x=�z��d}��(��tD�'T-��Dnʔ5����LϾ����Lϧ��
>#w�O}��w]�<��@D���1=6��{�ѸK�����?���Џ\�߅���S�=����f" Ѩ�z���B���t��1�����_���ݸ8Xu���('��l)jlDY���������D�Ňq±�\�����+��sr=���n��n#r��x��֗%�C�Q�Q��Y�-e�F?$7d|�T�D]f��-3;� 	m6Jd��>xe����Yꪣ�ZZZ񧍋�v���o����k�%�3�LN�5ɶ�	g����U��x=i	�1|�p�fc"�OX����ȃ2�H�T)���	��D1�$�a�l��n�u�뗕����� Y����8L�v�=:�"0x'�s�>X��s��iF��~2�����>nȆ�Uwa�!���$�C^)�x�k��C�SCu��,�d�:q�^���R�5�ɸ��a�;���D@��2$�����E$ME�ھ�Na����[`߾�iO����#=��6�Z���=|Ȭ��X�`aaq�A�<���Ed*�Slݾ%����A<����|� 'iJ߰s�S��' �nK����I n�֝��;uHU�Z�.�(X�|Ay�6J;��P13�b�Q͢�]�;!�Į��x�(�,�^��5�U�7	m�\pted��$��8�v�.Tуȏ�5O���J���@YH�����	�ңAq�X�D��ɫ֖�Z;��<����֕���p{���idpeK�́�س��O�@���l�6&9�ST=5��G�A��%�b�|���+�@C��C��4^�]ə��
�ʉKXn1������a��,�SM����wMr�I��Wn��'��k���j�E�5oȹ�Dg�4 ���Q�B��T�X�7�W�[�B��#Z��{��/",����*���}|�3��j��	�O��
�����I:��d���I�`C����-�y߃�-���C�h�|�}Y�4%dX�-�����O�q�jE�VGHZ��ЃJ�8;�ga�Ћ+`l�$�1P ?��r���Ig5̨�|�,Cص�@2q�&�8r���#sR�6J�X�$�&����B�I������y#'�Heaq�"-����������X��AQ昈��V~U�SE��2�{6�٣:�'�%�[�p Ԡ6ձ�?�~aBLV]
t%�B���D��Q�5O�ON��Ƨ�DƵ�
��n�N����z���`#��i��!����+�O��UP��H5Y-�`a1� �� r�fΊQ�6�dZXv#��䧔ی̚�g��A�3��V�/��*X�ʦ�[:'�	���k�ԫ��$r�P�`k��4���KoA�oc�����C4�#�$tj��%u�z,�<-o�u�R�L��{����*Q��`W���UT�Mku������Xˏ`2�ib�,�:��ښOW5��E"	%RZ�RZ��|A��|þ_�+�/��xI�$��}�9h�4s6�#݇a��휾�r�Ү��t�q�Q�u��>H,�&�f%����XSzQ�����k�>\�Q bH�W����]څ����`�����;>��",�+F��վ��h�W������e�<"���(�ԗ˿���LX��w
��?T��Y�܊�"J��� [G�Dki��@��V�������7ۥ��l��\.�Jb6��g�It֢�K(x�Q����J�W]�F��+�H�h�W��U��][�v葻&.�6�������ikH*խB��l�2���԰�b�)Gw�$�ѱN]�{�ż+�����@4Iǂ��.6-U�kdmT��}݈�CCä0uH��6�JJ{B�"{p�6�H�6P��S���.�i7��Rt��o��z=��W

S���%��j����!_R��	�;�"�Nl�HD�%?O����*�l�Έ��g$Oc������V���uW,ɖ_$�^灘�/U��b�~!���ZL��+�bִ7�Ī?hI�
���w�e�g�V�0<��_�i�,m'����[D+L�l�x!��*�"=m�lȊ ��&f$�O�u��U]S�8�p@DtJ.g,^�9�	� "!�h ��@��I~Gqg�Tf�-vO
�h%خ(��x��W_��ܷ3�s�>GY>ɧ��\i"laq��-?g���˕��K�(5��gQ����o�^�1\�r|r-\�� �{˛ �P�<�0���
Cؾ};<��_���5�5���g�p��>ʁ����e\&�{��;��k�����P�:�ı
T�j��2.8�/��+m�Qd{:jITE�.�e�T�`l~�$K@-�&���g'��c]GU�c0i6�c�Hg3�	e9%�CV�l��΀���p�|R�p��䦢��#�q<p	a�\7����	�؃]��x�]�ɀq��/M���d<(
�u�&����J2^ ���a�\D8)-�<�^��~9 �"k�Ÿ R`Hoqx�;,��тv(=EΓ�m��ǿ+��*��+`Ҥ�I�F��V��X{����̕6�&s���d@i$6�$�nL8�b0F���6�Lr�I#!�����l{;q�5�A7jh򚌢�8��0�$e��OFID��5�ET�8w�É��Ǚ�<Y��Vw�
�Λ�Ӧ$y��c9��ؿ?lݲv��݇���B��J"/�(���|��
	A�b-xv4�Srжm�Z�!�s=�^b��p]�s��?��8���9�z�h@3�5��_�j���b0�zǓC�B��t	CZ�"�?+�ȗlL;��ɔ1&7\%7V�q�G?� w,8jɥ���ü-pѲ�a��v�b?�ݩTF@���3OA���9�?�
l��y���lV2fz��H��ėodW)�4��1E��	.�h���?�b�����].eѤ�#�
��XE﫵Io|��7��X'j(��R¤���Lt��7k��Esj��yC-,�k��|v<��D�C�����^�esՙ���v)�9�h�GX	���Z���G�Ɖ2<
��.=	�#�E�8������Hd���1��;���z�W]�7���X�ڥ��@����y�NՊ<�;\���z�>r����YR�����y��dw�hp��{%JHFRפ�/99|���mm|����$�Irh�[�"��G�J�,ލ�I'���sfO������I��Dbd���nTe�}7�w��M\_��eVSk'��h�����'+�"��5�b��HUm�LKC���jç9?���Nߣ�K>q�׀��$��JQW�GI�>�&�Дkb5W桽��z�yp��Vh�= �d�ۉ|
��<�	�����!�� ��b}2j �_4N?�2����@~ ��
Y[��-��<�r�8��\��#B�>����FB__?d����08.k�)C�9qev"}U"au�C��_(r�^��Њ		[�C��$$-��Y|�Qr!�I��!Ң�o������|�1�W�f��J6��[2���?�"���]k�#H֖�y8�s|��7��_fd�܄���������R��9Z@R�����E���N4֤faq<ϩՂ��t/;�1J�q�R$�;��n�Qy=�@��� 4ژ��sX�4M���,�~��3�l*����_�w��^1�Q^�kI4_��������"�(=P��d�|S�����.�y�dMn���U0g����6�"�J����2��ߙ�"���r�o|�J�8m�>spZ ���|����� H�GR'�c��\.�"��c��G2���zH��X���u�Ass�k�J��s\����$/N̮R�窑�D�ũ��c�;�䪪���L���FHB��ދtD)� �����?��Q���(�!�H	Z 	���Ny�������l��0'���̼���{���ﱵoӡb���ڧg����jv�0aP��^�┄@���Ux�������v��Ew-�!�7���]F��l ���D�m�P�2v�o�h�u���֦C�ϭ��T�'y�i���S`���`�7b�8$�5�Ԅ��Z���8E:�v��M���p�~�),m)�������0�˪;�U�X	F�*�]{Y�8�y���V�{j�d�v�В�\�q4�/#�{7��T���o2F5(��f��RY

�r(.�����P��K�,T���漮(S2�R��AN�	CR�u�uqדo t����g3*��-�=�fx:�N�R����aQ=��<�%4���"�&>�������*��%�<]Eh��u`�W��R��+�٨�N)/�J�5g�U���uK���R�粼z��9�Y�{��Ѣ�^�����f��x�\��_�+��pB6I3�R T��,g��or�j���k3q��g��'V�҄�J��N���W�.������j��1t��UUE�nu�[��������76���tD;��v����Դ��)��u�>	[���ZU���6�8�۫�^[G��|O�,�&���ן�t�D�\BA}�<7�����ӈ�x(&LX/�},�-^� 7��w�J��OaT��]����`��5{f�^B%��C���,����>������u����,^X�#ޏߝ�G�* ��
(gE�v�=v�	_;Ǎ���>�E�V��+��ݮ`tKؔ�	�'�k~�9����O:�yu�F��W�W=�������SN�y�%��:�d�Y���;O{��(I���}�����Bc�$�$5u<s�DHk���_x�0�g�$l�ێ:d5��4l5��.h��@��U��[�V5#��=8�s�Pʲ�e��dK���H[��hT�=#��z��n�n��P��?��qF;� �ĥ� k������)UP�hQ{-W-�����`��v�cm��(�ⰡS����^{���r�j�e��e9�V���x�#h	�vy���q9��<���p\���`�� ����G������ǖ�'���O�\���M���~�����k̘&��'�`�M�ŏ�+,Vo!�(0JQ]`PF�B����� ����^7\�+W8�{?��~i�� ���N�1�O��uע"	�-\��Z������̹H�����pL��Z�)'"ŝlǊ��|��să�5xC�A�����Z��x]�l���%Ti�9hm�9�^�֌0�)�^׭nu�{�s*>�<.^��?���s�*`�j�
�U�!��I9�3���$�q����JZ�hinQ��"_X�f�Bz��X��O�E��<����X��ud.�f��f�ٽ���[�Ӣ��"���(eE��
jb��&�R����
,�v58����p���( �!���(�e���F[K���R��!#18ca�	����-R�i���:�b>��� ���
<��ݘ��� �����y���aˍ����m�[�}y+Z�{�����n�����R�x�I8��}p������KKv�(��j�>&��QW�)��ۮ�h�������/aYK(���G�����Q��G�i/(!�:�$����B���ë�V�*J�XTm��S]0l	-�Б�Lg˨Pt��rZ�T�X�LAr�phU��+��1��m�L�@�nu�/ӑ(@Y��?BS�b���8�����h�AS�zW �i�`�} ]�,�E���(�z�jV�ty����9(�MjH�rG��upY��7��GrL|�O5G�̈6�zqP�s�$�>G�O*?�_�aL���Dt��G�%�F1\��-�q�d�TeT?�Ǫ�p\��:uL��?,��m�JwS��>3y^{��ޝ�$W��W�9B� S�	���n��	l���8i�ͱ��͔謷����~n����jb���ﯸ[l�#�����S���o�l0�<������^.�
d_{�?����?�
V\;-�b������4�8�)�Iuo��=�x�Y�?LZ����%*��*d���p��d�������gҶLL�h�1���������ɚ��x��/_��B(���V�����Q��3t|�A(���SD);����	��`y�NEP�o�m����)zhtrh	�Z�[�(�J�nu�m.�'��W[�?B-dy7r�=�&l��sU#�[0e�h���Y�A�����%_;�0�����k܈�A��#�X_:�h���j���:�~��F�H��l���C�BS����̡� ��>ִ��p����k������*��
��,aڀ%-�ȩ7�R(Z��2��0�4[hEw  �2;��w�b����p���!����ci]�:]9f�����p��;��g�x��i�&Xe2�i|8�y���q���aW_�rF�M�����$�Žw݄1M���ܞ�J�}�l�I�(���/Ͽ7�r�$��y�u�[?X�ti,�t[r,4��r����Ah��"AK;�L%9S�Xy�ieHˉ$5�jI���T�.l9>�d�ǔD�S�6�))���\�o�7�j	"�0�u�x���_�� Ȇ>rhY��H��C�1�i��A����Z3�n�1�$85Q��;�,:^i�����s��i�;o�-Ȳ�PD����"�o��se+az7���E_ti|d��ނ��<���f�x��q�#��ύY%KR��Xu~鴋�!\��Z�b����=�~i?#Z��3��/��V�[q�OOƎ�)z����;�fɈ`��O�Z^�u��E�[w Ra>.aɯ2�Z���LZ��f�eْ�Ƞu���K��DU�=����ǫ/Y�f ���'���;�|���%!0�g�֭n�c�Xh��]�ı�	ݧ^	v&%�-�)"��I� ���+(�{DU�c\�m���UTw�e��,#ߎ�����_dߗ5�M�#[:�eGE�Kh�Y/X���� dǔ�ȋf�^OK�:��n9���б}:�ל�54������ò��d.����b��ph;vMT.ia2����d�J���k��wj(�h@�Y�� �*4��Nc�GF���ĮY��N�n���p��^��/��\q�$���J2�wj��6\W�4-����H�L_x�-�py	��$۵�pd����ϱ�~�⑧^�U�]��|F�bE�ouf�ʲ
OB �*��F���o"��i�vVQ��e�ă)2�Aj����y�})���4v�\��e ���[;4�TP��h;�h� �e��)2�HD��E/���m7_7NAtCO{�ނ�խ�M���7&y�:��s���ȷj ����F�w[�YU7Q�LB��ѝ��m�T��\�z_�+s+?v��/"ߕ�3��ή���j7�mcذa(��iꦎ>�޵�X�+��[ڶh}�B/U^O�LkH�xQ;NI�܋���2��K�ٯ��}�[���N����� w�҉[g���m�&�}׃���[aZ^�+9�i���6��m?3	+Զw�as��x��gP
S:��(9���S�W�?�&�������'�W� ӹ�>��A��#Q�߬ v�*�k�ɑ:(���� �E<�$"⁬�m�?�fr�~���W
ZW�ԂnQ�c�M�z�7�*{�K%���ÿ����)�K�#=��ԭnu��2�vYҭB�M�@N�(�K%F�s U �e3W5]Uƨ�D6u���$�Sqɏ����K����L�#��h���w�t	���\C������ݎ��v������IeuÍn*�u�;�y:�eiI�|��:�+��E㥶��s`��)�6ު@<X��SF��ؐ^��3Oa�m�CVMu6�`C\���q������~�>7ZfJ���Tc?�?š{N��ߋ_���ah���s�� �c~�.������cp���*�{^���C�Z�P�u��N8Y	f��O�sl�L
���D��μ����%z�nǒ9o�>�<��]�'*�:�~�TP�$fv�Lt���=�ݏ@m �VA=�����BD��к�m�X�$��M��~wŉ�wn�;[� R�Wc�|�~��=��Z�D{߯,���w�|Ґ%��k $���2�qC;#���#	""'C���Ss�����xB.R�2��p��rђj̊����6�8�h�(�ҮJa�%h>�p�쏵ॼh4`/Y�Dd��Eɯ�ۑ6a��ZL�ԅ�;�n����JY�����n�'�;n/����糯���h�"��j��\���(\p���ͷa�3H���̦'�F��:��Ͻ�ˮ�s2#Ѹֆ8�[��+/�QG�����I�tIJ��$6\��ӂ��F�>�M�T�YuC� ����%�Fey[d��6�E��9�c����P�����(hm;��K�1�[���Z3����j�^�)�<ƺ�QI�q��T�`Y^ԭnu[V˛�g��s��%�}51R�!ϱ�Ψ�M��A�q��z��Xk�t�R�����)�`Jm�6E?)K�?c/.�|�<t�/Q����ME��~�+'t�`_.#���ês��HR��w�+�s�(#�z���v>��yr3�{��'����Y/���"ZKL��t�rL�@� ��]�P����w�y�-�p)�˰|Q�!��;�M��n=�r�gY��,Jj�U7E���:��٬��I�M�u����~�M'5��N��I,''4��M	*�����ђ�;R����y�V띋m��k��G}����U�2�AZD�^�v%X�Wzuaߪ�[[���g�T�}u�Χ$���GZ}�J�M�Qx��~���zwv�^�%A!��$��Tȫ�9�U�JI����[����/ԭnu[FеdE��j�OAuN,7M�'G'�-�<�u��B	K���U��-o�r5��T�q��:z����Њ��������yK��0h�񗸀X�զ�,mA�4��&ڣ'���[�m��E���,Z��RT׭5����^��������`I�J�h���(,WV�m;�M=�ւ���a�hKB��z
,<o̘����*��.dͩ���;�*`F �E�Q���p��,k��'�>/g�wd���y�:�o|�D�Ֆ����K/�TT�����Q_�w�?�y�y(�,T��f��p����ey���NĴ鯡h�tfb�2��-<�!(�����9uT���\Yv_>�4�����F�q��ő_;A**5�#L��T��|�ZUgZ���� Q����dJd3�%y����+��v �yJ�1��6b~R�"��H�I
��`��$�H�Ӝ�]A���K�{�DKW��d�i1�u�[�>Y���3~���&L'�T�I���VF��N�X�ճ¸בc)!�N1���~�����QE��}������֕�'��:��"V��;W��)�t�h�Xҧף��7�h��$�.[�e���b�#hͣX����~��[�<�j �}�YXPĝw܂\F���C��Ny+�w?��B���S��=�V����.�B���#��e�D���a�RtD�M{	]{���P =��kO� uZk���+.�2�5'�*Òϼ�����&[ԋ�'�A�s��/�8���ۯ�������3�y�o�C�B�ܾzvG?�]�^�[TK�[�B�L�[c�����D93W��PO�;��H�V��,P�"�l6q�۷��z��P�s ߩ�5'On�.�a�}�4V�h�:�h����Z橜,X�S\+����V2�@����fYn����"1V勞B�4�Ģ�i)'��$/[�_.S��B7�AU�gw,�7�ugT����+�M�Q�ط
�j�%j�}����z�P&�/�N�DF��+R�X��zύO�@�>E�]Gȶ����`ÌM$p�lo��_~}&��:Jx���K�j`lH[���ƷO��j�(�Ǌ��=8N�,I�����.@�)��u��V��9p�L�f΁�f��='����g͗�x|o��,��1�y���t�A�?x�＿7��7��"��<2�<_��W�Z1�Ir-�#S�}&k!�����ș�,/�ٙ��Ĩ��&E5{��)?ō=��^�\~�-�&^խkf#)�$V�Un%�HF̹�-&~7�T�e�2/�kơ�~c7h��l.X� g�y��ޛC��؎Uc:��1����)�<���$T��������]��alu�a415���� �U�)��1�C���5��HcFƊ9�YÛ���,o<��;�]4&{�>8��D�8A�ܟ���	l�J�Wo�� �=n�5��ͩs�y��&�7'��9��K~��ͱU_����$�U-[}m�rf�뎙c4�j`�R͋$8�_�i$�ѓh �p�I��K�6�/h`�6���B��$:�>ӑ. �H# ����j`E�ȎV�
�2ه��V��czB�%&�Q���˪���АP�k1Bl٬:�şK��F�{>�Qt:�����?���km���fP�/3�c�6��/WS��o�����k�¢��[iՐ�2\��3q�Q_ǨQc� MF7�P�#|,X87^�W��|aQ@�l��e��?Bk�����IJZ�������}���$�x�K<=���p�@.)G
jt��8��J4���Qu�kmS>�A�A���q S��y�ml��ah��N��~S(y�$c�39̜����(�˴�9� }��V��,j?`����P�.f�	f����\�H��O���Y 	u�5W���k�����͗;騝J'��T�L<1xQw.���`{�� �&���F���jy��7��6S�"	��A��e��\���zP�y���x~g�_���4ǒ|7�[*���0���ٷ$v�{x<ϋ��\_�k��g�*+��	�U@�;��̛�ٓI�'m��D�xoۊ����%���VP�G7�]Qհ�Ǆ*����P��X;��j]O��Nh-����`41\T��+b
�������W{2�*cB$^JzWb0�= �|O��6&N\c���W�RG�ꨜ"
^�;n�BB�o�>��`��1X�d>�x�u<��%�K�t%���-u;=7�EjL}����s�͝�/�U�[���NЀ�:�B�Uu��$\q���'��:�/!Le�����N�^X)F�K4�rDϑ�f�}bG��L�,>v�i;-IY�%]VM!u�,�Q�U���Yyf(0]�h#Yg�u0eʔ6@TT
������ҥK�h�"|4��
O �L@u %�q[l���j+էNDSS�|�b�
,_���f̘����@����ƌ�s����f�m0y�d�{Ȑ!�=�����«����ӧWk�1N�<�IH ��v�a��6èQ�0|�pYn���x��������?2y����&��k�ر�݆�,[�}�f�1�=�.\��]����&L��I��{��O>�$��(��A�П�
'����H�d&tmGQm�9D��X��=�
�,UO���kڭ[� eV��6T�W��e���;&154e=��ZQw�ͮ ���g}
�S�)�aDס��-��!t9M��i#C�~˼ �=>��5;W�!3��K�����O��W�)੹p�	���$�ݍC
�ZY���x��ih)X(�HG�����"R���b܈Jl�r��93Hy��cc} ,�%b���"�wJ:5��a�%�� �%[����4('��tCo2�W�>�k�J��myZ�qu���F�n]���9�������{�裏��z��������/����l�+�h�F<�@{��jy(i�>��Hp���߅�3g���.�삣�:
n�ax��s�Q�䷿�-^y啊�u����o��m|~�ϫ�m|Ϗ9�ƾ��/�㟷��^z��i�~-��=���:z��J���}��`��;p�嗣���G���i����L�Si9�7�xc@ Q���~D��ȣٞ/i����n�/͕� ���	b]��d����zH�����m���K��s��M���2�r��n�3ܠ�B���ϬƲ���MP����$@�P�C]p�L
􂫟�T�B%N6C4_�j7��S2�y~���k�c��12��U�
4�(M�A��]��x^K\#ףgiFu(��~�ͨWVxi��ě��q�|�F�iNK�+J��x	�mB�5f����:uW:6��-
�
P�ch뺻!�>X�p�{��}�0H���Q1'.���S�CtRp��|IV�_(5��L�G�)��G�(h�XP�dWZ��s��߁`�&|\�ɬ�^C�1c�`�}��A�W\��{�/�����/c������d� �P�ȑ#q Q@����a�s���o�6�ǒ��3�8S�N��g,�'&A=��\r	.��2\}���/���^{�?��x(��k�fy���Ń���[�SNO�9����\��O<�"�N�-<Pu�I�o�&�s>蠃H~���ŬY�*�]u�o�g�3߿��o�#�����_w��+�4��c�h~��k��C}�B��?�:r��8Ey)����"JAQd�4�	D��#�M9�L��qJuvL��T뉳%�>�MiA�vݖ.��6�����F��{W<�	ꀌ� 
��jj�g��:��	�'3�Y��.��t�z�"(�n��%�8ϫ*4�4+v�W���Kٕ���|���W��Nbxn����_�Y��P=�$�GY�R��A�!'�[�@���jS�hyI��i��0�
�a�vu��^����A�R%a��+"���3Ʉe�.uv����4�S%6�|*�u[mu��2�M���$$3�+	Z�?묳p�7���FO��"&� ��}�{�(���'�| �:C��d2��e�a���{+��|��W���I����w�gϖP��~(�Cz	>w�u���}�}��Gx��ڄ�y�<�;�8�l�xkk+�x�	���*1b6�h#��0�m���Z8��q�	'�ts=����n��N:���J5C�����x���)��`��7��>�q�p�y��_��\�����~�u�u"���Áda丐k���)�j`de�褐*4���!cC�V��<2����*��f>�z�E��Z0�R �/���ǈ��c��NF)Gڸ'���LV��(��9ߤ7��iy��8Pθx�չ��7O�:��ՑY��/�=4	���v�1�k����ڶ��wiP�\M����ELR6������2W���0p;]��8� TF�%�3�����m������ M!gլ�P!��������)u����%x���a��<B�\�u�wY��=��P1����3�PF��V�B*��ߣ�L�h���ʎe|��qh����h_fѱ��j��U��v�V���<�����x饗%�̰að��d����}���,�Fz&i&�'iK�r�!�ww���\w�uz6�������v�M���---��O��<�sĻ��8.s��cڴi�=�o<�\����?�1��~��4y�8��\�Kꁜ�5���[ŋJP���orG	�	z�/�G�=��ӆ�J���?��ωs��ݎ+���-��v|��Ӌ�h�� ���-��"��Vr�9�M7�T@(ϝ�c#Хg{ Y���^5���(��*)��Q}Υ��
����!�j kT�L���)�����",'ZǢ@�y{p�:�[z��;�a0^�@�U�_�M)q>9�X���oP��Q�G�kK8���[+IO�#�X㍈c�Z_��9���E���g����,�n�ͮ�%yC19,-z��c��š6Zw֛8F5Fn6�}����l<��˛���Ex�W0���8��k.�P��
v�����d�E�N��3	|�>� �rC�:��ܻ�3��5�r|j�����U��3��I/��>��S�z&Тq��c�=$��o�3̫m�����&�������A�Z����;�w�}�,o ]R^��^���Y��&3�M��1�Ùg�)`u�ז��ad���O?��Z0I���N=�Ts�I�+��ο�����g��G?�^[5���w�}q2��</3�?���򼸜��2�'0}��G���?��Ob LN*��I(�N���|0����
��7���$E���(&�P�y�Ts9��1�Z�L&'!�ln�Q�?n��FI0[�d)�b-˖��yZV,A�u)>�p���b�V�0��Rʱ�*�¥���s$�qR�J���:V��llo�I����8��oi}�����+i�Q",/G
}������MR���@���U�n���Ǔ���6�
;5b��%Q[�T$��J`���VE�<�'ϲ+����!���XɼL�>ZN�,�/����y�$�Y�����s�DC�=�5�G~$�p��l�
,]��.V�
X�=��y%`�I��g޶�L |�@��鈣gF���f��bj9�7�jT��F�g6���JQ�����|�i�loI>���wϒB\��$Ȧ�$v+��!y�0�]�:�����)|2b��1:�9s�H����<���X�;����#�$�2��d�zr�Ɍ�$�Jn���o��7`����P�䱚e��gڜ;����/��'���s3���2?t�P�\2�kC�jhtS��������5����FP�d)��9~���4�Z	V�ћLo7�9�����C�1��S#���R��"�V#$o����M���N�[�N��~�na)r�eh*-F���h0&G�=o3�ur|�p�c�3����p�5�v���*�����2V�D�����V������:��sI�d�>6)�j�W$�4}��;����&T'��
TO��N>/���|6�nY����f>��O�g�˃-��xo�
}C�2�΀׳�&X��@[��ԫΠ�U��Ϥ��To�>W_0�
�H��wVt$�%��\�_���ŋX	()�d�E>(=�i�v�x���3�i�1k>��e��7�}�{�mo���+9����e�<��}l������$.��km��g���?�y�{�ܹ�%u���؈�fҞ�aɘ?�A����ۖo�%厸E���R�NJ�S
��al��]_�`�������߁8g���2��33���3��� �[k�gj}��bw �	�	B�a$�Ͽc�nd�p��Y>�Ͽ�?�m ������k�~U\���G����:�nj@��*D�ѹ�� ?��V�^[2;��H�+��y�M7�W�Kr:/��,Y�d�GW^�������N&�'<`�@e�as��}j�&+4%����o�S?3UB����{d y���:����o|z�������Մ$+a�8��zFlI�#�`QKV*'Y�h�-)="e�(��P]���JgeY�m�Ϝ�V��}�͔ͤ����w�QF~G�(��ɐ;�������3���cRQuh�?�T�⋅Fh��&G��f�N��h@(=!&����ce6�9f*i-�(�}�e�j�@���_�\�4k���m�0�ECz�W�����|q�}�!����h�Nh���_���d��h���v��-?BU��\�8{��W?���'c���V����D����$1S�^����L�1<Q���9�\u�U�h��=���L�}�d�z2do����Jf��j���3^F&c(��Ӟ����x��L�ɤ�'��	�N)+#��p&��(�eΟVZ�ŲJu�4XG��VXf|zV�P���V�>�Pph�Ъ^_={)�5�&Q���ժO_iA;׭nu���3lȋL�N�db�SL�9��C��Q_9J���9n�( �)9�4�$w�xe	�ȕ��'��1{�����M��������k��m,�p��6254�7`����O�y���p������Z�̔�����M���$���1V�D6���J�&s������DX��NkX�Sխn�v��� ��$=��	O0��4��!CEOӔ�4�E�Zz���EX^ �U��|�br;� R����c#ٔ<��7p�w�)jp��
��������� �7�sd���?���n�ϵ8�����w��;%���Gy�TC2���,�I^����Z]�t���S��m�(�	�eUG�?Ac�*V��.}[������;���E^��6-�~8��\<��УIUo;VV�+�$0bB�VI�U�/��@�(%�h���&:�%�!e��d�����LD�)����T�A�̌�3�'�=I�B�)d(~�uוs�WT�d"�=���=��V�1[ޔ��λ$�OK֎O���������D�&�C��z���L	�����0z�{b���� JJ)���]ԻZFQ��:ui ZP5/�m�J{��P��K�'�ҾG��C�uot����:�O�OH��:^����V��cAe+QQ�3Sf$���Ȭ�m�&dڵ�ݎ�7l�� hjt��Ug���	��G9��&3;��^O�P	Nf�^�u��S��u�ޜ�ō��d�ݔ5�e����}1�F.O.$KgRX����bu"V=b�ο��o4�>n��Gn+Y�Ș���JPk�e�t�~{��焓J���2ɟ�%�+=��R
gS�p���m4Q�f��CO���E����x�����_�`A��o����֪5�:X<�emڿ�t�V�wiu[eM�f��E�= ��+D��v�@�)U[�gè�	�ô��$��ٖE�H��C��羴�0�ܒ�H�գ_�[,	J��Օ۲- ӁK��WY#�$e�L_�	����  �O�������	B�{
ͷx�
Qi��\�ze��ֆ�I3��hkֺ��s���(e������	Dr���)EO)ۉ�ϼ�<�I`f����z����2$O'��'^yӖ�.uSG�KVA�Nj�ztt��Xh��*�������N��׿d��7iw��G4�g/e��:�^сl:�\����K��w'*�n�BA��D
�MP1ն�nJ�l���:��۪��4���m�4�4$��R�U急"�kB���5K"}� �EW�&@"��!A��I�v-�$R�N8 C��zb�Rʾ��n���Z)8��JF3?�f<���$��ѻ��㏋�:+�{챘<yr\��@�|�s�=Wj���/�����JZ��u�]x��e}��&ՈX��y�\�}���E�����
��U3�I����ˌ2�o�����Ӄʲ��z)<Vփ�:u�|�w�Nyđ����%Y���$Cu�M���[*�
QT�j#s6�%GM���-_�U^TM0cz5�0i��r�$� ϡ�I	��[�u�[���yg96K�
n��j����K,Öbar�<���8xw6cU�J�NcI����W��Y~�x��� ��GTu��D^ռ7O'��ŋ� ���'�x�	*�$x������N;�$��� �r�!&�/�.}I3���SȽ�R��t�A��w��w�ϟ߭�5�޿�o���o�����$���p?���6<?^+�ߓ
ƣ��z����$0�^d&xq;q�U�����`�W,�!�`ǭ7ES���'���+�'3R�o�1��Ǟ�BM����D�V�>�����J:�ŵw<�g��Z������A'0+�.��_m~��;��j�_ÊHڃ�:�@��j�O���m�.zGQ�{u��ڒ����i����d]�I�&�ԍ���[@���^},���er\����Wf�sY�Կ��S<��anB��M=��4ȶt�Rn�	ZL62���xt���l?	ܙXu�׊V+A�رce٣�>O<�h���u�[w�Z�|U�κ?���b+&�j¸�������6'�%E�S�de�ĐQ�"<ۑ,~;��Ѻ}
���V��2ʖ��P=�%d���U���|��_�,0��(�PN���N�C�{'7�[#p4�G�,mP��3fT$�u$%��/����Ef�o��zj��������3��|g��������L�g�W��jΙ���_�:��-����=�#5��v<���LT:���%۟���K_�o��m������`�/�a�����[�@�/@�9L5��	�۞Ձh�>e�? ���mB��k�Z^�w�M����(遫>?�x��Ih�'fI�x�3z��ϝY�ƥ|g�}6���:�xQ0��Iz��s$��6`	F	h�_������J�	$k	Л
F�T"o�pY����Y�f��Ӕ��K�����K�+��Q]MZJ���[�G����$��I��SR�b?�X�dI���)��A�=�Lr��Hb�U:�l;O)�G��IUnér͆�΢]�w\��@��}Ч�D2"����{]��T~��6W�v����ױ�V�@-��W����$��ȕ�#�zF_x�x���ٖ�_<��?�X�E��1&�0��f��	���G�n�#�<���'��M�8Q����4���~f�'���2R_��z���?jT:�D�k�綱zA�^Yw�j޴�|[ [�W�/�ݧ>���>:FL���&+!ߔ8�Ne_)�d g�f����o�=vuC�aS�9���	��T�kKH2�av��,'1O d�M�|ҁ#{.9_���ٯ� }]&��T/QݺoqcBvY^�����A�'׆#'ڡ�s�#z�p�n��Ɠ��Q���1�ċ��tD+��%t��x+�mO�1�jG��m�ߔ�
�L��n�
��e7���T�����q_�äBO�E�]�fv�F���ˈ�3,��^{Iv��92釉G��n��3�\���k�Gs��?��B�~,���H��i4lio��wrZ�=���'� �aqS�Z��O��@M"�Id����6ׄ�as�1�t��]��b�Y�6n��Y�V)5��y��%��5�����;"][Ӈ��W�U�����c�L�=qJD�-�e8%r�(I�-q�������1��D8�Z�A�y��d����\c#�Ɔ&���?��Ќl:��/ ���Z��(at�Ʊ��jg����=ӑ�e���qj���fS�vx�dU'3�!�5G��(u�xp���ysb�����@̺�^Jm�wQ��6̖��d���ւ�!��,d>�~�UM�tgA�J����e�j S�1�U��"�n�	i4��
����p�^�h��^
�[�F�4�\��A���U0$f��ͪ7W=ώLD#�mUdh��ɵ���g�^_�VJO�#v��ӛ�n�n �5f�|��ߏ��w�Z2�z���U��c��I�Ñ�F���MV�jY�d�z�MX�E��4�QÓ�	>Y��rR�����8��� K�)ߓ�"�CZ�k�_C&2%5[WWk[k�Z��7��v��c�	4��h����z9~/<u��������2ްP�o���w�~��e�����v������p�	�#t�ꕁλu�����N�x�E�\5I�}�L����N]�>�a��%Ξ���b3�7��:u46Y{"FWx0
��8cc
.^�w?X��f~�yzX�C8($�)���n=7S�(9�,���r�ؑX�ty4KEm�Y����R&��w>NԨ�S�5�6,Z=�]7B=���ׄ��4g�՞Ҏ��t�+�g�1Q�<��7�6����t��������嬄Ф��I���	q��片�xC�9N���@�����v���A�(_�G�l&�����6�f�oqY��w�e�
�*�����?��<?J2Q�F �Ϸ�~{ �R���2U��:ݵ���/����Xs���u�u뺙	�)i�:��T����ډ�D����fPl������\�@�K�Rl�N
=e{����� N�5{㸗rsX���C�t&���:�,�0��SH��S�s�����r��p�_/��!9XtB�E�V�|��^-"��|�*a��&a{�j�[���(�(��Ĵȱ8Xs��1���&Mœ/���3?Ċ�R�������&�m�Z�;�$�%�N�7�-���m�m�`�kg�l�f}�'�=��N{����4���q~��y��/���v�&*�==7�m��`����/��4�0��>ok��<b�k�� �t���Eϓ�9Y�Ǆ��=_�\�ǲ0b�O>zj����˞z���q���z*Θ�g��ӘQޙ���b�;�� N
�3��,G�h���:�,��2�^~����䳔��mg@/��;��c�y֣7ׂ�\�Q����i݌šs�h�d���CJ�� �KD<J�x�]HK" e�މ���(1�O@�e���}zy.���l�N�'�}zrI�yceh^���ǜ�k�U�{6�އ�t�"�H��Ys�Z�[������*������L����4]�}5 y�da�ݶ����!Ū2�xK��>Ŏ��P��0M�-`�}�������1gy�f�5>ϱF��3aq����	�|�m�Ά'�f�'�O
XT?x��TIa�T'[�4Vc2FZ6��I���-�Փ��iK}5���眴)��Z�����F�#P��S�U�����p0���' c-w���3�gΜY����.�zL>��c�6m��V>�3Y-iʔ)8��#��>���`��W\��D�C�,��R����9�y.�j�|�ɱ$���2��L&q��O?]���jP<���]5�6���~޼yr�f���t�Mq��7�g������.�s:�֜`u�/OYJ~v5�#^x�>��H.%�d����=?�o�%l3u��iP�ڼ���Y�p����yJKj$a��8����'s6]g���VMy������䪿�ї��� +3��
Z��|��x��R�����qu�;�33�v��oc�:a��I�H�O��+��9
�P��ycƯ��6�sf�.Ԩd}��Z����ru��� ]st��u3�l,��Kr��U�_�7Kr��FHK:��dqq��:�/��������^�[s�#��֢�쾫]]�O�%�V���滸����}1LXP�\�r���N'�W�hq3K&:P���7�Ӄ)�g��������O��Q)H�ꤥ�C�O��n�O�9�Bպ�.����"���Ჸx����O�(cm��%����Iv�)�N�&S���(��JX1$�ק'���cb�K<f���Wm��ΌqSIȀQng��d'�����62i�� �ۤ���Mv�Y�av�d"s������r��' %_�� �?���m��	�	��Z�|�Ü9sD˔��療��hmlh�uZ�>�K��0���5a�q-|jf_��_�y�wc0���j�P���G��P��b�-�4�U�U�F4�dR�����u�Q,r)�G��u��&l1jk�e��q�����O��v�&�	�(^Q'̢Z׎����Je�G���V=Gͭy|�(4+�Ub-;�.�5� �������%�s��0�ɉQk%�c�6�|����W�J��yؠ���+���MH]�x���}�5���F*:9O�a,�SۊQ���s.��q*�G^�ǭ��H8�X�V-��#~̕7ނ�n�^��~��	.rg��M Z�2���#���T�;�zb3aM�ԏv�X�Q�- ڃH�Q�siGY���I�)�R�4Z8�,8�,	���h�䆚��-�=�e�fj��d�0�0�M�1B^��K�"�G���G�}��В�6�A�M����]/�.�=�Y�g�C�Kz�}�U��8�Q5�?Z�Kv���h��&�����m�k��:��*z[�k�<O�Y�q��y-��Y:+0�䙕���O�[uM�Ȱ�l��gq����I�շܭ���:�7�n�1����jU{�3QR���ѩ���i5���Kp�aފ򪭍U�u��'U�J6�Y�����V�%ok�NR���%�>���)���g>p,�;�3~�<��UX	D���(F)��ϡ�aP���>����,-��2�N�`0`�Y���Xk�dn"!���z-+�(\��rS^P@.c���Y�e#��Λ����;��p'�V= J�Gh�݌��-��W6�رtC��l�$���*3�c�!��@D�N�q=���w���m��4Z�)��TE�P���<��-�B�$D��h�� 	��*5���e;A�GKm�P~JEx�T%FYV�7��w��S}tV�}�w/�5'3,i)7ʲy���d�Sې��բsJd��t�N0JvІ/�3Kp�S�p8���L6��Iph�S��=��S�'�7N����p6�-�
��;���o`���e9n��sV�|��eI����w� ���}�w܁���5�w���3����H�)���%u����u�)[:b�0�e�cYFo��.9��6��&��L���7��U�V�ϡeK��FL�LI*K��e��ĘU;�>��O�iMM=F���������U�O�o7*�	�1{ޜ� ��A4�-�l�v[o�	�򹭅"���~�{|���h�2(e����B���Y�����Yy\]I�����1N���O�ϧ�'[�-���lLXk-�)G��\p;T�Px���"����o|\s��t��Gt���*rn	�O��CZ��G��;���Y�h��N�`�?��l�;켗\�g�=�{��ƌ�Ra9r�֠
�"��ͧ������ڞ�f$�Y�誹NF.t�Ί������\\�[�YMQ5F�M?�j��<�:���fR.�^A�*��͒�NZ�WF�r�=���W������(9H��qjY�9��Q�%)�p�2jPo�
꺴���z៤i��28a+�
yd�ڣOە;��:�U۬����,���C�C�/�	1�nB�A�N�v�`a�`EӲ���J����k�ɛ	��[�N��l���%i��?ܦv�P���z�d��s�:5�㦛n������$�0�M�$���>��f8��9�{��y���x�|џ1n������4t(��1Z�AS*���%�?k�p&_x�Ŋ��q����C=$/fғ�ʐ7�.y�|���d�#fƿ�������&�
 �|��e eR���>}4!W훉d�}��7E+���1���c�٥�a�8u-�L��\C����Z[Z��y�z�m�P-���W�US��~�xY*�Z�<��J])&����Q�Q 91��Q��5o��JR��o���y�R�,TF��J:RVc�mG���X�р�$��V���D#�#�~uI�EO���ӈB�������_��_7�?O>�VBKj̦�����/|ʂ�Gy��ս��8����jߌ���5W�(p{���1��$6�#���A��ߑbC�Uޢ�}4��n�u$ٮ��4H�+��+p��'6�z�m�a:�B-�tݱȅ�Ȫ����NB�}z6C�t��kTi�z�ɭRp�)��o�36�x\qɹ
�e�bt>J���]���>� ��;ECf
4��^8���!2��Y���w�{��?�W��nT碀���jsi{��W�m���:�f��߮�����T#n�|�3i�w�M�[[q�G`��V�hs����#��E���0����㾏�/��Z�3M�򊋱�z�8���0㣖ޟݢN9�.;l�M7��*� fw9�%^�* Z�n�x"k&QsS���s��������Pt+��r�A
�8��O�3�[/O�B�#��.�%z�� O?�"^�������D!��vI�0���1�G�C^"̈́����Z�Mt!�%rޜ�J�R���x��)ZO�Y��U}�,�)a�h�듬�D��������I~��PJz~���e����{�&�yW� ^����(�>���Y�,����]���l㭷ފA,ϳ;�Xi� $a�<ٱ�*� qy�6�&���+�ԤI����`=�ft2���ݍ/�w">�A
p�������>�����GGa���H�����
�M����-�?p/�j oq�	��],c�zRkރ�[���x{�0?iF��S�kk	
'Ah&�t>�.]��NVz�NC�A믿���fԷE�c�Y��@��N��iH5❂���=1-�nD:�o�p*.��\�9()0�J5��j���:e>~��뷫�N�Um��N㗿�)N�w/G��0,�-����6_W\����G�%p�V���/:{n8�P_@
.�5.�ߞv2N:�8��ђ
j`�W��'^�!�n��7X�<5K��(�����kO4r���hc��j��ƪ��a��F,]��%��~���^Y$&�ijtо���г_�ps�h�{�u�7��%�47�h)�����;xࡇQ�mt�X�`�J��x4�7 ���낇B�t'j�g����ڌ�����D���ߣB���X�%AeG�ʓ���b�=d��G���*[l�T��I��AJ��u�	r����7�NwGU�����{�&�^ΘU2c�/*�i%9���
�h��G�PPhB?)1�^{�����������_���g�54�R��h�JZEZz,) h�JY֓	�e9�Q�֒�@$���y���U������s�4����qȗ�����x������xL�~�-�c	g��2!_{|���E���,ȕ��6��nO���w�xȏ$5?��}�pZ"{W�G;�9A�`rJX��G=>�^e�K#��hq�%��쀜�M6�����K$�vW���t;��u�"중�Ʈ���=��t�\�yL?�k�䌶aǮ�-�v��/)�Fu�o�å�ݍb*�VՠƏ��6� '~�
Mj�I;%� ~�w���\��\��n�s�(�=��3~���1n�x��_��c�+� ���o͞/@g�Ikc����ɩ���\n0Ʈ� ���1��Ɵ�}O��� ;��f�l��
�>��sX�x��n$��7&��RA:a'������+���?��g��=E�Fޟ-��D��@�����,჉��F:��$S�yM�R��c���8eohO�d�'��tV�����CN��V� �X�6#ϸɪ'�<2��z��m���du'�����V�"U����Fs$I�^q-O����r�K�o[����ЙG���ɵ�]%���֌���/�)��8-Xr�a�W��tEr��X:��U��azѶD�>$���YƧ�$�.�7^�����/6��>�]s,6Xs4Ǝ�m��_>���7��s�����H,���$%�Ej���zf��������%̛�����\=JT�4�ڑ:6{�eK#S���u�V���N��6ƍ�@�dB[��(�D����}Rf7�i?�¦S��Ŗ[���GuDj�:�@]$JC�3)��u�ŉ�Z�!*;�j�V�����{�)G������n�|g�l7T��y�������=�tJI��&��f8v�-D૧�O<��d��F�����G�¬9���`�����> g���:�!���'q�q{a��v���\�����l�� e��k��7��5	�=�,�<~}L�<V<�3�zG���z�R/M�g�8+җҴ�Zq�����o�� ��UZ�Px2�̏�?NX����m�3[���T��k�r�������0�!y:�F�\��G��v�Â�k��/�&Q�UGD�9_(�i{�J&�����U��I@�N5���uf�+X+c�:,���\D�X������j�לO�|LB���>�q&����K�<iW�c�In�=A+A�:̙�n��Y�%��J���T&��C9!Z
-�-�Y����F�̠���>NcF��Z�)I�>��W�K֖�&)�-�Z�����w�ВU�2� �V˩���o�W�O�	]�NJ�o	[xR����ӈ0X,^�ְ�8��S4(��E@����Yx���p��1��8���ř�����O�1ǝ���P��p)6_7��&O³OτTdb�!O�NēO*����1�ӡ<�t*H����C�Ǥ���]54�����a�]�R��jB���Y�N|
��|<3�q�|9��.�m�d��r@hP#�kx�T��/.��AC�+�ЮQm�.�eg1l�X��X �^[>_�Y�<F<r�v���ųI���u�[G����d�ٸ$#ρ��V_��nB>t�Ǟ�#�<��V����2��m�C�Ԍ�����oǅ����u�{�=���_�%���5�(�>K����6������w=�/~a����꫐j��b��6���{�,�� ����-2ï�fʁ�{|Ͻ��j]�J���=v�Lx�-�*�(`�Y�A!�T:��g�}��'d`2O��9��t�M�Z;pe;�0�\�ƠL�n�-y�C��O����k1�_�Z9��EN�K���z$>	s-9!W�g�����~;����	��� =�LNt�Q)�d�*��v�%��V�JrTY&�����~V�]��� )�G�����rXd����ɷ�J��.]��iE��i&� 	3�ּx�|�f���j=��w�מ�ŋK`J�@�\�W��g�g��82Mh�"I>.�}�=�|ڙ���`�1Xc� ,j������7�{}�������)���j�)�1�(�'��2Q���X���'�z [o�ҩ��P��<�)�P�F�/�㡇�ǐF�W��4*]����0��E��RQ]h�,ՉX5z�Z�nAPc�j���}k���7�X���hS?�,k�ſ-�z�`1o�J�^��w�s/��$����7�ǵ�z o��L8�KF׺��22�4d0e�$X%�=��p^��ڮ)~%M��&�=�}sw���&����"��x���f���p��xc�4�i�����L�5�<�?���>s�jN��`�q���i�9�C��mDn���fv���qu$���ڬou��oUŚ���>'gI3�ҜБN��z|xS�L�E���ldv�j /�gP<\��^c �{�O�o!&�;5y�K�h���K�X�-����y��$M
��>k�X�>$�۞�g�C�-r����^�>���2���-U�s�Tcb?�J��7*�L����m�i5#�;���υ�Vك�If+ݪ8�뾚�5���l���,��QޒdI��Y�L
Eڪ�%�@#�`j�Af�js�x���pl9y(޽�	)�XJ�WS����'}rV���UD�҉�I�Qx�^B���S]����٢�0���{_�o#�����G��S�#�f��}[_W���1���d�Qd�솚���o�e~1=|M�����o���M���h)=����B�E�~��s1b� ����S��kY;@�h��￴��cf��M�E�bA�!��w���W���G�_fZ&���n�Qh��9A&CA�>�_��x�}�8��Ga���~�0��ﾍ�y��t��~i�(T�YO�zPKxOHȶ��"ah1��F�萹kR3�f��<����m�5e��/C�Mc�5��'��u^�=��c#l��Ƙ��Bl�����:��̔�.����v+��׎�$B�G7�6^��oj�������2�j�(�:�Ƌ�n�qy�Vr@��R�F�k���u�F=xE��^�+�p��"nrv����q��1��c�0��{�&��A���4���H%B}m���-�>�{��v;�_������a�SO��۪}-MMkn#���.Ay�u��E���{U��V}.�C�Ks�Ȕ� ue�JT���w�kIbf��`�m���<?����ѧ�A�ڔ��u��"��deU@��@@-9�?����b��qġ�	=�;E�֑(�������d�H �TP8�%N	�RX��e�/�B�<�^�<�@�:�P�����#-�W��t.8
�D�|>`�A=�X�Sځ��.�DaW^z�-Y�7^W][M=Zg��8���`����8�V=;�9<��|��h�s�������{�����1f�1�t���կ�K.�>>Md��C�Z�l���[�ms�
 �����+�n%�i�%D}�.�n��4(��.:��{ 6�t�1h����l�0�7ߘ.��C��B�ȄE�Q�m.�fC5:�\�!�W�_�9=p�����!}����o�%�Fߙ���k�����[�dԫ�O�Rb���rvh��)�����ox���`�����[숵Ə��16��.v�j]w��8�S0c�b�W�Á��Rn��{`��6C�3n
-j�T�%%�1����XT(b�}�F���˖�cl� L��4�K��������aҔ)��뮷w���H:�l*�ο�Ä�:��+��BFuu��n']�@'��y�-��
�LJ:|?*�kv�:+l�Z��NN	�PB�_�x�I�H�ڎ�,���ڦ�p�%�D����k����
e0����G�+3sN]#���idU�,�H?X��#���'�Y����9�(P`�+����GN��g!��*`e������j�D�bz�dHXaAA�V3"6U�8�U����g�����x�G��������g�����\~����;U�؀�WD6�U+��U�b�'��|zjJ
��y.�]˦4]�ж˒���/�楿��d2�
=U+�r��mEٹq�S%�X�T_������x^��7/T'�3%��D�(�%y���/���fu.)���-��u���@�}�y7�>�Q�{��r/%��Q��Z��?���lz`��Ȝ��=�y�4'��@��Q���ڔM���/��>ZL��OT� ]@���ZM��L4�� \�󼝦��d�,.��ױ	�2͘A��(�s/��VN-�!_X��~�d��ꋱ��#q��N�w���3��^��1o	J�+�fǈ���F��GA�.���o|�|~�o���%��/%"�r>@2�l�G��tA�&A�ߡʂzRdYWG�R�ڐ�S���}��6֞8�F����e�1�u|��l5rД%w�ɖFg6�@�}\�mn�*=���{gښ�@ML
��x��y=�͛?G��]��ܖv�}�� �}�m��;����!ۈ�+�}E���d%ԥ��s���?}����]uS/��f\~ٍHY�`���?��b�H����cO�����x���k����zU88��2�����#�V6Z
�*(���>����L�&�r�l�M������$�A��I5���B)4�$�N0�1�1��{���S�{�{3;�ZU�`�^�֒vgg�̼���vnsg���L��v�n4�Z~�������i��s����n����p�>{�!�tҔ��l���W�jq�J��1c �S!c�qK����e(�;�˸=�P�eT�W�2���h�y	�y�tkD���Q�_�@���s�g������)uX������:]iQ�HB��5�{OJe{�P�f�P�bL��Lq���@[;܌���CO�|�.��HN�s��=�B �AL�%�=F�͏�CV��d\Q�Q�SH[r�TV��Lw�	-��Z0�ҟ9�_�XD.]'���L[)a=�y�^2�ΰ	�K٭�}��ۑ��R�>O�/�-�B1�J�G�c�҅
Hd� �<i�F>�!�L�A�á�"b�mV�|��l��x�h>�ӃεP�"����xu|Y8�*ϝE����,�+J���E7c��L(�)c�<�/tO)�n�d�
<��h�~���PƳ
�R!�8�ct��dm�$���g�q6N;�x|}Ğ�r���.��2m�L���#����ь,ͩ�<vLx��������ч�3O:��p}�`�R<3�i<��Sx�9Hg{��v�q$���<��PtK%z1KR��QUDE��W��HM���I��<su9˖��{�����4)ZC��b�L��e��E+�C���v9G4�n]�|�ey+[HydH�b�)\��n��.\��0e���&�\_��eS��	M
)�Bޓ^�A�K�7��ߵ0��c�z�D�T�V��RΧ���i8�7W�[��F믏u��a��Ǉ�?ƈ�C��A��?/�C���b ":��}�@/���Ӱp�"8V_�,�'�)`���V�l�m7�&}�O��!�|MB�^{�v�����V1q�G�>o	����+����b�0����/�����4��P޵%�i~��w�B ����ʲs�u�]da����ㅘ���f�>�?	߭M^s6j=SV����6�.h��HKJ/�	hU%R�I��R��D7��(hk�]�l�C7t��4�"2��A �)ye��K`�'����uT��_V|���H�P�hZ�\Z�ҍ�p�+��:L|����E}�#�f)^7#��K�kA15�t�A�^F�I�R*�S�=:�oHچ 6>���B��y�*��A�I1ߋ��Zs�\6�-n�ݪH��T� -��	�Z�(QP 8p�hϋ^��
02R�3��,��@׌�82`�};��g�e\\��0sC_K<�<�Z<]����<�;�֬��3I�Z!zя濭�a}�g���n������{�Q="]�W������p��7�{��Őg��`��虩�E��|p����wPt}<2�Y<��X��y���8�4�6�ft؉�r%��֣�U~������!�bO�j�muA�"S@�D���RSP$�NC)��<}Z�����o,�|��-����]f�1-mx���}S����称hY�g�ᅗ[�e�4�̓8��s*����5�<� �G?�L�N=�n,��k*��h�EW�8���>1�gͿ�!���eUH���0*W�洄��ЅRL�)�D3�tJB�l�?=���� �^���/�L��Q����w�.<�HQ�w��<�4.{�$���SϽ�#�����i(&��
)��V��G3���y�0l4 x�3i��sD��w���s���$�W���.0�}��>�r��H% ��j^��J,[����e� ���w7�e���Y�bĴ.W1��h����9\EX3��T�!��K���WA���j1L.�M#ŋv�}�W�	ފ%8�S1uA2ny5v�n���0�5�~���W��hq20l�a����4��u3-��K�=��&-J2ӄ-�ʅ������T�ei�=�����脿\7����;�ݏp�~���틫�x1~��a�+H��//�-v�qG����K/U-Fh7��
<��(�r�=Xݍ��;��q�٧�\Tn,b���k��;��f{9Wף�<����
Mt���?�n^u�WV���C7��#�E��=�<QW�ʿ߈����rC�C�^�z�m��u���8M M���_^t>�|s�,��5;�����p�-W#K:����W]�{4���G�TZ�_'�x<.<�4<��Gpٟ�.ŵ���f	�K�BKM�R��%�t�	`�8u���]��[@{��+��ī_�k�+�nf����v�~b�t������@3�˨H�Sb�#7�m-HsT,`Z-�l,�$�"9�e���J2���,�j�J���M��)�0]K$��P��C9ΐ��O��j��'}.:ͣRV��A`�,�&����6%�4�O����)�|���M����d6�W->K���B0�/��?z��&���&��&{v#>��)�t|��fti�l�ۤ�l��g�n3���h^ь?�.\j��k�-��K�I�=��q�ߔ����M��=�N��v��ʿ����]���dm�s>|.��\��A���$�7�� �c���k�t9���ۣ�v1�/���E����������:
�>�P,�sύ���lNsh�G�j�ʛ��)��_Voh4#�w)�`��e�<��B���+k���֨ͺ��4Y�)��f���n1��ږ��
OM+�ݗ9n�
��Uݜ��v���1���+6���P�	H�׮��,�+���q�?��g）�����Zo��V����?��Jԑ���oM� ��LR�9�tI_����
��?���?@��3�S*B�$��AąI��~�e��+��?���b��ڋh��F=�t?�R��0	��b��H]d�κ�㸣��{�fk ~{�q��/��矌���%Kc8t�y�H�����O`�ۀ-��w��GL����gO�,���u�5�͸�����hL�,9�e�&3�tx
����G���+p�C�@��#��.��T�M�VJ
U���z^��������'���ѿñ�1l�=��k�����<��X1����.��/�W���z��,<� ��Pɧ�k�ىq�)'�������~�f�j�%6Z��-f��1�:��6ҭ�CY�U���UFk�J� �(EA��4�8�$ PRUX���Y. t�7ub�ʯf,)^	�;��Z����[x:!"�jhL�6啗�c�З�r�T������-C��(����%�D��A�؊}B��ߌv�E��xm�7v�@G^mnR}�]�A�����isbq�`h`��
�ȧ�����ӱѦ["��˔%�5���?:n#�׷wF�^�$a> �bY�¤i��(�vy�ae�m�*�m�q�W�.XMGE[<<�̚�`!�z��(�B�Og�ЂK/�
[�#��ǅ_�s.�P��9���Q�-1w�,\��F�YW&miR��n�v���׼O�-di��Vt0s�ghj�߰�@�O�s*�J.֤Ǥ���KN4��
�FR��K��*�uEr{�R(�U?�|.Q�Pu�0�6��Ji�I�JȖ�	o�����})�̓�dr8���Ѵb.��O�ڧ�,&O����g�r2��vz��q/`�˯���>��ں�0�47-¾���_}_(�"��%�K�+R�t)|#�BږaVU���2T�8IZ@�rGm��T�E賅��_�B0sx�ٱ8��-��o��:-�}1u�B���r��x��%���㿃���7?���S��'3��_wއ�O<��z|���)��B!^fQ����%����z�:n/ة,ƽ������sbgh�t^�+��i�=�7W_sRp	Wc�+o��g^�7i]��p�[��;��?�0�Pz��x��'���" .�4������]\�g���G�+�m��� /�F�%�
	�$�FzC"]Q�/��W,�먮e�7��>�X4�b�hm�64ccW�N�ѧa�݊Ԝ2g���~���J���*�i6\��峦ZÇ򿓆�j!�·���]~n	tK��Yrv�#�ܕK�@s���M��{oM��N��e���L<�����v8易��+e+�O,�<��c�:u"���H�6��!O�Iٻ��^~uV��M�*{9�w�Y��S���4�l�uuXM�9�� ��?(��
�� }�84��O>	���8�d��F1�����q�]�a�Q�B�^5���P*����8���p|<u6>Y�����p����9^|�Cl��m�ƄI�h6�ց} ��*�JzRV�'4�V90F������O�����O~���E�/F�6S�RTކ�!��A�^�9�ܩU;�r%^���˜*>�� �_�JU�Ahؗ>��޻n��/<��M�ȐQ��ga�������X8�3�R�������_������B�\�"�4��?rv�C���������4�0e^��B���N:��\ :4�B� ^4��{��%c<�nE�J���%���@c@��[D2,˄)i\`�A�m苽���˛����	L��=Z���&�Ƨ�|�<�zq�����o�\#0ꥱ0��j�e�˒#���~���w�,z����3x��!u^��si�o�����^�}C��	K�Mŀ\�~DR� K��=N��4E��<=:Ʈ��?�旸鯗�������9'^���d�V`���1����@���dm�(]�$߱x@5SDI��~���EK8]�,m�s9T�P��i�Uv�?a0�W:nE�XRK��}�c��|���>���z��}����G
�E��2m���+�yH).�e0jv!���V�T�pU L9���|	���{@�0yQ�VT�:���g�t��1d��PHc6���ѐ��l�l\���Ff�馛*�#���ys��i{����OV�������2��(�I������[\ �ʞ�;'��]��~����de�� RqZ��0��ҍ��B�YbOF����������%?��DJk�?��78��}1���hni�_W�rHBU�������֛1ꎿI��&3�I�������)���&)(�b���|���j�R~�"�x�_�bƋEebN��oD�4�w��j,'�(�]v�%��6�@*�U�LNϤ���F�P�����:���O:��Y'����y�$��ē������|�*���o�b^�t��'�Ws#��"�R�}���9�w޹����SH�a�j�iR왤?B��p_�����dƹ]�������e˂���t'ٖ�3E!�=�o����%��o���?��o��yn�&�K���*?4ʏ��i�l��܀�t�����%m��pq����sQD*��:��1kaRQ���.�Ho6q=	g�*dZ�(�LcLӽ��=_�(��2T�a���w����n��NA6E����;9��,�V~I�k�i_%���� ��d)g�bf�/	 ��0�mM�郲�#���N/۶�uf��CG�C$Zx�\�-��f/�9�BW��	F%54bZ�j-q���NT`��ZfJ5r�?�
��Xս-b�IF!E������3�
-8v#��N9fw���d.3���	�����}E�t��wJ�R����Y��T3�ɡm���t���ƼB��-tᘧ�L�n�B�����d(�;v�s{3��M���5���
�3E�g.[9��%�)dH�~4s	����u�9x�wQh)�5���XK��]R��(:�A@���!a,U�ʊ��Y��Ӎ���"�";����Mwe�.6F�O�F�-]:m�%+
���,w �'�r�ˋ��6��vq���q����o��V͗�آ
uYxT�,�m1�d�:�#[��7M��!
MK1�1��?�)�-�8�3�AK�4z��3N8/��������m���Hգ@ڛ[��(Q�[,t~�|mȐ���nF���B[8jY�{�l���eP檋�����(�6	����)~���M����Y�q5l���>��p��܍��K��t�JB!4��X�Oe�]�SzN�̃�]�,���k�L��,ā]ר�%fΩ'`8}�44�dsԱ���0{s�*�	S���&]Iיo�k���u��̬��S����8�\N;�h��/�i����sVJ.$7Ehη����:5��i$��f���[��H��+��S�%{������reǺ �A��Qx�J�wX�� j)�� �x�7���H"P��n�o�B�0������釴��}F-J��D'nTt�*���I"�MGޢq��.��Þ�K�O)6DU��Sh_�g���ѯ⨃����Ydm�iQ�K��h*ob�&d����쐔Y��W�x�7��K��4 �J7\5��jZ�N��+�Y�+��~�Yh��ȸ�����mw�Ͽ��A]��ο/��K5���A��yP:`ԓ[������V�<���n�%c��8wN�.����b�%�
/��W7��RJ�6))��*�uA���˰ɦ����؆F���>��������ٺf͚A ��_�b�d����޼��M(hC��BӞ$��(�7�]@g���k�JɠPڽr!��>g��9���jk�4�/i#�@7Sа�"�K�vG��6���y�d�P�3�S���d.��iH����D��!�[�d.�y����>:n(D�����WTh\�ʹ0�+��34c�!;���˰�}G��g�ŔI�+.�5"�a���3�v
M�AZ��]C�`��%xf����w㞇n�Wߌ��{���t,�U[���"�=�4$��,��!*�×Z�ηLx��C;���6VxVU:M{{o?M"����j���KΛ�<�为c�1p�>O��c��+�ɘ?k*�'_��}[m<@�O�Y$����{f��O<}Q1E J��/F�7&�\����2��ii&����U��'p��NtS�1%�_l��Գ�����eSDٜ�u�Z�� ev��=ŕX���	��j�\W������܌��D/��#��q���W܄��\�M��E�!tC���ا��^�ଋ0{�'xo�|���3�`٢<2<��C��w9&K*���8����3�Xfce�4�wѲ<�����^F�I��q�y	�#�]35Q�.j�O�Ԓz��,-�^��Q,��e�_�{�y%�v�q�y�.�C��5�'�g�sf-s	d��HT�qݲr!}�!\t��pķN�#�y��{�#vv ~���
G] )I\'��W����ǥ�я/�UW�I����o��;����Eq�,&��uw��p&�=�u<��C��:�?|o��v��WH�*�rP/���~�G�v���'���N*���/C�S�F���Z-0� ��?d��Hc	G1GF�rOj25 H~�̻ކt���(z^�ZP2�#��'�(尕����?7Ӈl��w�����A)�[��z{. �����=�|,l���k���)�H��F��>s�e�u�9l�*�Ш�8W�Wt2.�3g>����M�U:R����m��^ⵧ�&5Y;$��
1s>8,���Z�:u&;�\s�o��K�K"�0h���?���g��2���w�w7�|�Y�Ch&�x��g���/!�f"e��f+�c%\ ���OP����?��V�'� ��t�9��_�0�]�I��P7;����4�RaǱ(J�jN�B#@h�lvVƐ�ӟ2�}|��e�ux���$u@rJ��<|�/_Fz�^E�t^��唕���߂�����^��_BrHO^|я�e2sO� d��	�
v���8�����[��o|�H�&�#?��Lx�ڨQ����	|6k���/�����]��h_v����rn���Y��A'O��_��
\���q�=w��s.F˲ S�ɪ&5Y[$*F�?�����E�Ҩ(+�5sNW@���UR����O����.�"��Zɨ�[@�-��\��d]��3�g��A���V�m�����\���K�Iu����<L�6Ӧ-&�L���r�L[��<��[����D叠,A��G���-B\�$��#�1�CI2���yt�V�g�	-}5$�$T��d�d8���\�s��?�ߕ��2��r�
x$�;�8K�ng�<�Ț�ᄣ��m:ה�9��C�1r^i��/��Y�F�U'=��D�~I�+/i�hƴ�`����sd��t�>Z�&�A���O��A-H��Z��S�ž#�*���J���?8��
�e�VL��c�8���!��h�(��aVRN�J�E�mz�;;������P]jt�.1c���Kc1|�'�\:f�;h0��7m	��ٝk��
�4ԓ^�$�r��q�`�=�j�l�O^�#�+.�� j>o.Jj��qOc�G���F:Ss��d�~B6���;��3��-����B��OZ�UN�y�ɲw�Q]����j��f���g�d��n�����i/�"��bě%e���.>�ӂ���ާo�T�2C5'�7���U@�,֔(�>b�Q�(>�@Uc%��EH{��
�6%�a�~��� �IM�8)ͳ$�H�8HQ�:�?��H�
J��l0d5Uڑ�����SʩT�jQ�-o��U�&�R��PWr?�W��R�N�c^R��B
�a��ʱ�86E�rƿ>O�,�g��$��TG5�q����ѕ�� K�?�g`�'_S.չ��nXJ�ǉz�i�EQ�e/�)�E�oXP@vY�Qq�4飭=���?7i_�⪚�X��X������I�JYפ�D�ʬn� [��s�)
*��}���D���C�R�e!l�r���-i����S�ےeDy��cEX�^D�@� �@�Hy���$��Z4��"K��j�75�IM�X�����%�߸��V��LTՆf"*~�V���
��3ձ1�6J���Ռ�tYB�ߨԱ�H�t��N�e�ճF�٧��EE���<�����2���8#v�����ǥ�uZW����6
B;������gJ����+퓃ra���� y�����)�����A�~�&5Yۄg����C5�aIM��{��uU*��V���|������޼���@ךi$��Kn�Jg�39�����I�D,����<"���W�l�J04�/ȵV|��zdI�������e�L�*_������O���u&I�5��nKD��%kS�~�+V��sB�ue!��*�U��ڷ)���n+�s��%��/At��L�h�Ǟ�h����s��L#A�w+�#oGߏ�g�2TV'���Dab�e�QJ��2T^
a���c<c�XXjR�5Ix63��6s.���Z�*�*]G���0H�>�B�f��YEg'���筶L�H�1S�L�"�gbҧS��Cޗ1k_n�#m�px\�_9 ��'Z�WF��+F� 6ͨ�v�`<��r�{E/	~�WE��)m�R�]����% �'oW�1�h�� mW�����p���Q���B�s1��MJPm�T QA(y�������'�4�*y��4	#7�캧�_���VuϞ�|en����ɴ܇(�(�Om<Ǳ��00ʨ�J{�ǭܾ<�́�r���+O(SX���(��8w�n���m�y�x�'���Z-1�v��tFRn��7��P���t�8y��_D@����3/�W��U�J\�R�ϳ��,�0JO��Ѫ釠J:������,,����#�@�e�%�[�]�R�!�nQ=��}NR�_-IX�"��?Y���N��o%]�%�'�0J��|�y���T��$�G��˷�vj.vs!�`�������Pe\U�U�5�r�n���<j)����1ϫ�[�1ZD�(hZ�?#��.��U^x	��h�hMjR��ň
<D*��V���H��x�5�8w0��
t�J�֤&5��WC�k�ne��d����6��[{AW}m�њ��s��,D���۞Ǭ2��V�Ш�[umBMjR����K*�$i�(~�������@�5�]Ij>��Ԥ\<�\�0[DX��麮��u_��E�M�A��KO�W,�0���T	m�о���"\�1[3=kR����K)1��v������"�STnFʢ5L�1�q��j�S[�jR��(uu�p��H�&´T/�F)��JePt<X�-��Uz$�PQ�0H-�'\	���ㇰ�9�`C��.Έ��9Gԕ�d�j Q���d�# jE�5馬
4�������%N���<T]���v1]����F'�AjR�/\>E�&��|zp��YⱓN�߇�<��b0�6�Dݨ�v�r��^�r����I��ܸ���Qd/j*�q�tMjR��tVZg��˚ ]-
�}1k�������;�<�����[�p�$;2UP�uAʁ�j���"uo�YMj�vK"3�.T�L�?��h�Jۺ���d7#�e�i3�#�o��+I�������{>)ˊO��Rj��Q���pi�Z=�PT���IMj�s����L�PhEN\+n�v��Xt�OX��tr���͸�Ռ��Y�!��_�{6���ѫ�)��yV6�`���Xޔ��*��|%�xN�<�5��mK��J@Zѩ#�U�k��VN�
�O:�:'�nB=��\Mj�3R�B�6~�D��	�FӀZx���	"���
:�ЖK�S`���=W�f��-#-�>���4:8�����h~�0?)����`xϊ�uN5�ҚG�&k�����j�Bo��Fh\���-���X��d�Dݵ��w�����l�r�OH/�C�f4��15�b$���J��V*B���Ӵ>�<+�~�����x]�Lz/Ѝ8h���7��K�܉S����0oi�PEYF��(�IS��\�(����ѴD�V�/�;��!<�Q�VJ��V�]�5��꒤!e����=���#�����q���|�W�MJG@+(kP���k��j��Q)���� l��Ԥ&5i-�m�͓��S���G^��9�\�Uy�͞��M�͆~EO�+�8s!]z^��֤�t��?����E.m�.6�1b��w���A�(��� m.C���q���};lڗ�1i�<����X�wh�d�&���t:]���(_�z��|�ۤ<�W�F� �F>�w�凞g��duHy26b�п�e��ݐ6�m4ӣ�I.ѲN9]�v�Z��1���/y-�� ���׋�eSUU�|�5�ɪ�O�S*��4~�"�����{�~���K�di
�\�O���p����j�?w��{M�@ϓ@:���<���{q%��pذ��_/� �J�>fFB�Hm���l����.�b�AYl������:�E�kg����i�纍��8k�bJ?2e04�~d�	5 jR��#q����i*VE���U������b�%��0{��
ʕb�7�&��*�c�"|�DI���n���7�&5�HL���{�-�\��:�,��m�=k��t��{�y��D/�u'=�l�F�,�O��s��ڢ���8�
�1dP9l���HE�n���e��0?�*P*ڧi�1�^��b��w�}�g,���4W,����G���Y���^ }�g�	��_>ĥϹ�Z�Eh��g�q�Z�IMzLĢK@����el�Mc�#�w�,�x��yP�s�n����,� ǟq9�X0,K��s���-��'�\�^�W��h�"���ɧ���Q��_��L�Qt`��(��#�КԤ����Y��_w��_3F�mf��$��*�fVQ���~=S�K� RB�f1j�5Y�	�1�tH t�u�8j����&`8.�/K杸L�fF
ł�l.��)��b٪�ޣ�F� Z��)}h��3Z�~3��F��̊��
�i��h�/�M�z�k�/��S�xȦ,��B:aӦS��  �2MYX�����������-�"���vʉ�u�l����tIe�2h�yI�/C
�؞��c�P�\�"��4c.�zvtLh�Ya�&��r�"�8�d4�C	�$���y�瘶�X	��y�Dead~(����e�&5�ɪ��������OD͊�f���t�R5��N?J�	MI���S'ׇ5Yx
��}����3Z��+tL>���r̋�#l���y�]�X�t	�{g�y��&�� M��=��a9��=b������u�x��li{m�q�MT�g�	v�z�N�D��66٠��݈��%��\���pyf�[���Mp��ptyA^���b����U�*��^�C�ߗ^����[ֱ���I��#/,�Y1x��$<���`w%ے��]���l�}�7�AVU��J�XG����s������(����Ԥ&��AXz%D��E�ȣ���oF���K{��m��}�DR#)=~ͮ状͢���
�����u{e`�KaZ��=)C�5���|����`���.z����1�>�(,Y<w�qri�@h�D�9�hy-蟱1l�-������7P�'�V�6�h\G\�t*=�eyh���{FHy�!a�Ͷ��7�Y@=�P2[!�iZ��� �t�s5���g`ʜ�h�m��oٹ��;�� �~KT�ʨLBn{����Z�O:�KM>�y�Y<+x�h$J�@��H�����i�畟%��'{5-ːE�3R-I>L<���������a���ut�P�5y�YL�	�5�ɚ A;�'� Ѩ(�]ݞ����/㊦�rT.�h^�0��T�)^⭦�#0R�K2�+�B�l��{�`�1_7��}b��u�0~*���8����uF���H0T��Aج1�`��ӛ+�N�G�6Oh�@�O~~)}#-�1E�gK7?_��?�ѿ�Ƹ���k�D�L�I�?D��QtW`�-��O�b�2W���=[���V�JO�\��R(�L��|��9��/�{팁}St��`���-���΍3��:-r!6�Ɛ[b��0af,lF�W�C琒�s.^T���!V�ɡ3�
+���58U-���{v����sdJ<�f�;<Ќ2	����RF4^�/BJ���`�����+�a�V�wԱ�����ӈcj��Ϙ?���P{G�甧��M]t��}��/��h�u�ሮO�r����`Ҕ��{�VQ���]��E,}��Mפ&k���F9�E`T�&)f;��>�F�6��"E:�!0x���g;�,��Y��S�L�����_<Bx�7��ό�&}�z�؝=��g���͗���#��y�|fC��U�}`�X9���8b��,X��O8�7�P�70c\����`X�`-R��;���:�fҖO�*@��`���q��~�З�|q���l�TO���^�RVo\p��p����~�{#,���X-b��a�[�eG��ڭ�.����d���cʤ�&��.�l[m��-�.��4.�y��2��6Z�9#�Y�U�ҁ�9�'�o�;�s"�&D�t�h�&߸p�s1�H�5(t2-{s���-L �Y�����Ga)HI��$:�����ЮmR�hm�X�h�4|��`�R!As�#���!U3�S<�5e>�1:�[���Po��^'��:�C��Q[U�ң/�u�_�°��&5�IM�a]����rl�����_����l�7  ��:4��_�c{����s�*B5Tkf�Y�F�l���o�Mm�o{4���V������#�oYR���S��}��	��t�����w�97�~��>K@cW%���=8~36�x2�+�[�C�#.��=���l�����H�2L;���9cG?���¼�ix�p`o��(<��c��7�F�hɣ�/%����rBwڢ���"�K����1K,	!�	���;SCX\å8x�!�|�Ù�3L`���3#�M��Q��e3���I/y=y�y}AĖ�E�nt�ԅZ^|���<sAjҡ��P����S̓��]���nt�ОC��K�"�4%_5��\����Z
"Z�[QW���_GFa|�҈���E��t�a�b:MMjR�5U�O���[�}������B90��+��G��B��v:��6��n�)�w��#@��8}K�s��̓��'�ȧ`54b���{g�����'?:���>�<�\����]6��BG��Q����.\t��8p�0�|���H�-��	2�q�Ȥ�߇@�R�LSL:�hj.`˭����f[��[�y�cp�-�����E�^�=��S�胺�I��]���v�X)�<��̀=�.6Y���#Lg��7�g��W
�>�\X�f���y_$T`�u�ȦiY��H�.�Ｙx]_�h:�\?0�Z��T��ęH&�1�Lre)�D3�6�s0Ä%`&r@�	qF��%�a5�&������"�!sFYlP����S���i��fż�A�3$��6�N�IOh�:��3��,Q�"Z��D��b�*�޹7�t݂�IMjR��]t>��Rj���2<��ch�wXp�4>�� �̚��_�|���AX��لO�"����p�z�tL<��x<��s8��c��O�y^����Eˬ�n���eY�;��k{4/��'���G���n�M7��V��DB鶉�2 �t��>�8l�>�e;�Vt�Q�ܑ�,��L��h���/�SvL�ֻ�^Y,w�vi�JU��#�>�"z��?j���PԔt��4-J�X��A�����㾎u�CW��V�,]�cƌ�̙3��0�0�s��L�/�!�o�9�೥Mt��=lU�K�c��h,(�/���T����*� d�^qP���w��9��lVB�>��9�w�ɤ��=�ܮ�6����v|���(a:��<��
��v,�L�����Hte�p��q}5���S��C�A�QH_�����߶T����M۟�URw��
)K@�<K�����&5�IM�d�}_h��5d�M��R)�,�yzϑ*Sj_L��bK"��|p:aJ�i�N���b�-��v�9�;���ep˸A�z��.جW}n4�,i�c/����?���x��1ݘs���.���2Y�E�&�8J9us����� �%�?_hKb���A����9��P79	]46da�����D��������h�A�{���E؞#
ڽf��\��²�0<���݀ƾY���e�#��s&-fAѡ�D\��E�n������rwԄw��.Q���"
CyfS$��G�"���7��S�}�P�G��q�7і�[��d�g�쵅n�GV����k��>��d�H'/7�3؝�Q��&�]E(��v[`����&���gU����,�`O0B�6͈�[�>A��܅�0n�k�h?�E#)��u;4�#�z�h~Ϫ��B���J=��n�z���1��F��_n�g�5.��Ԥ&k�H�:�g�;����q��q>����g�RE8\�D˽`C�u����Q9��p{I�P�MC�gx�k8���f�&,Ԃ��u�� �M�8�0�y<?�Yθ�_������g����!y��2U� �*o�	Ź_�өJN�fiW4R��*  ��IDAT�9��C����e�83�G7V�(t��Xo`��|�W�iQu�L@(������3Σ5,M�ؐ;���$_δ�8���~����+�E*�:�P����t=��-r�=�)tGdy5U�,w��t��FǙ'�]�^}A��_����=>w=<
n�x�Ȣ�d��"{����sNö����O���y>��	���x��pإ�jĳ�nA��8�[�cz�&��6 QF"�/CP��08��#÷�=H�*�����M,�}E0�B�G�?g�m�k��ꫯJ�z�L��z�aZ嚆L \�����Oc�V@4T���/�	�Z���j�����++kS/v�MjȘx����ˑ���?�N�ֱ�.�XV.�c���1z�q�C��: .@ѿ^����k��1�1�/u���i'WTW��5o��yn��X�O|�T�����&LzϿ�}u}̜>/O��}v��\Sg������a���B�U�6��Ny�.^��u�ШW�Z���D�Y.Y�4�*�M����/H�\
����)�@���Z3n7F�7(b�!���i����䥴P��Yg] ñ��pԣ�R�,T�ε���Ŗ�|�������z+��[���fh��o1sߘ%U���k���Y�	�˟��|c7!<����� z���Rw�=��ɢ��a�}�-�{��`����&�g�a�~���]wǅ?��z���,�i��0O��aM�J�Q�n�i���IUm�DW(��-H[����juѳ`.Y�%"�h�>ө�N�Or�V���5T��� �Y�	tr��w����~|^lW��1׎N#5���(fTvZZ$�ڗ��)[�u̻>�}�0��Wq�~�a��A�1d�~Xg��1l��q��g���_���.&\�[Bk��d/v���8R�@�!G�<��vNr2w�q+�W����M{?�x��W��NCp���o�G,f� ���E��ѱA�M	ŷ��>R\:�t���J���3�u\Qq_�M�)��a���
�
�r8���xi;�fϗ�A��R;0ڨ���؉�2 :$g�e-[n�rff�R�j#M�c��l��~"鷝�мz������"Xx�Ig��{nA��8��C�(Đ�����f�T����a�����G���*�.��{Ƿ	���\u啸��6�Œ����n�q҉'�H�o|Q��~uɏ�ֹ�J0w����"�Ѻ��v�m�3N9�Q'����C���f?�e��Qn��A���M������� �l�:eB����KL�v�*E?x���"�,aR��F��w&N~�J�,�Vć�Y$��"�|��kh��v��(�/RU�U~4�PSdXtG����;%r`kU��,$��V����]�U�:C�k�[�<[�!�!���1i��CA�MagyB;__ψ1/)k�3V��tW$\ʋ��}�c�G����0l�:y�� ^���l�(u&G����ز��l&-�l��ٸ�_�q'���z��k�ƛo��������w�s��F�����8������3�_��8��,Z��--��y�G����_��b��^�D�� �v���Mc�"]��}C"ʲV�k�����Y�	�'��B����ً����D9��9��ﺰR��K��LŌ�T-@�!�oFc#������+��X����\�NsC�\�F�S���Fh�uEx[����g	�;�Q��?��W����!��c��!��G��#8p0�XHe���(�� 0ڐk@�l\�ƹ��WwiRXY+�0~?�� '̜_4��?L��k����O�v]��o�X+�-��/�1/!�$��n���'�s�n���g?���ǣ)= -4����)�Wb�ܗ���/����|\��E7;�^�xIzM�����C���0��U�����b��|���J��ko�f6����j;1�~�"3�ys۝�୏?�\�J�<�������B���V%�m��\�h,��c�Ê�u������|���1�Eť��� ��㪮���@�|�?��1h�Hb�-�IMj�uQ�����˦c}f�։a��^{@p�t7S�_�O�Bz-�<�����}�n�t���E��y��f���˵#`��q�/��}	m�}z�ceG�\qz�#�ה@#*���k�5&�/y��{������O�氰�Fa�����_�KC�;������n>~eJ<f�V��;TL>����߆��*ˍxx%��[��~O���qBۈ�J᷇���:���$�|-	~2c�0.ͱͶSW��@5��G�kQy"�*�1a�>}�7U"��*��Bģ�b����7w*i��d�*�`�pW�v�dp��X��f�mB���1�@��u�dm�U�׬^�L������/m1ꉇ1ꅗ�ؽa���p��OPY\��W��%����5=_N D�"k��8}{n�%v�a[��ڼ����'f��H���E�������9%�c{R9],.�{dK��т*@4�
O��w"��,]���8t���	�X�n��Μ�S&��������.�,Ty1��F���I芔��#\�	� ���ɀ��BS�}��Ԥ&k��#%��p�>�b�u�5��m�}}�ƌ.���@��OgbҔ����V�,��K�Tb2���iB}:E�dK3����E�繘Z�)�`�Ίj=p-�Gʭ��0-m3{pΩ����n/�����c��C������F��ȿ_����
f�S������\�3�s��x�)��;Gv����*JZ&N����3X!T�܎�B����'`�mw���lTcd�pT�Z��N��1�~�)�i6��p�:]����YU�)�nK�	D������Ũ?�R6��<�F�[�u�~6�`̟7�է\��+%�'��X���:x���/�aG��|��zM��L�~�/I�܎�J�Z9�l(��W��0S/<aͅ2��LRE	D��u�q�<�W���@?�.��/@b3A���m Gڤ��K��e5QCy�"�(1&e��iC����X�W�F���"�ayy��`��_�芸g�-R�i�"�ج�2#���5�6���'t(�0L�D�U���4�>zfh�Ni� Z�x��jT��Ѯ�Y��Ԥk�;�o�1�D;��@�J����V_�^Z�p�Ѷ,xk��LD��)���Q�-�-7^��K
�:s|���M�e����iZ�����X��������9ӈ���t�#�"rV����<�oZ/%��_&�>������GPp���g�vűs�}�.gi��x�I��t%��e��Hf^vO� �D���.���1o%�/0�WZRYxm��"�z�aPh��;�Fof�*�{�d�;xⱇ����h\���i	?�,�2k��7S����EW�[E� N(Vsg�MB[q����t��MK�Yu���P[f=.���������o�$�=��@/��gN����^��>F7��E�� ��a/N���I���&����.]dU�"c��ՀY��>k�w(�5&�epC�٩��jJ�3�䕓Cq�%)g��a�˄٥<Ĥ��s���~�K�UX��Vx u,�b���B�,*v��^\�'s�/M��,��k�J��i�l��{�k����^�qJ��k�ͶS
�V�<^�J����0�Uꀝ/&�IMjR]��ͰB�Ŕg?���8Zщ2��
��,����-<6Y���!F	3�0���v�a�����Y0X�z�O�5���^��p
�/��ύ{��
_����y�u����G���G���Эc��6>x�x���2W���i �<�Է>ő�}v�^�2��F�%�\�D��f�]�Q�t�iU�oNk�4�c^��9b0�'�Ys�M�Msk��g������3�A���Q���S�M�X6��w��<-���Ԕ�����O����O@� ��({��$53D�JbU����]���KHR/��̞=]���E�dYs�ͭ�9/�&@W��y�.�x9�������>��?;o��<�����{�3�s�8��s�Ѭ%0���L�)_=��'��$��͸�'�9���3���[رD�A���^�i�p����{QW��0v;�l3luK|nj�`8�B�C��kR�h[��rX�sE?��}455�v�}��9^}>qt`�]v%Л*�����XX����1����p#l�o��Z�Da�qϣ�ȵk�פ&k�h]�HǶ��ҚT��� ��3��N;���[o��$#F9�N��;��<�\+G�3'=�
	fj&�L�-�/�f��민��GވEM.�T=|�ӹL��r��^z-V/q����0T^�QO=�c	��z���o�%��Ы7
�h��sšc�^Ђ	��C��zZ��h������m�
��:4���ࣥi%L�@�g����ؑbJ�\�Of�dN�*ږ�!��I�	aɩ�MQ9y�4|"Ɯ�#bb��y��:t�4�,?�ln��\��+W"�3����/U󦪦�$�v��pk+�c�ܶ9�-�ț�F��#�2�����6��7��#6۰W]�+�D`t��D�;o�c�-7����0���!T�i(7���|3�[0���b��$h���翘Q)�PQ�׊XwC�<��
zT!]{H��cT�G�X��}��v�~�z�N����Tm�R��|yZ�_]�cT��!�����wC6� �[�S��?d�`yύ��5�������9���}�\��WF*��^N/��le|���^]���1/�Hӊ�}NO��A`� �=�U�����]cm����:;GR�n�����m�����"�XB��$= �@U�K#>w��Xd�G��H����3�%0�!��|
n*%I��ı�{o��~+L�F���B�����[���ĄW^Î{�0AU��+�K�o��WGw��C#��ߚ��>}�q�,�SMR��f��qRc�L�B��F.g&o�
��]\ԝ����Տ�2��U��+m Q�9�[1UV�7}S:}�ƴ�M������$=E�\(�qŖf45-�E��#�a���k��$�j\,�����2Ȧxʍ̦��������zc�\�����ݗaຽ�+`����)�l�%����_�*��e�T_�(������(�����W~]�H	J��e��1&a+�_Vx����} l����#U�G))=�i�9K]yE8>2)[�o��)2R����B�����pOy���ǡ=�>s���2��)�БA�����J�|I���Y��F=�˾������E~<���V.܈S>��*r�;��DA�j�I
��5��J�DT��S�k���՞��L,�gGOɪ��vZtE�*�%��-a�1��
��X�-�ᓜ0�p�h1�@�;�
�A@40%����/�� ;N�˦r(��E�!�M`5�Ơ��(f3)�6�h.-Z!��MSڋ�5&Y�Љ�4CEoy5X�7���o����c��ͺ�^�c8��<�_�tJx�3�%EWR��Y\�md1峥x���7Jڂ$��ųs<��lS?'�_� Ŋ֋w�'�D�~��Y=lې�!m�����o���
�NA�S!��J$ B�fD�,/�4��q+���<2��if�����Y�{�pvʐ8/#AդK=ڤo�~�[t2�7�-���"M$nOE�g��D�a�8_t���q8�q�7N�Sc_���o��e>�<(�Y�-�K�b5���aN3J(�U֦����P?|��6fbn$B=ڍn:)�r�֏��,A��l�Nڣr.-�V8�p�g[�,8e�#0Z�dȃ�$���!RN< ����K�@��{/�v(i���J�BB��c�FUh����lE.9��c�e@�z3�b�t�_���N��T�Uv�Y�
�/x�s�l�h�t^̊�@S�l��1J7���)�n�*�|�x)U���i�\-y��8�����S�t� ��,y�c�[E,����iZ^\V�<�m���-߮50(�Ѯ���������]m��CE��w�,cs�қ�[JU�O�,7���s+�!;��R��Ȁ7u:�:7.��@r'Y:n��#�.Q_n�����c��dj�X%op���f�y1]�|Ƒ���Yy�t0�^�� ����E�E̢\�JԚgz��,K���,��	�9�nQe�L>�4�wa�gѷ��&��;��;�V�GV�����p>�����N:uLNR�4rnxC�9�UUp�C�4�L��x`�{����k��vx����2SR�����$�:B����X9��9|0eƽ��f#}3M�4��__��V�J�hص�;Q�4��Sfc�ͶCVz���������Q8���
���,�0������w[��k/�s�h��K��O�G!�nL�6O�o����΋� Z�ruY�0�Zn3��V,Y�Ӧ�A@�{���f+\��ߠ�����b��d���	0�����F������ڑ�}�49d�`�7�[o��N=��4Ͻ�6�&CR<fB���B^�{t�S�X�o,�g�T����U����JNy�mi�%4I��bmy���;#���'U=t�Lv��Ӆ��[�'ݧ>i�K��%a���f{E��G��gm��+��b�� �2�%[�s���2��P�]�4�20�\X�{k�}I�/�?d�1/VEV���~�鵽M�]����t;�&gn{��J�S\�}w������Ϩ�.�e0ʆ���f����L�e����;Ҩ���b�0�}&�Ꮈ�%����pA��J���~�X��TfF}ю��wտotc����J'��Q c�ʢ�1���3}*��y3�`)b���TT����$�I��8���^���}34!�	�����3�	�r�h�(���A-X���6a�)�R�@�S����~��(��G�@��� ���0f�S�����E��^&�A����m���+0e�bx��XK�A]�=�[�^�9#���ԣ��g�m�_��n�������;n��o��^pΤ��7�������M�fe��^��t�F��K/Qvo<�F�b?�g`�ܥXI7���w`ꊰ���>.��k�Vx�f )@���g/WJG��Z�l�.�_m�����I�e��p���(�}ɒ�X�x/~���K�M��8Z���S�����G�-����F��a�9�?#m�΄�;�Ò'T.O����m���Kay�&��Ә�,l�ۭ�:�߉~��m;��V{����3N�lF��lؙº�W�^�ȁ	�N�$#Q���`��^6�L���w��)�la�ڭ��|��"p�z��b`c�b3�Nĺ�fa�M6Ġ���o�iZ�h�dr(:�/^�9�b���xy��j
a�����H�&]�1Iu�o��EB_/��6<boɐ���O�~�5�C���c��c���(������1z�h4�J#cq_R� ���������	Ϯ�;�tW؅.�:��y�I8�����&��R=�XO�1��0�{�q4�u(iQ�N�Y�����Y8���p�Y�Ŷ��;֙�}��<�z�I����p�g�C{�g>���}��Um J��d7�D1�'ΗH�އ��ʦ�2W���>��[3o�<�����x���ī�%�_6���8�;�D�ʓKϨ�`.����B�n��XE�O��������s&q���e<�m�;/�Q^d��ԁȃ���:�Q�f5	U ���wpxh �Mm$0�������2)�>F��JA��>�k�wY�M:^�*�C�^��v�Y��McZ3^�O����+:>�V`�����.���L-_���1�]�bfΜ�e+W�o�>��fh]/���|i��@�$�Ҽ�.X����l���&I���5hN��BS��2OS�c�V�	����{�T�P]h&r�I{�-u1�q�>�#g*Px�G<�����ƿ��D��B�N���C�y��>]W�L[p0~�L�l	�	aK�Y�
%W�,G4��#*��p�-���v�m�׭�e�F�����n	#w��%����1c��1��CSԕH��ioV��#���z"�AA*���I�ƋsndZ�k8�J��*�)
7����g��u��'T���������ď�z�GV���<�����S�6H��ݑ�}n����}�PQ嶱�Pv�܌�{~��w�i��}Gu�R����dπ�V�0Н���U�q�+{�|9<��+	z}�!nI~�ANg������U��T�Ҿ��4�"���!�[���}7�s]e���4�Թ�ZJ���Ad���{ 9��J�T��I�`�ss�Hɒ�,*X�(+ۖm�^y������W^K�J�"-Y�JT � �f0 	 @�<��������{�{z�T�LOwWիW/����R͎b\�-�����Hf}p���!��~�	������Uj=t���:ق~3�2@L}����i�5�A�dob�{�K[f1�e�P"�G�H��'����ެ	��#�@y����O8�80*�2���� ����!�"�o�o'�x�T�[��<�쳘1}�����ƒ�P������+�Q-��K�P��in�'�6ܘ�u������+�Ղ�s|�^�QQCD
�^�-w��x���1kf7NX8�p5g�Ui}�����A_���5��z�Iy�@���?H����l�V<�t�2��p�,�Vb��h����/$�����Hc-�Eġ
*f�N���%`=���lI�(��1��,�A5���ۋ%�͂3�B��8���1k֬�����O<Gu���u�6s�l���D���׻�9w�q�2�P�x6�l܆�5.���-����f���Hs'z>�%�Y�	����8%}�\�"ő0�-Y���9��ħJt<�o�y�u�mVΒ�{h�;����l�`@�
�Kʊ]�����]�,ty�z�U��gpYE.5� Lb����;[�,z&	}���ni͓����-���d,�en>'z���U�U_�T�+T�2[,�$�#����: d�3����wHX'�0��d)�2�ҥ����Z Q�Z�NG��✂�����ۮ�%1�g����zoI�@�z�n.�V&HDY�x޼y3����)�����{��t2;�0�p��9sf������bƢVXelz4U�f�K�3����d\4&"�etQ���,K���
m�|�5U=�u��b	�d��	��dp�+u���x��I��*I��;Ͼ����4��>U�Jp��1�\v�^8R�$27�uVJL���Y��1��uUo҇d)c��)6�6��gI�^>�9&�Ah�� �<�L̙3G,ֵ��M����d�����w��p�Ϯ��iӐg��W@i������'�JzQ�QeZ* �� i�C�5�}��UF�蹴p���%̙1|ڍ�7cݦ����%��/q�g�J��U�`��>̚2I�I'Q��,t�غ} ���(��^��{mY%��eZ.8�� ��D�A��w ����u�U�2�-�P�����+jg��i��q�T�5wԇ75 �ƌtv�Io@9l�����X�u��lq��j-ʬ0����G^-��|/�� �)��r���f���ʱ�m�y�=�-�he^�6�?��ua=G��Zӕ�l)Ÿ�����R<]�aj�y\�W�~fvH�ti�XJ:x��U�DQQ�wB��㘷�[{���!�C�
C[Dylٲ�~��%����0��g4��N���������[���#�z��~�lo�����i�)Гb�YcY�ήi��z j�))�^�������S�� ����۷�����y,����m%�ʒA4]fY�<�k6yl)�}q-|�\�����-'c%Y� �x�߱�p�&K�e�ibnQ5V���%��7�����ٍ��Ҿ�>̟7_@��Jx���ʖ(g�~�-[*n/��jc;0����<PЪ[���\��&&�sG��v�x�i���2Kk�/�@y	%�Gu<�t�Q��ښ���ch������+��ekh���<��>ʥ2f�[��\p��0]'��$?��?�4]�ў;M�j�b
-���K|i�����w`�M��+�h'�7I�q�ޏ���%\|��pye�,غ*%z�ꍸ�w���ͤ�8t����;��sp�T�Ӷ�I"�T��wD�P���N"��$�u����\t�����Q&�^�v^�|}�A�-�D��+z3e��v~�q8�c�×�s�������S/�"�7c�j:6$:^�7�s>fR�=�D�i�\���_�������X\#)E�x�͌9ꬲ�O4}���g�)�	�������E?m�̝;�CC2��f(�7תB�(cI���t�iR9P>�`�V�v)0����d�hRqA���5:ߔ$���Ď�*��d�V���~�r��8z���Dt�**v�@��ފbO&%k���K^؈ǟ{;�8"�O�ӈY�N�|�G0��׉���A�բ�����0��˨D�f��2�;q��3M!_�FN�{v�I��dA��c���ϵ�$o�k�E.c���r��mx׻�)ڸ��l��p�B<��c�2��E3����s5���{�I~�J���Q�i�O��o�(���9�h���m@10n@�s�׉��y:��b7m�r��2w4��\�ע��D�rg����:F/��Q�+��DGs�]*Jw<W�L��
��Ȭ ���W�э�5Ԓ�`��Ze�+.aV�=�͗�$�D��,�1��r�+��#0�@��m�?�ѹ�.j�O?�ك��x6��B]�dd�U�,:V�]�qj�ca��!H��+��²u8�#!�]�8M��.���>���*�9��S��M�Y�9����)�d�ԯ���p*��h���+�_p���#ɸNlFǲR[[Ƚk(#qU�2f:;]��w�4�������K/UF�n����i@z�y��?����GK�X��'�i�S�guՔ0�}��k>n��kNrZU,
�h�qҍm�*?�
�>�2�̜��f�ٽڭ��� ���a^]��m܉-a7}�#YX,��#�O&j��,��VDeT�0�Ƚ��4 �N���ق�n��`�Ne�i(�C�.c��8Iҍw�R�2�n�h����S}
�sQRm��+���}d�"E..�����I���-eom;�� �*5��F����WՕ��2}�>�z��2����e����iL�:�NC���@<�V���-�8�� [�����@'#,����d��l}Oʪ�*��V����铲T�T�cM�\L�JF2����$j�٥���YmwCF_�a��Eױ���J�F!:�3�N����-��O���v
�|!�Ta�M��q!5Kō
�i��\Y��f��*��^.nz�5��	���趙�BO���G��	/|�pɒ7�G̝3k֬��
���x�3e�{F{��I���;Ui=��a��#��#O���k���L���
�N�����#F^���e��=V�G���|�\�sYM=�9F*�Y6YKc�'�<�
i�R��*���(�9wuuK���7��E���
�G!��U��X�{t�F��ĔO�8�s?�y�Nfa̅j����N�ܾ��c��|�t�&O@�8/WiY�u���8�s��#���(졅�*�P ��jH�6��1݉�Y�eCC�{�^�q�ql��82fi|�yq4���P������߯�ť�
}!9�9A���9n�q�WcX�N��!�(£��b���e�g�=滅;�%T,��J�c��f���D�3T]CY��Z�ɫ���V����'ךE�r���\�S9�P�P�ɨQa<�q�Ի��Ǒd��|v�\w���E����m3�'Zڹ=��<�G��X�1�6M�p�n۶m�ǳAahhH�[\�E�R!�@&�5�L;�3\{,�86���Ǌ��{�
f��`��x�U�D��C��BZ�  ���D_�-4��ԏ�$�c8-�Ԡ
f�O�^Y���F�3�N)�?i���gI<���)v�Z
D.�&��t
~ލ� �# ��H
O��XM�\`4����PaXM�C��G�}n��s\Q ��UƤ �����_s�̗��Q�@Z�B+�\1��SO��mٺU¥�S��M���P �ٔV�����~,+��*^�t�:X�Emq��+��'�rxS�������,O�kR!��r���
�x�
72b�v٩E�-V�H0��8}\�EԱ\Դ5l,�NU:r��,�^���%��֘����"�|)����LhϦ;g,1�:��	EQ\W����U�����A3�<���aE*.�ҕ[0z`��1�A�
T<�!?DJ�X$����^��9)C��cƤ#�dwoc�٢i��h-֬�0��'B���2�����.7$D�j<��X[���/d��	�O'N�'O�=��#�!�}�/,}p�,|{5���+h���Q�=��f[�x�c*#;����5�36𣶳�[�5B���f�PE͆(%A
���kvc��4��֯[7���N	M� 3�7���=��7�E%�ց��f~�N����{' �e�VXC[�S��ƔE�.U�#� KjxS-U�R���6m�$|��"8���`�{g�
���G9n��UJ�qYDق�m�Vz1(�����
m�T��Y���)a���@��� ��� 6U�?�0�9=r]���Q�[.���㏏�*z뭷���Gek0
��Ҋ>�=�^{iƤ4Zi�jȉ���M�ij��6'��ƁK��4N�RL{FO�R�?�֗]��7���{CP�~.��n(�U2���;$�h����h��s���-�V���y�QL�:U���j5������my0�E�]�M�2��c�0��3Տ����*��T��z����.��w>0B�#eʕ��30:|���HrP�hS
�H^���i���4rd�$x}��Q���I}�' �c�K�+}5RTLeNּ�:�j.�i�=�N7G��� ����0�8����y��g�wO�oK�}� <oV��B@�T��6("���0z᱕�ݲyvm�����b9-�\�F�i�y��5D��O�QeZjE2�|k�%��^������.urtFx�4<Mn���mu@��Z��w[�m�lM4U�K����-Ĕ�I����t����X�BȻ�����c��/d�SjVՎ��S���$f���)�o}�d��N2��:��Q2^���If���߼��٭dwfc!�[J
�J��u�KiH�ٝ����s���y���gg���;B���u�>s�X*آ�B[��L�1
��ju����}�i��?J�x���e���0ښ6����o�U�cK�5�M�Q��J^N������%J��ua6�$������� a&F>@���W�꾟`��q9��j w�{��@��0r;��=ì�[�5l���}}���7⒋�,��|)+kK�k$J�����#��w�H��dϹ6�ٶ)�����{�~a+��nyj�9�2�oL�R!���bf�ط��n����2e
.�����Y@�����Oa�K1c��+%�#�����[d¨&�m~z����]�kn)Q��a��V�^��?���b�k�'�j�fx�������������JQ&�`���=��Ѷ�#���$Ja�G�7KũǄ���}�ݲ�^x��y>4�A(3"�r�-�b"|T�xϝ�t.N�yv�u��U��P��X*DG-�w�5T���4�H\W8��qS �B&Tx�2<��������X^Ϝ1��L��m۱u�6��܉���oR�зw��B���MT����Ͽ�$��ˣْ5��(�����Di7��o�1l����R�0|�ુh�2���џ^�ѝn.#,*��ñ�@�rѧ1&b���[�$���'I��!�97&�@�ɣF{zz���~�3Y�9��|�l'l<`o��
��a_Sq��[d�$�v�RX�syb�L�P�3�*�)������S#R+iV�e�L���7��@jH�y�[�n�����@�HJF�v��} ����9�崸�X�x�n���8�@�]R��U"�|��3��W�)-��9�\%w�f��n�8�%�j��kע�c�k�qJhN�Ժ؁���k$�R"x�JhA���f%)Q�L��Ś�p��c�y�f�CY�8�%�^>;�C�t�6���_'q�X��3���Y�L�y���&c�঱��$�,��IR�ؒ�$&�R�t�uU�5v�j�yZ�����K�g�>�d��na�)J`�澾,^Xh�f�}+����}BL�:S�����JZ'�}e�%�*�>�;�g�b��^̡>����;�n�vl����v�OC�ǥ�|/��@1V�n���m
�2�Ҹ�[�wA�Q����xc�⠁Y�A7��(��b�,�1�3��\yd�^�M^7�����,�KZ�Yp0����Z�8�g��B��L��y?�q{�A�,q}��ʄ]�S+^W��trR��QP��y��PV�����%��2����L箉u�bŎ��&�qp�d�l5+	�+[�fM��Y�ʭ�ɧC�	��ڋ��I�,�*�q��PJ����mS4K�J����M-�,�N�,q�t��(fA6-]�ъ��<��\Ov�?��d�!ژ��ҽҪ]Ⱦ-�b�엜��d���	N<�0,:� L�+�\�dM�~s*,WŜ�W�!��Z�8��/���~��+a����u)O_v��@��������	����d�൳�6����v��&r�B���S)+�<�Q�sv3��~cŀ�]�/3HakQ#�����o�S�o@4���Q�䐭sD��:�1�1{l%��0ŎؽU# �q �kR-jl�?|�
[@_�,�c�Cl_���vZ��\����^̘ܕ�D1=T����R��.?�2j��6m�j�E�1Lli�1c:�<�!�R@��玞[�*��&cF�Y�N����c�eͳp�|l� ���Q��"n7�t�օ��; p9�q$&�I����i�釹X�+��I����v�8���8y�L���3X�	`}ׄ�D�Ċ�P����}c�1W��_�b֯?f<Y�t.��)�G�`ϗ�Y+�	S���J�,���z�C�!1���B�A�ntsO����� O�k���Ņ��sb�P���b�����vty`i�PYYʍ�rtр�!Ԁ]�2;,'�G!E7���N�wK�&�))��%��d�#t�.��*�I��w,D�6	���V�l�p�BlW�cE#��S�#�c���ps
;B���>5�i��^t�r��?�+�Z�O�f̱�'�0�T���R��X��HY�m�L�48��il.q
���PO�lܷ�S���qi6��dy��=R�'	��C�8�#p������UDC\��T�L*���z"]���)����U����-���^ـ�5�^�XP;QƚZDe@[풜����g!���:�N7YE�"�gV�_�cx�jC�F�֚DJӎ}U��M��b�*Q��X ���FJݐ�]��b�;w$��W�Ǣ@����4���-$P{��_~�h�4%�%�s̶�}�s�)蓹�_s��ZKZ�k�҉QI��u��q�j׋*�G))�MZa����T�C����Y'�O�y8�@�K*!�c51<��3Z☶� 㑔Yig��I�! 
���t�Ϋ��֩N�C�y������#w�}������f��������WA�h#�x-SR�KI��I����B�2��m`��@�U��v`����?�5}���a��\�\Y������jI�ҡ���&e>#]2��,�:p���m�N�*�~��2������<O#�o����1I�j�3�q' e�v����^.����S+-��kL�E�K�`ʼ�ǌ�Ը��5CNK�I��8N�3�3#���yBv�ѓ��y����C��?�N\����/��84��m�CJ-)���b=�fp(@�RVq��ݒ���|��g�-��9�{p�OQ���$7&[�s�p�g�sX��� j�D��	�l�&p�uT�?�=��N�\\I�,��ι��=Y82D�{���T�XM�86���<�z�;q�3K	h��X�E#�;��Y�n��>�,����D��Y���x��߆
ϭ�yڼ���x�'m�QT�ER��I�����%���g?M�( ��:�Hcm͏)�o��?�\���=���̶;��jh �d?�z&�,E���F��-�N$ڏ��7:�IX�����f���3:���8����������b�<^��O�A�|��5��Ս����ɶG7�$��4�<D�ꂢ��?�F�͙-Z@�7�5[ݚ{oR�v����%�&	Tw�c���+�)�M_梇0�%Y2]T�D�,�G�����zz*��|�\l"+DLX�yY�;|6�m?��}V�O�[��Np�h�5�	�6ހn~���7R�޼��!�y���ҩ2���Ǽ��XH�/
[�,+ӷ����twHR��N0hHf�lmHr�%�Č�K�~���mW^�]-�Z�����gM���_��=�Zd�� �Ф7�,[I]V����Oary���n�F�ZD�i�Ʃɰ��d/����[�&��L�KI���P���|�R V���9�Pǌ%s~ym)먛�*�#1�|��e��!QV^˄W$�r��ND�C��,zct&L�t̍m����7��m۶m۶m۶�|���w��9�g�f���9*͵(�6�w{H�>� �(}e�
��#���x|�fD�����:H^�2A�'���X���:��ohB�d6X>1�W���No����ZWd�2#RG^�
���6ӹU�<tW��	k0����{Hj�4��ވr���5�ziѴعw&����1D ���� .c��U�ɓ=qϞ=q@�� Ph2w!�1r�l�w�4�͌��#U�GiB��	����t��"��B�\���
@،��@��nF��[�)w��|�`3:�]WV�2����7�\�[�ZA0]ی�`,5L95���`׻y֨ǱH�h2�D�����֭O�R��k��xk����Ln~@mh8F�ݬ�~���D2�϶��&�(�F�B#+��������q|��Gݺ%3z�=�,޺�?�}	�m�Q�NЋ7��K&0�
���Ao*&۰o��ฏO������#� �i9�����D[Gek8��XyUd�a���<�[����^E^%�c����#D�D?>w�i�o��'�5X���=�i��E���zLa�̞��ŭH�x�%,Azb�yS�k��Ɂ�V�f�v�˶����@���o��f|-�� ��#G4�^��fY��t�x�A#߹F�j�aT��/�^�7�;Lin���毹��b>���mZ�G���[��p�Q��ӓޯk�s/��7!5ю-,G�!�GaK%��;q{�E�1x֠����K�г��>�Dj�i�'CǶ����| ���.k�n�g ޯ5���z�W:�D��j��g�^�}�l�>[�&��ďa���
��b&�屈�u+I�7��rWI�S��[���pB�4E�L��;��7�Z\L���[V�+&���Uk*��p$�\��:���Q�I���
N�v	Z ���h� 1�>�ԹU�v$7 I8]2�&m|$�k��f Q��u��j:�Pe��>�-#T��@__�d����	iZ����20���ڔ��Ϛ;T���-�K>S^���950Ó��y�d)g�v�$���f"���,O���lv�U?�9D�V�\z�?� ��= �S���o(Ե�Z�C_�Y��xjO&"���.��&��u`� �X1iw��$+�P6<�b�s��������O�����#.�:�?%1�3�G�lr��]a�z��>�D�uڲj�v
P��G�������D�Je����2\�v�&ԓK)��A�0��;H��9}?d?�Ѭʟ��T}O�������2L���u+����3�>��dEg���D��k�=�=��h#����M�7�2����j�(�r=j������r���~bp$��;�lWm�F3R�*��TB^�#���C���w@0���a^���n-�e�ƺ*?i�������M�B�1ht��J�5T%dVu/��
��+��Ⱦ�-��;S��8�H3��+P�4 �2�z�_z���^�@��jg�qq��ޝ�c��{̶�k�]ˊ��<�i�*f%�r��w��t_'��Z[��]E,�a���}���)}Bhm�+�I�'�4�[αcC>�e�\��4�[Tf�M�CP��p�6�����oJ a����G�>�Z��!#5���fJR:��uyvR��t��b��,���4ڗM]��6�5�4.T4�����D�'�"�M�[��7��ŧ�w^�S3�D� �\r�a�rF�=��%u�������l��`sL#V�� X�R8�f�a#"�#
Y�1G%�F����g+���/�jR�J�+�}t�� ^iM�̟�:��k��ZK��3������������0����ّ.h.l*-�Ă�H$Ʊ��L�����������eb����z��~���ca��f�<$_	�d:M�)X��=�y�F��u+*2����O�[��Z�s���K�h�GU�V�;��|l���o��V=i�?7&���nR�:)UjtK�Z���bj�v��w-��<�S�$d	�(�~�#fW��d�aS�|ߕ���j\a\`W76����7�^F�Q�l��Y��M	q�]�WXF1�tk���c���=��a�|� �_n
�QniN��ʼW��]?h�<-�?{�f��z��>���W����ׁ�Q�j=�������7[T�I� �ɂ��x�q��H]�t�̓�j=k_}J������l�l8���ne���N4�y��-�j1~��~� KE�F��ڮ++�?>m�R�6�C�W�yooZtެ=������X���p6 �>�A�ܿ~�5l��±%0�w���0H�����?��=P�%ZiW��[`W-fowN�M�'��{���nR�Rُ�6_ɔ��E2*</�	Y�q<���Ԅ�s⡄�ΊjB�FcD."3������E�y��\�ưo{�x��YX�����
�"�.���0�i����^5�d���+�_.ĞmG�CU2���t8E�H\I�B+�҇��$�S�7���6��\�]��z�*V,�{�P�{K����DҘi�?�6;�٬֢�5ً�ri�����sP1ȭ�[\�Y�/���CG�5�#��TH/�hؗ��lU,�L:8vnyv!S�s��Lz8�]h�o�k�g��{K��<�����9��[����qi��k=q��K]��:�]�;ɣ5�䪄HO���N�k5;���' ��1):�e�all�����ʓ}���((�1��b�dj���(�nwh�����ӽL�*�;��A�'�����H��T����8�l2a��&'K�U��av�]*�:� ��8bD��D���Χꏻ��P���֟�>��P$���|b����	.��g3Z�=�DZ�����F�c��{�-~�_}�%m ����i�������}v��F�#|��&��������"<d���2t�/�γG������S�U�$�Z��u9��ւ<a�����`�"�T�Đ[PUm8M�R���{��+��=n�4�8X!�������W���cI[b��طS�{3��^�9O]S`!7dѳ�WeM r��K���pX�>$H)�}����I3�K�:Z���03Za���ԙ�\���5=���}��H���@$nT��v�Z[�=v{|��=�D����r�RG���Su��r��K��: [�bNm�T��c�i�I���9���Y�D|�3�SF��ʙ8m�Ѷ"��)���n^/-r�f:!��������MM^���WmAZ��׋P�B��x�&����rmcO�L�[�<N<D��#��=���Rƙ��]���B�n�)�!C�#-iR��>2���uoIbݸت�;�?& kI�cq!��`��N�j����s�>�J-<Wl��"� 57��`"���A�	���R|�8��"׭�)J(�CT�?UB��b���r��	��mv��>q���NR���R�?(�GR�6Q��ةd�!��R�߱�@Sq���;�D-�r����[�'�_⨧h�5BU��m㗌���F�ϫ�#�wD�V?N;0���缷!B�[&�z��ؑQL5��\~-��ĬRg�7�^��G�v��ʴ��S��eN���/�k:���m7=Vj�L&�M�������e��O�( z'���s�������j�>	�`�^'��p�BZ/���sc�b�E'��&���ľԴ��l�|��N%�}�ءx8a�1SI�8���qA�k��N��A�:�/���`����S,�_U[��Faѱ���4H�[b��S�/�"[P(�A�ﮏ��Uu���f�'�ap(�m}��Y�����=�V�/�[�q��#spِ�3W��.0��NK�>�Tz��_S��u���eK[�$� C&ǟfǑֺ���)*b5�
>�M�5��[	��-��x|I,U&|�/��p��ު�Y�=�6C��$o��.I�e���(@�9��!�ݤz`�T#he�n��|����X�8k��M]�IUNm���B�A��/���d~g�	Ю�G�Uy�n$n�t֠�$��}׾,�Ɛ#B.�Ĕ��wb��`f!IE�<x�6h�g��ʒ&6�Ì�mv��)�es�����.������L+���C5��iku�B�D�˘�p��
+�/�4¢�a=!�'	8���|4��6��]�acP��8�UO��1O�ؒ.$�
��"��x��$˜�z��JA��ƌ�Jq��������y�,[�Z����H���D��$��r��9j��9���CƇ�c�?�Kn�������h��SN��N��vs����-�KT\r��	^Y���ް���A��WA���j���vU�v8M�;�t�!��߉��~^ u���@ZI�?���ۊ�j���o�au�}�|Ќ�)]��׭}��**��������aV�������,����KWǹ�ׅ�/����_�޿�f}����D*��z^T�T�ɷ`���]3C��@{���#�`���kxS1�6!�$J$;&@���&%�Q��f'��S������62�?�̮���~�o�����wP��P�2�7�̮�֤�a{%�u�P�x¬��Lz߲���*�M�j�y���Ī�����tu#�|/Ր�j]��l���ⳀJ�X�կ|���&A�d���&S�@����AtӒ'I�6��At�"΄)V:���Z�����W^�C>x)`h����� ��� R/Ǫ�l����{�l��ʟKT�x�KY�M�%Z2匲��q t�����r�`N\/ o��&��[��� L��u\��,��,O�8����$��͖��7Ĉ�Lyr]��D&���?CԮɸ��L#�5�p��}�']��\��A�� @�+R������]6=+Z���ݎ�0&�V�zx�˹P�;⃷��頡^�̛�fxq�pj~���o�~�c�ao�iI�-�����VVe*�|Me�)c2F=�1e��?��AR�0,�
9|-C���fr<�|M�+墒M7�p�!%���9D�{�%�c�L/'A[j۾������RЗ+Öd١Os� wi��RP�����L���6]v�\_���4���D�����)Mz̈Tv>��/��3<R��W��{] �T�lx	r��Ag�X����=x*5��=p;��`�D�l��ڭ�L��M*��)5����A>o�=OW�����ӝ�o�J��[�Iԯ3>?��Z��m�7����؄��IK��[�Q��S��u���pp�U�W0T��<"��)@���(zS5{q�컋���[zr #WA䀓ʂ��`8�׳$�߳K!$�䮻�Č��U���n����z�Z�x.?<�,��f�S�8����" ����`�²�TTh}�m��zc���p�=5p�N梜��w8GbhL��BE�QF5�R&j�m	�6��2��eĔ����m)��3��i��������m)z�vQ[��K������Q'+�b4��V�w&��jYU���=�K7�i�
�G>'SY�~�d�&�r ��z���CYEl��W��D����<΂�@�ޖ["t�໿.�!q������*e{��<κ��o�[�k����Ť�=�Y�wн%2�0�6t�ۋf�ň�����L]@mG�cL��0�M6y�e��LH �������6Aύqӊ��A!�]��8v}�~'e��Et7������K�GW�;ܗ_�u�	�T��C�1Ȃu����8,V
���Fex�����j}$���%�$̂7��r�Qވ<f�8k��3�.��z˂sr�J�7���n�Q��=��:�f��5h��aj���oΆ��*� �y^��RW�����Hv�I�;6{M"��r�_���9�ɡ�4:�@�u0#|B������~���>o!=#�=��HZg}�nv��$wy���`��4���I����ۭh����M�� �u����]�V���p�\ٿ?���[|ny,#JHj=���MR�C;��T���7z�m>�J�1�������(���q������3K���L�$أ�(����$f�9A�LTٹ�<g���%W����_�:A���L���V�q;*2�S�~�bu!�n�.��
a�yöQUۙ3��`�O@+[�#h��zQpܢ�ֆ�Z~�pvxi��+�;������w[#��2IB���*�� ��V�ZX~�Œ ~P@�T�|/��b�z^<MEB1�ʧmpB>g��~I2u>I[RM�6��ݮ�I�#�,�Se�2^���d��+�!_@���
��z#[ɣ����/��R��N08�mV!��+ a7B����I�	R��8�+�}V�y�6��̞�c��e�����=gn7�b>?�ʂ}�h�m7x�&�޿c���x'�&�s�$���E��8;�.�����w��߃<����)D�\�����p�v#����F�O�T �þභM�͹hit�!w꛴r�k�7 ��}��6"N��-uP��Q-���d}g?��K5���0��	�ZA�D�u�P��Nngv1��yahu
�yPo�Oi;?�+7Z�n�t���<��'��٢����28�0$Rڧ���ID^��Np#�{���y)��3��B3
i�F
��n%��^�G2��ZSR����T��6�ەY����ˉ#�K�	��w�J4.A%�0�������h�P�G^��ir��js�
��S ��������Ŧ�";Bm-`���`���J�G�l�#~���@I��B��2�Z/B���V�ף�ˬ�ܟ�IS�PY�P�"aJ�a���0LW�dd�T�'�j!߄��ֆ@2V_/9�0����9m���s!|�?g
v�7q��exam�~�v|*��O���y���|���(x�<ɑ�f���A�2��x��⠭���-�;[D�+���)��kkz_�F���a����*cI�o1��f�^c­�w�}i&�U�|�g��oR��l2^��v�Bu<�\w�3�(����թPdګE�uԾ���Y�;n�?�����6��F儐!��G~,p�i���8(��Ҏ&T���=���:"���t��|���� >�C�4�N����r�|��"@7�&�W�:]�'�K[�<�Ydc�
���
|�Ȝk����d3�L�ep?u���6�p��,+����[�kK�s�Ũ���7�۠EO��c�$�4f#�w���e�@ײە≌�������Y�8d�ƯL�5��]1L�˪��vqH[]�{�-���M�}�Ҳ��(
��C��
ക Ѫ�Uv}�A�������#x�o�~�?�>������	8ǌ��Rዒ�~��x��Fb�b�97�f����:����E����bR���2��zˇ�����D��G����=H��
�/V�7���u�����}I7��;mh6?��	!�^�]ry�A-ǈ��I|d���TTsC�xO�~���%C�P�i�K�f��_Ċp���X�]9{&G�=��D�^k�{��ۆS	�˪66�kj*$��㛘���Ef�v�S�@������{xx�Ӽ�9���z�����]<G�%�_��x���իm~�3���Ь(xH�cn�wݬ�'[{�gL���`ɕoWs�+ٓi�Xp/�8_O���D��Ԥ��i۸�ԥ�*��^��QrXC�Ǽ�ج�I�#c�.c��1>�nu�����]�NC�3n��ZO�=�t�#빰@�HF��ؾzѕ�����9p��4�^;��Y/�?N��-�|$#2e��@�>���/��{ى�rFX�i��IV�;�ݫ��}����E�u��.B�"��P�
�팆X���SD�Ju-$�ƒ&��e��s\��h�T�t�*=;g��*�u;�T7�4"�"��G�Oun[[�*G"�.Tv7��ʪE��H���t��2��G�MG�\��Gs��|tٵ���.=��"W$�^<�����Ѳ^�<��[u�綑Z��_��\y��ɼϳ��g/��%���o�ݯ1��S-[QI��&ymye����wY=1���a���-|=�'�<��_�|�?�h��-.OV�����n��R��Y����o�M��Ej#%�`&
{�8���j኎�+7�)\�ƨ��M�%��c8����o�����<6.)>�w~¤�U�������%��9yg��z���Rx���$e�Z��u�;�H96�{����F���b~¼z�j��1i�
�=J�+�J������l��#�?�ͩ�s�I�(Ɵ��3�˲�e�)kҎ��@vk�Y�c���������_&� ��,��3�~ƻ��YQ|��vO#�`4+O�*öNY�]��8�T\W�E�4V&����{�9������f^�G.>4�!'�i��ܶ6�G�5�|v�߯>��^-����AR���Q�����A��r�O�(�هK�-O�c�,Z��u��G$ﷅ���#d�+G9*ߑAV�o�L��W[ˣ�0+����U^9ET=��ζ��'/��;���+��G���E4C �4���?�#��u�s����N��
a�:��/fc��~��<�R�Za;q���bΠ�ϗ���.�Ͻ�k�������k�Wv!Zo�  ��D����'��s�g?��xW���u0�'-08���i�&��v���RQ�����m����|�-7Nr7��7��[2)M�������<�_��G��\Q(��S{�ؿ�[\��N����j���Fd�n���n�	Ȓ��kC��e�ק�ҩ��4�*��ЩF���Uy׋��^���������i#ʙ_��{^Q�QjY�ϫk��(���T�W7��d��_}:U,qq�F�m5~���@��z�B[��9����9�}S���yYy�ᅮ�H���B(C�{������k0���f��ԃs��0��F潫�~Z����|��P	�9��,N`�����A����[���=šc�Y�z�į&���������?
o ZKr���	�c��*&\�~�2���Ư��c�Up����1�^xm�P"�{��u��w8S��3\����"<[
A<Тܟ����A/��G�w���()Y���FF_�^6�Ȟ��H��K$9���gp=x|?kOju�tr�k
}�|��Z�wo���;1љ	��Nv+[=6֭�3���e��z�����Y�n`�(k�"��2�/wmJ��ES��G_���E\���4ӳ�'��m�j��s����%�NrZAiC��|#��so;�R��&$پ�B��%�z�z�q�4�f�JFz�H^jD�~�l��&Ή��0�*NJ������SO m�Oo�=D����B��W(���@�k-[Vp��a��S�#K�����w���0����`¢)6 �nk�!M�Z%������t;�r�{,W��5>@�B�r~�(LM�|̵x���؍xŐ��,:�3�o����|�F���*&���+42�M�|s����K�h��6��Y���r�1��SG�ܶJw�܅��;��΅��Ԋ��:+��c�%�z$��!�r�4qM��PS���"�������y9�D����-�c݅�i_�I�VN֭��gL�KI71n �S'<O�r[�u3P���.��� j2Y�[�%���j�߯u
� q<�<:d��2��D����O�x�{<8.@�eߘ���K�n,N�hF^ۋ�_s\U��ʅ���eI�!��`�p?Pg{ᕫ�POU|�s��Je�_e�n�A`/��ru�A�t�ʖ�Ihu�Q�y�]�P��/��gQ�����U������E�;��z�( �^����%$�!��ԩ�d��rx|����i[�R���cX�c|���Hj�R�CRt#���iq�w���M�H��_[���D���XU3�s�|q�[򔓹zv7�ҿ�|�Ƚo�n�%|[��|#��}3�B���a�`��8���ᗑX�w�v�7^�ʣK��X���)[��#��c���J�ZSlN��˳��)���G7���i���$�X��@��I��P�?=J��&{�ʡ��7(Rpyt�9�]U��qcS\M�j�\5.��[g�}���2T���C�H��Fe� eB���xh�GO$�ߚ?����_3Gg�'R_0�<��Ù<�kX(� �ΐ�����L��V/p�9�q&���2���Bv�38V<����sf��I�A�������k����J�$��'��1�u��'����5�Ta4��Aѳ�cX���o"�ȯC��|?�`�Zs��-��Z�M����4�����A�)r���⋮NSV�ʄ����E���_8;A)JvW-��Y\�w��K�L�Kޙ��Я=_ �g
.�u`.*f52��!����$'�i�����:Oޙ��ɔT?�K6Kt�m	A�S%�G7]�!�f�`,�2�/<��󘀫B&hMH�GDF'�$ԿU%������H������P��	�+|�z��"Twnh�]c��+o~I���56�PF�,Z8YR���W�*�]=���-���E����_�tL��X�Wn�s�E��9s�q�\��iQ���Q��װ�n�K�q�5~�$�kT�i2ͷ�,[#X��U�g$�Ú�m}�+�s��ggS��!�bwY��j�?���ؗ\����j�$� ,)?���b�~���ϐ9Nց���"{��Uk�����,~	e���U�f>C�=tFpVg0�yrN���D~��`�����	)&�cLs��-獡	}���:�����@�W��C�s�#'�e�ͺ��3�R=�Z��|������֫�)���}H�v?NM���d��]8�+������B�:a�
m��ů�n�T�p�+�"�"�+�dBC���u�O�Md\c�ةc��t�YlN�p"��"�~P`$���g[.^5탤�W�iDD��4�w���F���.��%O<׆�A�[�!ޓm	���E��1�s$��?��c1b����jZ�cs!2Z����q���k�&�v�|߂ڎ3��kܐ�%٪Km�)
qo�) &չ����b�0h7�kٌ"Sk���$O�hk �Z7!�+#�i�Ս�5\3�t^�䒣B9/�x�#�)������>a���4��SJ�;��m�z��C-�EƎ��0�����������ЂӀm?Pmo�}�.�Or��}s�`7���(��Ox|)R�������|��e�$��B����Z�}��-��(%
Bs�<��	��z�X]��`ZZY
z����J��nwa"��Y<寷J
~�]�"A?ذnC�#�� x���7�֡:�+3l���2�mI�kS�o��u.�8�T0��ģ��`��(�������$�_����Yu��Xp�;s���'''����+�zj��O��U��bɱRL�]��6�$��0�i��7`�5q�)���Y�4I���{(�{��#�1q�X2�����x�<��Z��|��,�CN:U��[��Q���r��l��V]��]dBjkg�W2Ss����Dg~į��O�� x���&[���s�Crz�$'%�O������L��������a)37�YU��/�m��ZhV� q��*7"y�l}z�I#;zu�n���R,����:����+B��o�Ku��.�4��yA����y1��UC���Tx0�.��Y��ꡙ��:-�Z&�3�ɯQ�W�eD��o\�a����2@WgP5�G�!�17KuAnp|	�&2��	�����zq6��[�Ōu���Dh�6v�`a�paᐼ�2���_��·�{���7.�b�u�-�S��zvo��G�-�o�Ӭ��/�va�ɢ��B��d�C[�k�]ߟe� 
��#���B!�y�_Λ�&�l��I�Os�����`���t�t��L�^w�&I	
�yh�eP6���E��N���2��L���$:5|����w"&uC�(�;���>Ф���B���v��W	"�������3bg7�$����v�	��.�Us�T�r��H���t6��`J�v�*"ol��E��K4c"il]��y9����G�;̚����C�d/�o#�k�o�����l珍h���C�ҨB6[+J����r���)�&��捩~8D:�&��o� $�^S�*��z�g$���FI9ul�y�+�ͻYf-�k��;���7UMu� :�b;�$d�b��t�q���b�v@t"P�9�z��nx�9f��$���Kν;j;�U�XE8����^���jB�Ay�X\Dʣ[�=�)�ꫪm�ˤ��*)\�����:�D36Q����7�u���	��D�����|��I"_�yl�z��?bi9.H���[�B�����U|�#j�Ku!����.A��j�A��#� h�po��&��=����[`�����ݖcf�`�9�����X���",�Į���/4���HfU3����.[!��A��@�t��!7����?RC�8�\NP��^E�}1��|���ݭ�&Й����е��� 01���g��v�eu�vwr�_�e���jO�h.<��l׏؊X��MNl��B�ڇ�7p��n�QҚ�ێ+<��o���Xqv�yU\���a���O���kz��_����u�o�|�g=pk����P�
�
VΜY�#J��m�%��]�_�Zw^A�2�`P�N�n��Sڕ�V�Sk�|X�����q���5�!~���Q�c�Π'(��<�ٱ�-V��4�'�EK�����`�a�^�'��b��
��"[8�Ɵ�?b>;�!׽�`� N=Khe�;+���v�,�P��P]~Wk>W�<���\�>��a��;�*�?[	�z=��'trA]�eÖ����%�:������n1W�L�m�_��p)6b��3�gY���.�+��;:R��mkC�2�|��y	�Hw#`M@�\<�~�#U�f� (�����VC���m� ��
��Z�&�̷}��)V��+�g�1
*,&��)�T�����!����q�z�����=���h�pB��D�4�0�p#��#��h��M��{SoJ]~$��;��xI�_eh�X�]&�����q�����z��!$��-����V�񻶍�<��,�����5�xu�$���0��i��H�c�s=�,I��ם��/Fa�e`�� ����Ɵ^�DV%�{�Akhݟݿ&tɀ���,�c,q�o]�����v	eZ�"	�I��#��[��ұ�"ژ������}QU���#,U6 EMו�7�<�L����\����1(S����I��D ^E`Du�6������ ��7.�1n��a�^/(<��AĀJ&������=ͯװY��&�W\{��i�>ӶX5p���sM���IDu䂻�3rL�ٚ�K}0��:��5�^��J;D�;�^�Ϫ��>�DVk���Yi�oKg��Y��o9!�H����T�܂�ɘ�D�<�<U`����S"��A�_3Jz!P�*!�mFB�
1�3�3�yZ����g-'�߃+������v�x�C3)���B	p*�Ԣ�'9L7��`�*�Hg���e%��Ie�PR.Q��2{b���8���+rm�=��A������<�����-�H�ѣs\k����>z�ҬRO?���Ճ������$Ut��-��4�KbɪS#�I�������w4D)PG��0
��e�Ta��A>Q��a_Q�#��D��E�o��5�i���)ͦt�$T���W���(y��`�_"Rc�����	�+���O��bH���m���n��ׂh�����6Y��i�,"L���6����YI�M;��E���LM�D�q�(]m12�������7��1�������Qm�VIk�q���o�bv�O�	�Z�z��y\Z��a�5bO��$�G�)H�0���喳C�R�M-%��p��G��l�{�;k3�z��9�]���sɠ��7OSV����QD j���/m�>���Q�M��8�+�;ƥx0gE�D�L��l��jd ���W04q�O�hD�7��g�0��V�F�Q��	t��b*�l��p`��5�ț�A�(IPF`�:H� l�-�~��C�:��u�b�0~[bTz,j�O���l_d絷��0_���f�R��⤋aj�`NX*C�$!�.��Q�S�%jZ�`P�Ƕ��^�߶�H���T���tZC_rt�x�>�+�Z���BV�m��[��N�ȗǝ3��V��	H8#[ʁڃ.��K�"O_٬�ܒmo�G��$m�<��(�I��P���Mm�?�3�ü.�
��i�v�n�d�
D֧�z$3+P���O�\QS�i�#^ ��V�`����}��.Vg7���ND���{k&Q�� ��
�ݴ��������,��dy1�#А�v��a�'2%p#!G6(N,�F�©����ׅ`Ŏ�1��t�ܟ���=�������4���u���0��˝wc*�0��[
a[���ggy����mn��[����,�����~�t�����!�
\��Lf�-[��5��wzB��+�%+�҈ǴI����-`2�R-���?�d�t0ؤ�U�d�S�!�y����2i���
G��8�L؜ъm��ޢp�.�W� H�
؈���Є,�]�g$jOb�ţ7c�[�k��`�J����p�����ز(��������d�4��G]ԉ�ɨ�6�_^�,���Lꔅ�v������I� "��>!D��ʱZ�(ҍ�EY�����_�y�H�d�8(�G�3!E�R��5DZ��Z�(��Z�NFV��(�L���P���6g�N|����GN�>���+��)j#VO��*��
��C�����ʹ7e���Ƀ���z����0}��
�l�� P+��+���>�?��KqS�ɭ'������̜	��k�#
�*+�j+]��hUo�^@ԈzW�H�W93��_
�lLG����q�p�Tl�'�Q7�o��S�/@&�E�j�b��Ӿp���ݞ�ဗ���Q#���XA�QN�>*�f�.��o�"�N�)���&X� aT�jm.��WT��4Sǽ���F�M[<G	"4��V���OHS���K��[�PH���B���=~+�<m��ZGI��S7�rw'Xh�	�&�<g� X�^�wqP���MB�.���06��m�@�{r\V�d�¿�f�� ��]�@Os̘{���vW�Z�뷄x��������(oҪuDm�;$"�U�pD��t�-������*�Cr8D�_X���O,)��	֟����?1�c���f(�O�z��b4�{�a������uP���)��$qy��A�zO�^���� ���j�72��X��x�2ut��I�r�\����nX��EivonEX�ȁ5��d!���g�_�s�К�g��ԍ�)��$�ش3d�W���Fc"$u��<�M눸 [,ۥvT���'�FG�� �͊*�9�xO��x7�5�M�\\�XCiX�\��#H�F���M.�$	�w��Z�r�S��'0���t������{���j<Vy�8+|!U�
Mq�ȎD��Wn�|��Q�)Y��ǘ/wr�C[u$�Y�.�-��j�u�I(@�O���3�
4Cc'��yY�;h���)���N�{ӅE�1���?0�γ@Ӯ��B����;6:�_M�pݝĺn���3u�,t�>)vi��t@[�v�&B������(U���е}�~b��3�$-���(M��8:J�
}k0	E�c
��Ȱn��a�.ZPe�7�8�8��w�!L�����%�ZQo>����/7lL�]m�~�Ul�"HP17���+f��l� �������1G���ޛhpnR��P�*�HK�r��f�4g0��I�F���]���F���0%W�N��-#���'T쉡��{�04f��1ρ��$� 0���Y;�+�~��˥]�Rܘl���o�y7q�J��S�}{�Wa���}اXg����|��}Ӵج�?y����B�n_ ��X{��e*^#)=�/x���H8�%�gФ�w5�ܬ��lF�4ܺ޸��Z%�ʶ0u�T��Ɍ���,kU��#�#��,���7�bTe*7�%�.��v̫X���둚��'��V0�-0������E�����X��6/���{���4임>8'k�����	�_ur����]�ꃤ��)��ɢ!�}J�y��ԗ\|8��S�@)I�\#��|w[.D��FZ�i�.�y�Y��w-+���i4{�+SV\ռ$#~~֯���_LM�L��7RL#ɚKK�LY�I�Y��h}���SKsnz�d>�Z\5��? v@���\�����o�;3�����V�wײ%��u���Q;���Y`�:��c8�IO���&E�c�پ�3,d�X�2ЧKY����H�fN��g,��aƞ��ErU�p�гK�&W�_?d=�y��\1�jG'�D�X%��F#�q�#��
��#N%2��C�
�3�pj��T|^����
%Z�y�)����+*d֣@�>0-I;$��@`=�@�=�vJo&�"�x�!(5Iަ͸Hh[l��)KX\���/���X�������<h���@b3�g<#�<�	Ǟ����t&F�0�5�L�v�%����x����β&�(R��f������
��<�q��R������k��e�m�K��QDW��.���#��V߹ŅH9�<(�����D�H�O����PL�d.�|�J%���<��"0�5��V���ο�ۉ,�j�V�6ڣ�(k2)lqWr�<��PJ3 ��X��b����Iٺ�ʓ�8�eS����It]� xQ�9+;+"�o?�h�wS�b���3	�ǙǪO�P�炨"Ռ:i��^�q�
%�E��:d�����>�PC��r-x�eb�r�bQ��IdSS@(kQ���̽��8�#q��aH_�=8n�����3����1�w��,��.�� <���a3K5�9���0{�ˣ��](���N�O.;W_�K�1�M1Z�u9��w�o��������R�=��z�X�Ԅ���2��.z�*Ec~@�n~ݪ9��|	8��NʩF�Q�j}���z�]p�Is�)2��L��;ڻ[o�9f.l"���SQ#`��QqKì*
�<X~#��K8��0�w��JB�dՓşN;21��hmN���{);���.��P�O�8��Y���M.F��G.��� .���ٵ.��
DV#�d9�T��ba���ԗ�ز��\�D�aX�N�Ӊ�w�ö�����NaH��DZ�u�/�!�MȐId��,�+;�0p	TrZ�e眊�\t<�B�����T��NCq�����i��s.A�S�ʐ�
,�r6�����������`���n��Ohz���R�(9�F�P�9B ������u�wp�M7�ο>I6#_3�.��p�a�����c��S�x�ʁbۭ��U!\F@�j"F�r�V�a�-�ŗ���NM=n��N`l?b̘3�v�m?w�Q5;_0��Y���N��}vE�n�Ta�$��ڙUͺ�Tl� �kC �`7wA��-+�~]m�z�xf����U�����R����͔��7)��ב|��S�Ak��պP+�� 1�u���E=ɍ�,Q�=�"Y�����a-��IdC)�6US���<�~�� ��7�~�\�~4F�;\��O����[#p�ab`��T�K�<Z�.�p�X�8#�:���o�l�24	���r���-���2�ԯ�y_-ǹg\�%+�(X�8�?t$.8���f��W�'�4��G�;�b��kr�*yg�>=�Hn��#W���w�(�'e�t�Ol-��p:���/�r<dlU�`x.��膬c��Re�-��F�J�o6ad�"z�J8�����p<Ok\A̄Ϲ�EH<M�"�MA�/K(�E�3� �!k�0�>�8p;�ퟯ"(���X�'i����ڴ�J��tJqW������/yp����H���$3�1i���<C��\6�Rɏ��� ��ϸ�R�6�<��Q^�K�R܏�s��'�~���a�y�7Y���T�ٗ<������2-��b�^sgvD�"�&%�ކ�_����JJ)�>����w2V	ϓ��W(��t�<|.�;��X��sMY�mKް�� �wa��H"���ě���[㲋�F��[n���^��tW�"�0��%�;n<�;NBھ�C@��1�,�|������v��睁����E��
�!m��(tj��8���*�g���KQN��|��q�:����+/9���4����B:+:�uS�i)�_�jn	Z0�y߽{vG�.��˕^0�ҎpQ*M@2�p�v�P��B��=Ḽ͂ݴn���>=����.\ԖQu��spEҀKq�� 6 $�^*��"��L���	���G���b��z��i>���Z4�&�L�C��9?*M7{���#��>;U(�0@/U�?�a����I�������5�/�sU%��%��J�p��D��-���T�rǁ4�X��RMx����@*��f���/�<��m�nR.yΩ��	�$$�v�0�LE���r���HMe,��K�������:(<a�n^(�䳥S����.��X<~Q12�+&��E����p2����a�{���_p��|�a�s�$EE��v�}��=���w�Ľwߋ��JANq5Gu a9��RU�a:��i��w^}�c���Ju����]�`�B2d	KH�^��"����U�0�CA�iN�w>�4Fl�-��\z�Y��7��
�T�资���0���$F�������:h��F�����4� �޿� ,�ry��S6Ḕ('�௖d�=��жZզ�����왅4�CeRme�a��<v���9�h��qC[.���7}����xu���Q���d�Hi`��s�a���g�䤺�,pp�s�~Z����
���(�@Ij =8�0E�&K�(�]�n� ��i�'���c��u�N�\9Ɠ��M�v��E�Y��j���2k ��{A<_�a]��`�0�7&��GYy��>4�n7�z"핲Ǐ�ײ�ː#k��s��J4����"�c��hK&�B�����!�e6V���XSY�t�T�s��T"=��H�����Y�R�n7�nU�ISA]7v"����&$���LA�ί��#��|~n��(��vN��L�.wݎ7��w+�Zg2N������?� ^x!~�?��p���ԚbF�91�KS��}���s�mw��ό# :�B*�!lb��h�N>�c�͔8�2?]��st�Z�*�c��� ���:���y_B�!��R�g�a�.����xg>jM�� 7��U{n?u�X�k�+F��V���W#��*.)�R�|�g�C�ˮ���ѷ�g��.\��]	;n= �g|��yO۔VSA��Jr\6�;�l\}����w�������9 +��	0�u��=��r%�y��|�U��Ӥ���=�=q�Y��[#�s#+p���>���5����T���BH���<�@�����a�e��c_�4�g�>���o���c�L�kf�$���N�0�NP���vq��$-U�������4n^���?�UX.F���b��<@A��!�%[��,^�e_�j�>�%##�8}�A�yG���̙�,���^��rt%U�5�3�7o>�ʯ\��5��H"�DEz&;�[�yt̞�ᒴ���%]!�
U,�יĽ(�@K)>�]����x���0�����c悥��*���]�xV �t�Di$�
�J �V�}��r7�ybES����l��F��/��tL|1�9�ǰCiy��uE�N���	�Q�2E�h�T'7�����i��+��sv���3ov(���Z8��hs�d�il�fOC
��j@ots�����vJ,�Ƣ�s��>��{�BLP��	�T�i�.rW\@��~�u�뒃[\��`=�HI�8l0�5y&�LZ�!ć)y>*9.Sn>�s�o��:����g��gK9I���E!u���$0x���!C�����$7��t��wނö����Z��/$�����_��^�K��Mp��v������}Q�[�j�����8쎛pŏ~�1߃�곕�06Q��l�*
b�e�I���JaO���Z=#�%�e).Kh����U��d�PҦ |���}���*'�;.q�S�.�'�HM�D�T�On���7O�j/2�RF�<)�4$�ԗ���Z�GEz�G=�9�̒\���ф'!ӈ���&��EJ8����I@�4@� f]�?�'lW�MH"�o6��!N��P0{^���y�$�s�}cpǵ?�.;?��υ�����}�Q���@Pa����½fF�ι��vǔ�&���r�b��oY�C�P�O��a�6��������1v��H(Ůǜٳ�3���*Q��~�@�K���}}���f�~(��C�tR����y�Ey�+y�*��9��h�RYƶ<�rB����3Z6�4��aW��3Hm���X�W�ƚ]��F.�{�u >zo�X+�� m�пg7d�6�W)�+7�|W�|ù���f�鳱����s�x��7�T����E�цN�떘;{�N{�n\F į~v�"ʙ���f<��8,h(���l}�Ͱ�;���}�dG�K�`���co��Q����#O<��+h�a�A���Ug�B֏�&IdC�`ųtU�,\*��-�>��,fǬY�K�r�
���%ѝ�G���N�'0�M����J�Յ��"�6�=�J�IK�DId�K�s\�$�����-����B��/�tJ�|d���x�I�WD��\����2w�M��	��ȑa�;�JKM�҆�6�]�cA�Cې�m[��f��`��.N�~%�w�֬q�x�M,_� �6!��h&J��U�����3����!*��ͮ!-/+(`���е�r�Q������xn�Ј�I�y5�2�e�o1�w�;�?����}��_��{�I�h�[c�)��!�2�%�gL��dj(���޼��4��Q"��Eh�L-�9X>^xu�  :�;��q���у�Y	�/����#0hs`���`��X���w��>i����g?�-4z�3u����c�M��/M�AV�G����'�N�R�]q)��0y�!�6�t�� s�,��/N��5���7)���5�HE.1����h�����%W*�BߕPЊ�"'�����p��[�⺾t�ax�q���7>�M+8�H"�$�>��Yu24EYrT���q��c�oG��|�fAr�}~x"�X��9���}�U(��4�}��H:���ۆT�so���y #�p�<�lL��J�V(��̔CZ�3�&E^~=�1�YȚ�-��Q������!�$qG�O���#�O[�P��E+1�7s�r5C�TR��wޚ��w�O��Pm�#^�(�U�����#�fE�/k1���h9V��h%m�	��.V��Y�8E�YHh |	��p�d��c��#0�6�(��il֣7��R��I�˴#�#WU��N�_
��!Ͽ4�]p��s7���yy!wu���Cv�k���W�2�I���Ï��>�w�}�u4]$o4�<vc�+݋��0����`��SO��QH����%��*�ƽ]�4@J.�1l^�ME�*�H�k�,��!V2i��p�c����\�q�ܲҐ��}���3>H�M,ڪB��n�T

6Ir@I�5��/�tҔ��Յ�`���Yg��[#��L�ih���tAZ�5G�T[q�{D�-I�b ;i�8}�8�t���SB\�2hη,�=*u2�l�29���՛����9��ӏ!N�_�/0�����0I/��g֜%�յ?z�"pW	f��c��N����	b��4;Q�y�}�^~�9�|F�q�T���͘�~��V�
f�;D�*�k.C�%�6�N�s]�T��V�H���%yJq���ϓJfe�?h�P���3)��{��Yw,nl��/�b�"����|�rh^N���ϙ�Mo�q������'S�H>��8E��a�/�o���l?�a�%<b���1�ྴ|C�3�^*��bn1��\l9��tKx��W�Z�.�+�	��j\u}|��/kc��TE�����ǈ~6���r3�&h=�Dc.���A��nZ�b�>��)9^;���2I��Wͯ�8g�=�Uk/�SY#q'!�nݺ�����mz��J����OgK��CO�>����a�M����(�h|8{:*B�EtÇo����zͫ��}n��y��(�8��lB6Kd�EBGO��[�|�s�q��Ǘc����FߏW��M�0*z�f�a����Ek.�C�|�B	nSIjh�ep�fP$<p��O��k/�i'������U�|�1D���	�pL�h�8����3N����IJ��o��,*�7����5έe��B�'�����vht��y�H�ĵ8]�p������	���טDU�$TK%�2 �}�z�еG�W)Nu�X�RX�`��	<��[��֨��
]3zY��[*���X��C��2�]¹�+��*+����FD����Y��Q�X��W,�0p�%w�y7���r��xb�h���i��H7�1O�@�{F�!'����$ ���ϙ}	>�� �CE!c6���0��|� ^,h�񂦔��k%]N6&�e�8�;�O�����I��[n�&����I���=%���:�"[y�X�T��d��H��o�uuu�g{T5ϊ�T���cT�JJ�'� ޲�I琎��y�s����!�U.�;�D9���CSvb��Aa3�] ��Z����)�ˊ����e�P0sd9p#���l�"���R��=��x ��g���k��.h���ao�.J��'=P\@c�I#�낒��H��[F���'O�[3�0j�2��T���_O���Ƽ+�u�q�0�N+��.��n�o���6�B^'��ǐ�`�{3p�N[HtN���Z4�#��õ��
�v��ͷ�#��8��½έ5gϜ��y�b�z����I���,> }E#oŷ��s'��V��'�E_, �sb/��1�fêURa_����D�[`�I����D[�z��� ʊ1�"ʏO%���7$x����71��ö{�u�iEJ�.8tԡ4Ax��G�:9`F �z5��>�fT��w��k��D���e�i�o�d�Q`O���7M��*��N'vӳZ,b��0bH_8ܕ���D�J���F�P�j���{}kl�� �����DܣO�A���yԙ��>�����D�|VD��a!���rޖmG�U�G������a�ǝ���J�i1͎o���)?|=$�h*F�
X���NT~�#��&%Fl���� ��*�կ��_F?�SO<��m���� ��yM�8�<���0����]U��|`Ë�����dxEX�;���^.�X�����z�Aa
�i�Ʀ�gsWፉ�p�w`��UX��L~'t6i[�M����cH�J��suY֝%2`=�8�1�� �m5�n�z��EK�a��9�SdS꺰�I	��A��oO�K 4+�b+�kA�����ps�Yȓz�M�$���xK m��Q��^<��D�j꜂�L`�f6C�C�ja/�b�7�D���X�L�b��m�I礧'����;�=�O|��wš�ǻo��/�,�s�E����\�j1=�-l�� ��l&]\?��I�2%�L~t���Y��������1R\��Z��I���$��R�2��E��7��I�$&w�	��΍�ߠ]�#��
9�k�g���[�Ɂ˔X��a������nF�J;�HoD�3�'��|t�+e�!i����(�����.���H�%զ��Z�r*��:�S�����.6��u�X��dF�d��9�#R�@�٭�0�!u���*����ّ�&+j�rw"Ms���0S�9o1~s�m���o ���^uHg�r�4��i��C���G�8�H��Y�����-���S��>G"K�,	��1��<�<�4n���7t=��^�Y��髀�����u�B�!�ϴY��m��`{E�Ÿ���	#�F�S����(�A���H�Q�s0�g��f"��3r��,{?�SdD�MIA��,}�l���&������f����/k{D��P��Ey�ܺ3La�����-�,Uu�����د���^U��]t>�B�Ԋ&f?/a�%K�G׌t�L^Nҥ�ܹh3���(���E����&A�Z�&	�?��dK@�����7^�!���3������b.D���j����;�v�~}c&��A:�} U�` zX����v��F�p������c!��QCM2R1����M+����⁃tႩxٛo[G���x|DF�[����!��B����s +� l�;..����biQIU��g��|m��k���h#����\�ۡ�#��U�PiQ>�$%� Q$D��:��i�e�@�?��Ctձr+�,�1�>Ԧ��8}H(W_Os��|윬j��9Q-C��l7�c�w��`F�T�&+T�P����D6zQz�TT$�`��
GI����Pb�vV0'[�'!���b���l7� T|�6P9��n"�\��,)V�K�wp�h�Cz���,��yLMm8�fФ��K8g^Er�8�^ڈ'^���ҕ�N�Шk��Z�xw�K�F��h
G��Y�r��nxz�;����kF]+E?*j��H 4{�n]�ӏ"�9��Dx���9�@�ۀ4�@���e,<��c8�ȓ!�O�H��Lގ��VD��X^x�	�u!��5�I�;�Э�b�����B �JL��zc�G�� ~�Ax��8����	�¸WP⶞�}�Z����㲣w��'��g&M����B1tQr���}�`�f��iy�_/㻇nK��p�}�<���(c��n\1G_�@�o��V '���V�}���5�5��4B�\P�f���9 d_�ۆ"e���+�v�[-�B�~{N�Eq���;���jیtە���t��j��������>#8�U��i��������$��JT=߼�$J����F��Ƴkh(U=�,�RTC��漈Y�5&UD�JbX�=s��W-��I�߆�t������㨃vC�1b5h�4�
�z���e�`s�����Me>�s[Z����ۈ�u0G�,_8�q��f|:[��
\cŹ�&D�q����۞��g�-��T]Xե���a�~+W-ƻS'�{V��	��I��Pߛ�����N�-IM$f���My���,�1jK�s�I�k�fx�W0{��]�s8�;H�?e����r�Mw\w�5���?�g_���h" ݭw��6������m����'��_Ż���F���o���ށG����6�o�����>��v�|�C�Vǋ��%l' �E��ȑ�*�@6U��N��ǵ�k��ZՆ�Y6��uh�;�qu�!2ns鲗C+�J(9ߤ\�#Dz$�mۡ'T+��6��0��y<ìx$��\��lĔϻ���Kb�Q�3�]���sh���0[��$���"z|�p��F��ܥ>zfvھ?v>9χ%���>���q�B���E�Z���~�UE2��,7� O׿Dj���e�:i|:w!�CQ��hl��5v0��,�=�6�{�%F�����VHE��~	�V▛���=9`�'�p���&d1k�
R��@ښL�a�2��e܋/��Q�SN��.�k�_A#]����2�d��]�s/��|�8`����?ĕ��d�T��yr��+x/��<�?�z�7b .��R|��bT�NNΊC%��-�Q)�Q�A�T^kR���0sDD��BmP�b-;��XY�1O�V������L���u"�EKֽl�Ƹ�-m{E+� �765�ր���1K�qU�oMlCuxaoLU��ކ���y�v�
�Sj���'�H"�h�U�2��c&K`4��wfᣙ_b�m�Ė[�E��zUxV҉�7�S2x�������,�z�{�=�=*U�NE�?��<�r�U
��
|:�I���������e��������?�Qh N<�̨'s�:�������i������+�v�X�0q�gXQJG.Ta3ʥj+�MyB#%/]BL��:^{����X�8�C�M&p��c�F����|
����?����uvۮW��jY#0������c0c�\��s	M�^t�o��3���^R-���.�0��x��G1}��ٸ��`p.M�cK�f��T�bH)��� >Q_�77x�����,S�I�w�̠��X 6�\j��9�����io��P���PT@�)�6�z�(��� b�>��Uݻ��	T8��+�|�r8��j����ۏ{'9Ǖ?�-�G�M��c�
.�*�1�p�rXn��]�`A�{\�LGC�|�ԩ�!���Թ0�o�a�B��Z��Hg��
N$�D����U��?���.]ӱ�������)��0�â�^|c�llֽ]2zt͡.�A��ϒ+�hi�%Bo���s��t#���`���Du�F->y
Q�x�����ԡ4�-	�^��K;���Ǹ�_�{���|󾨫��$�s��Oh��IY�X���� }s��	yA 0CV�Z8q�j��'����M�{ɥB��K�'[/��R�$4T�/5C`��B<;~"��*R4a�7�'8�$c+�FNBf��)k��xn���ҋB\-R�	!K$���M��:�CL"_���#L��cA�I	�%W2tT$��c���gp�%~7�M�A��JYQž�*�З��-�t�"�2RJ9BNй��X-�{�����Hʋ���a�2B辺�n��sP	��t�ƿ8�L��F�JTȴ�ڶDc��J[˅��]��*j�16>��IKb j�i̵J\��/��H+�����l��#�	���y�����������1��`�H�0�N�wG�[Oڿ�A�v$�Ȧ+ma�����t��c�U�S�l\�"���E���&*�'4���SU����DQv$����C��#�TT��Y���J�+G�'U�r��/��>N>f��e�7O&^���c�HՑ�.��W��&xR`��-�lI"Nf��`e� \ܔ��IS��h
�i�Xc�Cw��b�m�\\�"�Mt|:�@y�,ۀ(E�jB�6\�-��O���Z38Hn��s�����H���&��ժ�?�&�)�r���d���x��#fC���/B$�)�Z#NK�̹��G ",?w�mF��ח���#(�
8s)�K��ڿ7|9��e�4�JRzʍ4�'�o*Z"�m�W����V���P�Q�5S���6Kr@���MRi��'� ��!�=�f!MB��G�1�B���J�w�C�:sP����ЊW���w*D��B�0T�It������l�2�T���tE��Id#Ë9��E��Q������uZ���ʑ8_� �DS̈��_��Q���,;l�Rd�Z<�@T盙-|Vq?V��/Rx���8��ЯGWR�MK�H!ʌA��%\\��W��p[�|��p, e�ׂY���M����E,x#�<���(٤z=�m�ұIeU$�8]�pR����rȗ��j�p`fL4JB�cp�M0�\#W���Α�o"�ϓF*�S��'.�0*]QYČqKv@"�{	�5�}|��L!�g�Ht�W�|Xue@S�c�G����ƽ�>��I/cKJ�Ȑrrhh,�^�����Ay�j�oB�E9Z4�{�������uU�wT��(�
ҥD�H#�(F��1c��U	j�a�$��iO�hEzB3���G�Р�ML��bh��h����b*�(.���LJX���J@7���T�F�Ca�ahpKҒ�8f�O�{х���4+�k��bPgR�`^H$�D�'i�ø2��֌yIRӹ�R�u�T�����[�xJX��ԅM�BI��j��$����o�sE)�%4�X�-	-�,���z�����E�pL�^� �&8�-߳�,H�Z>�>�ì��7�m,ͳ+8# M��s:,���=6CW2邏��J:� V�,�En�I�/!P�<����d����	TGh��� Sv�j(��#%>ᰕ�YU�:�|3���2P�X$���	�@jK4��q����Sc'H�cs�z��B��6��0���Z�}h�4C�E[O��^S�i�p�^���d�W�����!}%�"�K�L8+@KqG)#��C�!l������chM(^�PR$��*n���j�g��lB+T�a���E��N�V���FG$��w{U]�,�o&������@�Y�Z�s���H"5e�hF[�6�V�\;R0������#N����*F���������8�҅��-��p7��f�8�s��">��f�|��S��c�f=1"C���&К�'\}��gCm�DJtE�œc�ƈ!�c���#G���"%�)�h(���}��´���eȒOC���I�E�(4����>koHm�К��l��5��JdWeskD�;DԾ1����99W��7�P4>Z)���2[�����6p����
U�+jN�ᛗ�	���uO\�J߿�Ǳ��e�5�}_���w.f�OId���U@�x�e̳����Ŗ�n�Q�VfUGI�5�l�5�	V�-r��3�1��F��r
�l���}{��"'�6�/�B��b����=g!>����C1��mX��Α���/̃����(g/�JΎ��'z��h��Z��m���ڀ�6甐{󡔁���fd����p���Q������ A�p"�$�Nii��1�fh�Z��=�C�_��<�೒��Y/b!YKі#UH�trhr=��7�i�2|��\d� ݻ�%tmr���fccM�(q�++K�i�K��$��/���7����+�Hn]z<O9�(պ1�5_��7�����ܶ�[\�ω�"L�s���k�9�\*у@�%ab�%�H"�l ��$��2,�*��"F@�-C��U�WQl*G�	תvt:�'��,�W�(x*��^����$߸"�� RNvҒ��B'�����<Ռ�2è�'�D֙0턯3���^}y���Ζ�>ݭ���6�v<���W�����l�����h8�ٍ��G�H"����\޸�60}ʋտ��R+�ƀ�y@N��j���dq�X@4.O�
����<i�P��5*T(A��MݗY
t����D6m�dj+�U*��c��Ӷ.��n����R6����L�uP��è�/�W��Iޛ�*$l�$�q�.V�(���Q���y�����;m�tyC'Q��.�1�� �?R���1�+��"�f��"�=/"�j�Y)�D�\��������M[B�%̱�I����:�u�onp��S��L�����=�)2����D�N�� ��}����M%�H"�(��7�/�t�ʸ_}.1j|��1��I���h�)�d�xe��Jm&��j #\nQ�3�~��6��a|b���5"���T�(��ә̭��$�h�y�xLg�|i�U��zC�m�D��~�=/��J;KT舘tJ�e�����&���p�q�w"�$�1;O9뼲~�9�͙V��tB��v:a�9�ͨ�X�8vR(lC�H� ����՝�8�� 1������%���Fj��c�l;A�*��� :i�3;�&�aJ��o8N�kd~�I�v3ҷ(��~AD�$d�W�i�GɄ�)ʝy�5�s��Xt�1�����Z���Uxm�mqo�tjnP�}Up6+�b<��6�DiI"�)���Q��֢���n'5���j������s� �r�f�Rm�n�Dg)�;a3` �-�:�����Ī{T' u�����z�}��EHlcȭS0��k����J�k���\��G0կe�+�����<�߼�-��oK�J�*��G�HČ(�I$��K�"f�t���c���;)ū�j��*}�J�!-\'�Hg�M)��*V�w�W^����M������J%��1Lr�=_yC��lHR�	]]�괓DI$��A�{ �H"_�(Oh�]wK�
U;ɖ�n�
L�Vm� �=o/YW
]hi;��0Kl��%a�M$�D�'I�h"�@�4�a	���ϱU����8P3csÄ�-'�h����{��wݏT*%a�����	�0P��9Q�� �Q~oK8���--�A���,�JU`O�nH�#�K�|���E���RaZ��io����Ϝ�����{^�����5��7��5*�DId=��Byz��",�W�.C,y���r��q	���ы�I�/��u8Xm.�" 7`� e�,@cC�"��61�w�.@������U�i�� ���r��lއ�ic���X�x��g�|���g�����,5�������R���p��g�Y9&�hs���S�Xޮ�gq<R�s�Z&6��DId���&�HL���>)&w��'Q�rÖ���*�[t���썡[�T]x�R-Դ���[�n�������9&����1��c����^�%��r�<���������>}��׿�5{챪ߵw����6.��2��.�����V�³�>����w,w�i'\r�%�m�����eʔ)�馛��{��r�6�^z)��o��2���{ｸ����7Ջ�+5c;��ď�٥�����j~$�H"�� �����*��qk˶P�_C�ɯ�"V��b'��m8R)�DH�7����"�R@�hAZ�5�_n{I�è���^Z���x�d[����u-/�7ߜ�?�����gkvkGm���_��~��cڴ�xc�d�P}��5j���s�:�r$�'2.?�����j�y�����/���`�ԩhllĠA�pn���>�߿?F�-@p�����㏱b�
��~8��q�m���OƼy�d[���?,�s�+�e���I'���/�X (�W>�L*-�=Cxc�yC�Y�H/*nb(�H�`I$��[l3r|������F�u� "�״.�^�F5YvնZQr�M�F�'��3a'�5�	 MD�% �G���5mh�n^mъV �}��e!�K�ߴN�ʧ�.,ޟ� `e��|.(r2R����ڂ�j���M��Z`�:�������g�������*��26�6i��p5�z��~���	{�g�����C������N;a�}�ŤI�ʡn-�dpx�1��駟�G!�i$�3�;�Cp�W����r�ﾪ��W�K�.���%K�����O0gΜ2��_	,���� �N8A )/��G���o�������<��8���q�w�P�à���q���&N�DId=�j�hh�&�~\b�j0��1�hUf5�I����Vm�O��v�H$����Z�VH���6��¨'7j�#��o3���tS?P�`�21񕗰l�2*F����=��c!��+�U�S�� %/ �᷎5b@S���ĵ��km�Pu�������\���q~��/���w�C��o�!�2�cp�!�=z�ꫯ�o����:J���Xt���?��|f��ඹ��8W��a�P��q���^��g ��V[Uyf��rڀ��1e`�� C���?nW�|"�$��� k�#��j�O�_��x8}u��IEO@�]&�D�&����́r7�v�hL3�`�� 8��
�"��9��7����:L_�׻:,���oG"�%Pk9R�͠�:�%l��\K�MB����ep�����E����h���粮���կ$�����h�tHR�b�-�p�B<���>Xt��@J?-��>b�b������={Ju�i�"��{~�@V�	��e�>��C"�$���,kDyB�^��%�(նa�����JW��-+K��P�勇*�Kd�b����G�1a{�,&�'0T��6iĸ8<v��(GZ�2�u�"�`���{B��x[Mn˹��x�oj�Ơ�A�x���u�] 2�g����o�<�Hz衸��[%��y��;���(�v�a�>{T�6/v�u4]�����yl��_�~���ecƌ����`T�������~{Y~֬Y�}�v��&�H"�t��CtQ>h�f��i�P��ıG�d�-T}�RՒ;�h�6,������%��o
�$���T�G�e�J��0 `�/A����0�Qv���0(�E=W��^�M�|6Ьv��&f�.��h����d�� ��%W�O�>]�c��Ю]�������2�Ŏq�jpɠ���,_|�E���\�avB�X��)��H(��Tg̘!��,��S�����?��3�X94�~ٳ*��y�I$��O��#F}ߥ��/�}��=l��L�����t"�5U=��K�צ��¢��<>�~[C Z�y�1�'��Z�=W�y�� ~��*�f+Ţ q�f��m��:v�ā �3'(W��7����� 8������������^^O���g^��c��EH:��\Z����%�z7S(�8�s�ĉRѯC����V��v�m���G~9@�aH2�I$�E֊GTB�Fԡ���"kD	�:����^$���x��;����~q=�r�l' 0@Ͽ��j��t�舁�V�t���#V	�6S@)=�fh�v_+����(�ը�+P�+�Ȫ�l�m: 2Y<�H��]wz��%���e�$�E�\!������Ö$�H�r���F{:1�e�9r�H9�޽{��y睇��>?��0a*�+�2��|�͒�����L�+�ME�<ZN��Hǵ�W-�\���f��ƪ�ۖ@<�)�n�WD���	v�r�E{E��G�s����`�:#h�썚������qj��^Y���N;�7��7(�`/�]Eh��>�ߕ'���y?�r�i����W�φm���_���Ϣ�&�pK��u�'S$��^��_����\tĿ1��UW]%�L���Ex�$�]��:{O�.]*�4�fh��c��ً��ʅN����	0��O<Q<��B���U�L���g�i��7+i߹QK�9H�¶O*�y�;G�m�o�IK�t{�;�'mo���c���.���+������!��Q�4���dFS����G���Fxm,	�#"R�$�-Rځ]D^O��!�.Lt��@1����h�
�$$�&����t�&W��D�Sp���"Z�!�%W�~����j5%χ�9^tNL�c�A�v`���]އ��k⅞\��_��]c�[Q�H��f7RxCɯnPOƉe*�P�d/[ '����ɰ�{u-���~�SB�g�P�[@�����nx�0]��Z?�:�����=��
yt?��Op��Kg�믿^m/�ϝ=��1�e�]���瓎�L������0��#��7���xT$������m��k��sM㜥�2���_~�����v�ܹeO-�2�.KL)��K/�mQXզ�⚑�'zc��̢�ʔr� m����v5�Pm|}1�y�1x>7�b�S֤QFX��5���(�[m�i�22g2w3S�qQfsf�Z��O�sG��MȦ�6����/��P���4Gy.��.5B�i�K2o��P~c�D�>C��M�u�A�D����l.E�,Rئ�P����Z�"��4)j
�
fυMOl&e�T�#E���N��JU�]���@�<)�4��M��|��X��7��RiK�}�W�m�X	�����å�1��	��K戀<�C�P;�[��AB�����J�bV����~�5-TY�20%��v�e�]����#_ �h��4�sǢ�{N�$��j�J�E��7�9'/�E}����}�gϞ-�0�'���*G���z�_�w�+���}��۔�����mAy��2�t����k��OJH�c��{�{|�l�'ҍL�>:S=������ۻ2��. ��1[���53R��4��������{���SI��E�Ѻ!ĳ�gؘ>k>�t� �򹶣)N�D�ĲL:�>�}�h�.U���9���m�  �E�̜�3�$�%�H:�#*.�V~W�P%�`qe�i��S�Х��8�;GbȖ�de�t��?�%,\8ݻv����/O(��o|���<KY�5��fP�C��$�',�Fir��ӱs2HK�AS6�ES����t�XN7��`m�ڌ��h9Z6�߲'$C��(���,އ@`~/�,��b1�lX�4]�r��5��*�1X�
�f���IɦI"��i^���W���6��\R�l)c�,x?O����"��Z��M�ƀNw=b�ǀ�;q��W_}U��,·�?zg/�/���v�J��+��w�!]�4Xe0��Cᬳ������JȜ��M]���"��3�w��E��~�;ߑ|Q����j�������g�}d�>�`97����[<���"P���!��[��8�ݒ��}�>�s��i�r��aTH�"�����g��)S�/4�kV����>�q�w�B���ac�
b��\�#A����<��?�T��K
��,��<k��(w�aG@���Ĺ'���n���Vz��?�����=�O�3�dDu��Q��
?ƾ(��U(^UmJsC8�:K&.��*��z�.+Nöڑ^�#_l�m�܈T*C�+�зX5��B)X��� ����Ϲ���,�U0�S'�пo/�ۨ�8鸣ѯ�C�R��X��>�wݍ7�yi#�B��Э��C��6O�8������<��C�e���O�/�*~|��1��p-��w0�1��>�/ɬ�K�Λo�;�E�c+���;�0��L��qIŒ�6���B%a�`��[�Xৌ�~@��1���d���̤g�-�i���Q^I"e��G��ַ�%�����>�˩���q�b���<u�6\rYx�*������>��?��P?�W�C��n��xQ9��I��i�ر�LCC�T���c��}������9�# u�ʕB+�]�x���_��~YO�0}b�nLR�󍢒*�-�C��q�d�"r޴.a4��^Q��9f
�_�y�_C/:��YڀM۱LY+�����2��dÔ���KHYd`s� �����S�i{�`J%�=��b�X�H�FL��Z#�/_g�@����r��66;����.��Q˄U��L}��UW��ﾉ&�e��h��l�xt$�.�Lh�p����?8Ql�Xk{fDE]`�ݷ��5xoڧ8��`���POWn��ϰ��������G�-��d���4Y��LVlϗ���Ҳ^�����#���Ǐ��7߆��{P��E	����Ԍq%����)�x�m�z��d�{�����
��/].�	{7ò1W{|�d]w�(2v�(o4�r���T�W"U�=�\�������wW[N�&j�і��=��ד=�L�^t�E�����裏�v���x��؛�˲���gk<G��f`ʀ�������Ё����q���>]�Ϲ�D��ر�J"��{KX���(`K�c�Ǧ�{n�rX��CЫ4�X�*s��p�)G�J��9��?Hj)j�����5|�G�WEC�vE嫋� ��l��L�^����	D��cp]{u=F熓��u$k�Ⳇu�<x�u��5�h�O~�k�ݡܠ�uZZ�&�}���7�OQOnž�p�s�3�)�y��b����s�� �[c;���{d8)�}���ң�Jz}�+�����������~�����c�~]9�EH�؄?z�],\��y��A̝��T��t��gW�V��f��¯���.Ţ�Ex�,)�Fz(.8�4�e7\~ťh*6�Ϗ=	/t�2L�- ��Kt���.�JE�a�IC�e�\Z���[�00-X9zf��A=[�yB�01Vb©A�(r?y�5DV���@Ms�{�N��d�cs�m;l����f�n���X��>�T�8N�4	��z� d�9�P=S91�\�lYy�:e�	빂�������j�R�e�'	�odR+ȭoZ���A�(ǐJ���LjKL2��L#�%X��� �DɆ�Q΃������tL��ѩ�Q�}\�-�+���K�_W'�1Y+і$���0EM�=�d�	ee�C�a�[Y~���>��SN=�s� �P �l�����<�ˡxD�����<?�%߅g;4d.��(�����Z�鑧�@��iu��=�<_�[�/�N�ؗ^%k3D����I��ly���'q����������ȧ��~��Sӝj̈�'���� �9�YxW˛�񏧟�9�;�}ɱ��+��	�ǻKɊc`����mxR���r�$���}e�FJ��}� �%	$�9�Ǖ�R��.6;�n,t�&6lф�� ��3.q��b��ϖ�o�9;�2��C���v�
���qT%q������<�X�:_�?�?�Ļ,ŏO>i)
�����&�jc[��uM��ۚ+�^�K����r�r]IЊ��R��5��U+q���"�Xq���9b���4=�jI8bY֧^eߑ�.�&��ӥ����GD $���a���J7�-R�&��f'����Z���5�K�V�+�'���I��Q�����B@��"�s�'F��R�o����6�{�-<�����[�3�H��=�)�@�I���b,AO.'w;�5��w��c�Ǎ8���˟oƻh)���JE~(�~z�nn�h���*��ck��Y��r�_�`谡�r�p\y����w& t)H�b"ehY�!Mlz�=xͬ��(�p��	©�9E�7�褰Q���jֶ��u��(Nۤ+ʫv��ɍ��"�>;��>S"2�����6���ѕ��!��ͺ���*��_:��#������ږ܂ J�-�R �����g��Au���nnx�8��G� #�'#�oZ�QS16�h� �=�EK^յ��)��j֒A\�H�"��:����1��7���#MDZF�?����~cV��H�I�@T��WE�i�-�?)B۶з� �`Gd۵^m���4p�\�%�Ud��:�:���	5	�ni��F�ma7�)R���&YO6Q�<ޏ�r|��o�h���	,n��6����q�E��ݟ�6m/��bS١N�V��F(�4�J][(�8�fj+:������6�7xsYO
�`�pkK2H�I�t�`Cē0�޻툾�sKy���jw�����0BT��l-���A���n�) 1sz�Rx�w���m����j / ����ĳa������u���<7\�Ec�̨���F��d��s�zj��_�\:.�SED9��f:�T���;)'%��-�4��Үئu
3�ݟ��'�U ���W�l�P����T�NfIC��oi#*�X���Kǐ�PV�k�8p61cY7�
+��
kO�FsojP)"BP�S���*������5�ʆ�zi{�E���Vw4[ƌR��<\.��!�8*[B�j�S��u]H5��ȴ%l��\���W_�-6%f�����ュ�b��
w��hV΋anO',�#6��/���s���a J !e�i�"�����*r!�eG������&�IS��+}�}=���|:{�b�μ|}*)��Vu��_�K�V���ѵ�Jy��h�b�� �nlP ����C��p����8�x����ؐG{=l��a�ѳ��������0n�;h�5��Q�z�Ŕp՘�l�l�B/����OPܬ��!�kN�1��$�g��1y=��6����aI@�[��NX�窓py����Z3dܿ��`I҈�(j�F�A�,�Q��	ڇA��P("G�������d�Z.�wֳ��Z%���¬L���&:�[7`6���`�ܓD�Y}T�0*�J[R^n���H���"��b�l�s)U-o�fG��mU競��ë�霵aH�u��$"�0�\L@͈BD�^_��$��:?��o��O�Du$G�,F�#z�T/p����^w?�뢪�(r�ޙ��.���ntN��5,����Ù����
�{���~Gס(��4��QW� �*��8���ŭ
7Z�c[�⎱�J�L�C�)���y}L�x���X���h.gP�6�E�,Gº��چ���d�^�&a�a��7�	�O㫾�z��;�nT��c�q�57�1���E��=%�H��&��7����ŝ�܃��oN㔀j�ޜ�6.>�b�X�~���n��4�ٵS������Z�w�d����nׅ^�_]v��tP�1^t�䣇]��1c��Wp�E��tB�H�׿�F�N;r�/)`e� 2�4��$�j�l��yi=�|}�I@4r[G�k΍Z�l)�0;R��.�_Ă�HY���"6�+	 mDk��1z�N�����`�c�R ^Gڿ��b9h�k���F+�W�,�O�pK%L��!&}܈c�=��s+2�G%_�4U����-��90�\e������b@����>��V5��I��Xd�趌�=��I�JM��V��3x�<�t�$�Đ:%�\�a�N�`ٸ%>Q�bȀ�z���:�p,[�%V}d�]��ld���i�������N��Q 34HD�.�����^��Ӄ�kq����~�(V��K�û������kq�i�⾿�E!�p�5�Ŏ#����0_������{�h�u�e(r���A�~��^{�	a���0�[�ҶW�	H/����42����M$�Dِ��@�����f}�	T�f 3�U��K��y��j��� S(p��+D�Z?���MW��ǽ��>�|0{�>����	A8��s`���P<��A���!oeP�֞M���EFn�|��������\�C�{����\�UUx|���GD�o0�-���ʽ�m:������6������u�sh`$9+뭄f���s��F2�����W�Ԯ0jF�"TxX��;������*�iI*�G:T����0�)��v��LhCu-����E��{9B�i���ȋ�R�%�}s+�T7�����#�
�q�!�����ݜ�	��рz�v;��mq��G��{�<��A�����zr4��k7��֗���������]��'_�C�6�~�8��cHg��s�e���xC7)��7�sS�
��I��楳���PlP��\��Eh�eʲ��[SS�2f�#�
��s��)U���N;���C�i��v*��4�d1v�D\r�Hl���u�9��އ�=���h��漱<�D�Q?���HY))fpz���7\����S�`��Y8�S��OK�]i�5�Iz� Me���}�.���LE��p����v���鱯�c��$.�AI�ɩ����&�ym�bܩ��?��Y ����o������]��/����������/zA�r9�b���s��ا$݇�GE� ͥ��c�=��s/K�Y�~�1g�4��#c�+|����hh*��1d� �ޙ�x�'��s�<��������G+E!�1��_$�H"Jt�V��%�����h*�h�/�3.��J��\i#ֶ��q��w!�� �\yW+G�+~�����`r�l�L���8�������/�N{�{��+^�����l��[Æ�����h=�w]�&|�)c��!k�hpKHہ$2�������'�xrt���W��A��� ]���4i5��TD�.�#F��٧};l�W��ۛ����"`�#�6�l��7/��~�sEۈ80=�bP��;hf](��y 7l�����f��eJ-.`<�;Gb����u�z�
��,V��S��VJ�3.�m
R���m���?�~X�������λ��T�;�n�u4��N�����s.����6+�9����%綤ŏ9��C�*�ѿ>�?��?���[X��f���[�Iɳ&`t����{c�qf�D6V���<��K�0�Pd�<5��
ŕx��gq����]��r
��&�G�i�8��l����]S7�yD�����Q�GT&SB�\�z�=�`H�z�v��c�]�7��ֽ�^��P7���Qw5��w��u���me\��K����ӗ��mi�����QHXΐ"%�{���=,GWD%�_):�o����	�i"�}&�Lt^t��L�dD��f�;��*<44W_�<�ʏ.���P[�T"{M#�,�e��*)�b�iܘ�ɣ�p�!��F�S)<ibZ���� ��*���:�-�z'���Ћ�b)*>y�|���g�+�S�������$��PC܄ 	,��I���m��}�{����Ζ����i�ݙ;�޹�����W~�� t����с��
��~��B3�b�I�H�NϿ�,z�_�ï��/�߼���7���l��Ũ;m�;8%���x�a�̙����~��qł���g�s<~���
cф�ɱ@D�m 8J!��Bֶ��z�vq�j��&�j�Mӭ�o�1Y���9�t��Lӳ�߯�EK��_�eyMF:�*�M5����#�c�����H�,m�e�U�MD/�|����ó�.$�G�>�;.�Ԯ�"�Ez.C,�^|�q�FAu6��κ�U����#J�sk�k�}�;?���7	����8�����[gtb��̛� w��,_֌� ���J�G�FkLA@e�H��P����������N:]%K�����A�5y^���~���*A���PJ�����������T�<k�G�7k�qC�\���2`�7�'��de}d��~M
�>K��ԃ���b��6�p��VG����;��߫mv��н�ڛ���-�(כRh�<|A0jx!�J��Ֆ#�c*�7
�΅b9q?��⹧<�%C�^`�BH�TT),IN<���6���p�}w���z���'��l1x�9\u�8��������]�7�x�?�J�	�)nC[G+�}
��3�G�s8S �"y��L�'��%#��s��Ȕc%"u�P6Z`�k�}�Y��OZʹ!��q�aU����ى�S�x�ғ�tz��������l�oS�65�(	{�ʎFF��2%1G�#�$��Xb�;���(�7�ݔ,u=��]�FC�м&�a�Q�_ҡ��CCJ"���i;vo^�� �/���O��m�=���>�/}��v1�J�����S^�ppVk@,����ma��w����9���+�y�x������fK;9u�<����K^s���n
UA
}./&�<�f�z�������A�r؉b�r���yĤ%�6�^�d)�j�{��33���6�XT�]���>�x �G���%�̨�-�T{$�R\l�s�;}��>j��S�5�C����Ң�)V�\�~.�I[<�?����Ϸ�
�.�;�W��&sq�z�pՍc��$�,�Z��m��`�!���P�=|�������G���9_��7q��`�#��+(��?g��ixbt�qAI�,2�VDVk�"�q*����ڑ#Q)ds��&��(�1Q+���n[����V�*�"���Z4�;�Y,_Ǎ;"u����vuE�Z�rD�RLh���S���"RN�-�U���Nc=A'����ŵ��#���u�00�9G4�Ѕ�����p�^�Hg&U�9�U'Vm���'�s�-)���;��K�$mNya<A�s$ߺ���#�@<ĖC�F����R��є�iS'���+6ϷسF"̡>��"�Fk�'�S�s�h�,yN��7��[�I���!+��x�4�X��IF�ILot$�Bz�'���=��������VrrC���Z��b��H��Tw$��	.Ӷ//}����u0�:
\|�YĘ����#�ZX'vE=K�: ���N9� ���K���jW�}���o�����l�/�jήǗ����G'��ȶ��<O���E�9[,��[���+�o���S��7r���_�sy�nP>}��^�.l�8�c`	�I����bU��:�dŢ�ӓV,F��ec����)�YzZ�J"�\dК�:�Չ�Hyaඃ�,R����䑘#i��b>ޠ����<�<;�<_,��G��ck%v�k�b���^���o�%�����4��Ap��`Q��腈vCԪ%���^��x2�M9'���ݬwm�~����I̝�˩ �67J��NSO���y&鵼 ��u+�}�x��b�hRQ���uŃ�)��b_� չu(�Քe$r1�?�4��B�y7�Ӑ�Zȋ��W2�PE$Y��zj���L����
�tp�-��1Ą!�W,"G^vA~
%�ڵL����$F#~{�M0ꚸ�����#K�Gʣ���!T=�U��@. ��"ѧ��9���P�NB����d���&&p����;yaZ"ω�K奇\8D]�(�;��F-��āB}>uGr�(�	ӡ~�䵡<S�5ాq'/�n� �M�_����ƎuFhQB-^_xi1Jm��Q�.ᐵ)]�ۥP�Q�E�` �"�k7t�O/�N�5#���a�'T�� �ͯ����ȓ��v|v�A�QuFb�]�ayr!r�!����'`�9�䉋9<W�7�~0�E��B��D"$)���C�H��:aT)���(rPA3,��"��~ĺ���^�gY#�Lm�	"��4�rt��V{�m�*@�E�#��x"���b�LiYď(�P����G?�z�D߉�xE���5 
MbDv-S^��'uM�nΡ
�BzC-'W�P���ҽ�Z �����7�ơ�$O����.]G���p��z>i�Iƍ�z(��9��yKw��{/Lz���C!tɁ��y`i7EΕ6S�i�^C��Dr�R��Aq�LU���ԖK�ȥlu���I��iB~6��eR0&ɮ|i1I��<��r�raj:6J��$�yE.v2S���K	a��'G��#~�L�x���F&��[�d�qy����y���G������.~���"b�Bȹҋ������qJD4.4��¬z��HJ�)�-q�B?���ً��QR(Jۿ�t9����)���5"��3��"��j����S�OT!�f�C��	*�!�Dbme8<AJE���T��B���I��8(o����^�؜[��Cӱ�_�q;,�FBP�-�_��A=���b|_Iv�R؛E���(��&v�E#�4���m@��KM�{Fp�a�-�}�p�ۈ�%K�)Km�Nm��=Cw��p+^��z�t��`�_/-^r�6�WJ��r��gL=Qr:O����d����r���T�fձ�cG�8&�<7#�f&����-頒N�g烦�'OP.�;?r6����j�P:�I"W����{3Sϙ����8RD]�?�࢏9���R$R���K�j�q� ,���JK�p�R���/2�E6�s$CAf$�(^I��"���Jj@*b�������"��U��ץ���,���[��r[~Ю���ΡL{z(Ll�%&���x�-���"M>�r�N4�T�������"&���6e�6%��\�r�t�s�_�E�9pL٭+4�x��znl�Os*]-��N����Pޙ�8FRMC� �Y(��6�B��>jMP��	u^���q���\�6!I��q�<�V(=;��~��TK�Ir�@���*�=�<CW	=�b��/<~U͒Q�����K��H���;�U��?�l�>�3�(ӞK����ei�]�Q��[�X5��������fl����An�*7J^��2���(9��i�
qJ��dz*('�6� �#0%��8֚~�+�AAO���N���TNP)Z�+ERt*Cz��6���h$i�2B�G��	&`�VS���1��cǍCcC\�֒��(|���:�Z�˗��7W���o�=Z^���}}�R�C\��c!'j�xl[�uOt�<yAGj��JB=�krxaC�ъP"��"��(#���+YӲN�n&�ء����)�?�p@�z:,v���[T�
C��	��adI�T�d�WdtO�x?i��~"y*���|��ͪGO�?�"��?�:�Pӈ���8C��_�y^��&ˉ���]%�$W�i�٣-�iP]'h�U��+$�c������WF��G����o$��N�>������� 1d:W�@�n��I���Ѡ!M�1.=`l3m
�p
�&s�` `)�0h�Q0���Y���SNi¡�m͋���]�>�"���sX��]v�1��X�5ǎ��)�Z��n
t%��GD��o�`ǭ&s�<y�M��9�S�6�����uw��	C|�sk�@�� ����_���~������3�Jq��a��5)���z�S{���se6��Mu^g�~�~��>,#
�,ӡLX1).F�0��CT���(���b=���5L<�z��lQ��o��0y_f2f��Q�˔VN�e�rz��3�BM����5j״��x�۪�1�_|�3:ʉhEB~WT�8�<�0*��3j]��Z5ׇ]�iOH��(/o�	#P,vJ�~���1�����C�y3d�F���$�_#@�Ԓ�Hi�r���Ӹɟ�2���9G>�y=�کbҴe�#�I���o(�iE\JY
�4$��*���F�*���}Q*�)~�JoHr�2�]&+�6T1��jۿ(�'i���}h,�2l4:���&��ˊ���_�:pt���7�_s�&��5¾G����L#��e�q祌�>���n�H��C�c�r�,�&���N�C������'M>��^�a�5n4<X%!�2UȐ�g'��E �A�ɲq��pجx`��x��gX��t]��d�O���:�ժ��i}��,��P3�6�،���ϰ1!G�!	~��[W'B�����>P�T��8�(^�n��Ң:&�2_^m+�%���yȎ�H=+���5�i�^-@�-Q*��
��t�K� ͞��D�D�rI�f��f������7
���b��J*%�(�p��I��~vtt�q�����a
��e�!o�,�i��б�c��vÍ�ށ�V��^w�f	&�����D�:M��"^3�K�&W�'��'�i�n5p$�I�[*Z�����\�T��@��!��.=�S��I�U�&�	j���j~�v�	=��j�|3�p5{D��&l��*â�e�.gc�-F�³>��Mub����z,EDEh���0����-Q'M��]v�	[m��'];C�k����K�`�{�r��эMb>���А#Q�v��.:�c���;���wQ�T��\ա��#�!C����jjR%{(���qJ���!��d��|Yq-�B��{�H�_����Rw&���q6�f��>]sQSP* �_-�IQ��:Y�F1�4R�@���rN�pM7� U4t*�i��3uZ33���@�D��О���o��'�C��"rV��w�9�h��7Y����s���Y�z&o9'�x��D~&�� ����7��6[�?
��%̟�6lX�Q���K�X�G>��N׈ϟw&n��_��ٗ�	2j�nv3dȰ#�ΣZL~�Ll����q��OFI(�I�c�S!�����B{������&N�8�p0��p�iH%
��U%�嗖��-n�f)��Xm�ڄ��A!u1�L��%�99��rO�H�#�	���_z�6/�$YiS"���A&�
P�����[��:�NȪ�
�e��B:Kp]g��)�nS���E�	�z�J��;��y�������?6tt �wY�++ؼX��f�}����Xe?���ݜue�%6)Ғ]}C6B��q�qG�a�X�z��*K�К�i��(��
�w�̽0k��▚�!)�A,bOݐH�;������^��jG�-�;|`>~��J�(�V����U���M���1έ3�����Gz5�qj(>���:'�/a������G�ަf ^��ו��^ph�d8��lë��"�5�ge��BSH��D��Jʚ�,�m�)�]�r����e�~7*�����8Q����F|��є�&(�Q�������Ǝn�K�I(�,�V�,`/�4iPռɭ-�~��twf9���vL?N�`V�+t@�|��'�U�ay�Z���V��uG�y�J}�t�� ������9�
����F�Y(�}��>�W�+��<ʉmwRL��>�}�T�2���s�u��r��Cf7��&iPlGΎ�<��>m����X���f�g�cCm�EU��`��qږ�D��z����2����Г
����q��Z6Df��Iׁ�%�M���_��}�<\چ���v����&Q��\��eE�T2L�M��8�┣Gcޑ���`��(����y�UyDnr��SN:A�N���9",��t�.#���&��]=F:L#ᵷbҨ\��30�bT�$I1���	=�#�|z@eOn�'EHM�{2Da$��D�r-nC�<㓸��[1����͉U��Qb��s�)���?bm['JL�(��Z�E��t��?���) y�#����0��9I�ˌD�ܐ�L�S�5eW%�����/b���iݾ�qh��JVw�C��V^'w"�/ҺuKv�
#��!i��B�D�����ǖ��[�4��&D��fd�<�j	Dǧɖ�7�D՘��؋}Qs���/�7^=�$�F�����v��yu"�G�ָ��\nöb�< �������E�T(H�.��{�׸�0���C]N�K��CS�P�?��ȍ��(R0K���ia �J����IՐX^o���=sd)}����0e�����{=.�W�}�Pu��i'��lI����B-���Xd�(#�|�-#]x�z�e�X1<q�Q�p��o���_����A_�&E1�Obr.��xk<�-��zH��1<���1�Q�����8���ȩ2�`ޅJe=�SOý���ɉ��V�>�����M8�������LV�^~6���E���+8��%�Rj$�Yh�N�X��m@��ss Ӵػ��^Y�R��B�i�a-��~!"2`�6D� ��x����y�|I�I&��vm\��+Mq�v
~ �=�&e	e���t�r4mABq�����$��x^(t�=�g��*����b��e9i�[����闍EB�y7y�c�Z(W9���R� ��Mmw��&�y�BKV�V���.�sR�]�.�|��` y��my��)���!Y���/�~x4��]2l<t��N{$s�BJ��	/s��d�6�}��{)Z��Ø���u���4a��#y���Չϛ3b������t����N�`�m�"oCM����B;N9�A�DK-[Y���������9
��rF�-�d1�
�I^�������}EC���+74��$ǏLa)�p�U���[S�����Α9�~�%�=�s�����+a�ٳ���X9��PϬSC2�p���]\ւ�%tG#W7J|W�=�g�AU���э��Jk��$H)%m�o���kms���:�f�sA�HE�n��c�Qu��u	��a]����n�ͅzbY�|��ʙ�`<4�51u�q���;:����@D�e�ڲ����2���σCצԎi�'r�����M$��'>�F�*7�=zrQ�r߆Rcx����0{�67�QND�Ѣp�%�*ԧ.����0V��l�W`OTV�x�Z�iCL�9��vs\<��E>�#�(w���'Hg�+>���$x�Q���;`�I�P*�>�⭷�ƙg��^g�hi277�c8��\N=�4�|�͘����Q0��َc�:O/~aCReCg�!�ȗ�Om�N�~'{K��M"
�%x�"{��@P�U-q�����o��"3�=+6�Qc�"������q)���l5��9y�碉�0U;D�,]���E�F�~��K5�68y'Į�����z%�{vS7�G��<�,:�B��brG��KZ ���s� �����-KQæ�X��m�yσ��:R�Ɛ�О&e��Z�<��F|�S�F<���}t�W�r."�N��:t�������̰���OLU-��Б�.Q2�^p��3/��g���[��+�8�Ѓ��f������Gl\�,ܔ�l)�\?�4��9+��{�N�#M����5��qđG�F*���icp�H�2ф�Z.�;�8<�`���x1�:&����?�P�U��s1��I!����<�XD�X@�t�=�	�?F�7K���6��Q�pG�$���ZJ*By�m��fɷs܆�e��H(%oFb],��z�W+:�=��"MA��"{>I�p�Z�qR8^,�8��͡(>(�t�ۧ�"{��Pn&�@T��  ;4IDAT����C#Y�[K��.DB�B�v����e�G/(}�$���0�,ܠ��Tb��$�d��8�Y'N#��[��
�c��ǢQ�g�a��L&��=˗S2Zyfl�5@z!�=�Ѹr�����j�u�]:�m3F�x��e�ׄ<��J;���<a1Q~�S8LI�l �G�7~�x��y��s��ڊ�>`<��B�zI�v�pBNv�{��7�Q*O��4
�����)U������q{���Ϥ��Ǟb�D���EJ�<�.�?ñӗ+
d>gy�pW�H���r�����D������r��^Q^hE�~�$p.�/�-m2�7��,M�/�O����io��a�R*m]����-�+�})����=�ՎX�)ÐG:�����e���{�H�n�����Uy?T9a�Dc��g����D,��]v��9D^�:�0DG���O:A|Z�h����T\1g���/�aԨQRA�>qt��=|�%A2\�	,+�7mb�L�W�Sޭ��#Ʈӧ��K\���>+<r�m�,5+7X���;&m	��:�o�������SV�c��ӕ��"4?��:3��M���0�y��
��Io`�'�ӂ%�оJ�	��o2��}��
���=�?��#�)'���:"�_*�)^0sz�J1�]4�(;_}}���j�Vv3��ɐ!C��]f���wi�O�}A���.Z(3�F��!��FG/�"�a�Č�v�Vq��T�r�{c�&<���̎����m۶m۶vl۶m=c>c����w�����J��:'}���;y��~h-C��p���V�h������p�pҠ�/`�!�G0�rՖ%���(b�8��� Q�4�ͼ��ZV#��W,XM��N�<V�8��Oa0w�d`t�RUSTD"��$�,˲c�lYbH�y*&�%�Gs�<���\�P/7�y5/g=����c�o���~�Ul��zhZ�2�O�Nx���w|�}j�`Q������I2Νvu�Y���2�ud�E3�$9cpǹ;����Z�3��Ӄo
*ݢz>���a��V�@�F��9y}J|B���(���Q���.i���)�ϏE��u�ӎ�����r�a}�!Y�D�h���d��u��I�ݟ�R�h�~V�_8O	�v���:D��?w��Q<��z��\T �2�����b��%�(#Q� +/,�5��OC%�A����YH����x��fM���2��e�����]����)x��R	�;X�)E�!��?��&��s�$w
ST$�	�됑ԥz�S�s�¯�ʟ��	w�v�"/ǒ�`��&��K�B�c�@�f�.w������� ��˳4}(��;�D��\�2�M~&��I�b!�ːp��2�Du�V�S0B��{!������aj�Q���̶>�S'T�\f�J�O�,l�UN;�0,����W�r"�t����@(&=��X�f�~|�1 o����=Q��g�j���$I���qy.ƙ"YDI��8��DZ�Z�km��t=��D�0�jI��:�T��!�q��ĄLn�	o����Luq�]X!�F�-y�^�`V�/��-+�9T���ɰ��0q�+�9(�|.���U{�hE��r.mb�jq���U{QbΧh�Ƙ�ehS�I�VZv�h^��$;6
qn�Ƕ����֊v�9jFFBi��v̸Q��ĆX�GJ��v��T%�r���1�h�i����IEo���L�]�%h�th9�m���?�t� >E��N�g���8��ώ:!����H�=�G�dh��~�����%�Y��`�2>��?���zq���Y�������g22d��d�0�?�T��rX��&�^����u-��s�nHe�3vQc3�B��fc~�����/�{�Z"��S���k�XY�{����Nc7��`����q3K��|YZ��k�A̵����샓be�	'g��;_G���ٮՐ]�+x��1Dm�m��rRa��w? ��2˾6�<�1�-��̸ݖJ�L�噝9�	��]E��Prd5���/��d
�u��m%�&]��k`c]�^�8�m܉4����e[E����G�"i``��c!mOɷd�D��:�'4ѕ����n�v�'n������������碄�H��F��l6�߅�g�he'�8��RM2qK�I����`:�D\��FL��f�5�O��\*o�q��LkB(�;���hT�jT���
=%a���}�fX"#"[y�iz?-�IM����R	t�����Qq0Y��4HC�����P�4k�=�����ᝍ�R7����1����vӰ�K9Q˓V��π�.�]4����������a�@|�6cv�*��g�~<�W�Z����EH/i~�%`��z�B��(@�K����kH�$�(��ߧѣ�B��E�ʐt@⯬�07���n�}�=�?_�#D�e~F�h͙#���� ӒS���+-�/NBv�ދ퐃"2D�x�0�6�I���D#����80Jp�E'�E�ؔ�A�$���Hݿ=14[@x�u�(�u6��͠+�,��?FL@sp��[v̺T:�ni2o�s��q�22N�y�
��M7J"�iE/��ʪ_�_�����C�*wB]Y��N:�U���5�=ӳˇ@�˩]-����ڏn�>b.5b�Tز�/��Y\����C-�J�wXX�ҡJ��`�3���
F�B��lb��>���O���L��Hֺ���FZ	�E'�0<G����Lu-�1�'P�:Q;��vi�䯦jv��G�	f�Ѕ�%p	~%T��Dyت]�-c�5r*�X�bυt.�11��������kDC��E��b�� �l��gF�̀%8q�V�P�cĖ+�4���4�ʷXL=v���O烌B�cR�g��Aj�U�[����z�^�xn��e)bb�ajw�(�(Ml���6�5��W`W�
�� qX���늃i��ɺ�~y�(��5�	�����AX��;Y�V�(C[
�!2J�>����|'�wޕ�"��޺�ޞ�|����5q�i����'�az��4��`�&�~��(Kd�ٜ��ކ6,��Z`?c j뙯^��$Ͱǐ�R�%���P�Y@_B����"�x]�q^s�R��\�ɔ&�?�}�� ������5�ByT���$�����}!J��V�AONQ�Y�К���%)sIFLq��kV<K,�QC\�<��%Р:1&��X㨑]�o3��Ѕ�E�Q� ����-�]2�a]_�I��-ɲ���p��Mk��In�
��������G�n��P�	 �X�ܠ�$m)Q��t
ܣ���xƎ g�����E�d����1L�tF���W�x�q�ۻ	�
͞�ƴ\/V�;I@vk(6: (r0=�jh�o�>"x߽��^�� R*��++�B�
��%������VUh�g-�%��Z�1�SS~=e�ɝ��̦� �5�,�ˮ�#A����&����h�d6B<x����(2��K��E���,t�,�&w���ŵ%��U�魽����-�f!��d܃��&��t����q�����C�[�+I36&M &ߢ��fS��5v|]��]�����߸��0���\Q��m��m�0���ƣ�x�v� � 9�g\5֖4�LYp��I�^���L��Q�T ��k�\J�hH/��_�@��]���{$St�>��fAd)@GѾ&�����/�6}���_2#;��局z87.�LO�=1��=���`�U��x���=P4>�q�4�r/,�8&�D
�G}�����������61�js����RN�CꠙE�������?X��S������VѰ���yv�8Ǡ�+�J����Y�52��O3c$(y3=z���TŮ�)ه� ��PqSw�PyuM����:f�ҕ�[S,���!M�G���Kl7��eѣ�m6%08��� ��y����t%���9� ���~γ�`V��h�����U�A���@�j���r9�0���x��;�[8�w�
�C?Y?_�=�d����ecy�B��h��u"_����z�o	Fj����O���v}�.������
�b?����<���(��������ؙ_{wܙ<F�#�KP͏ɰ_
4j�4���p�1�m�E�ʏ��$�O����1����ʺ�<�g������p�>��^��;+��SM��Ԙ%�PV2���)�u�����!�%�T$���!-���7�Kl�k�R
����@�2>N�"e� a$���7���E���?ɵ��\�{��`��)<[L������~�+A;�u��цW�.��BX�拁<�?v/[��u�`� "݅�l�,����f���礀��D9�t���Zr2��t�G?�IS	���GV� �A��������� ���w�۸|3���U9�rY��վ��|7���`�%��C��߉��5����m��+Ô��VQ�s8@���Q�
��b��--�$9ʆ��㩴=^yQr
AÅ�����ˎ5��H� QAB����U���$���Bӎ�J�֢V��G)X:f���Hj�<y�o�<Ԍg9�Ne��U/��(q4hՀ�4G���ҩ�-�ep�[n�TC�Jʥ����FkȄ��t94�� ���m˃}�|C��1�t"����V	k��+6B��\�$�"F��/g%DE�ts��}ά@��TX��4��<cL���%_|)��D��c�<ٵ����Ԉ���m��Zg.�?�ą��ZB�f�'�GB���eטN�E�!��֨q���=Ш��?�,���拟�Hg��ȷ�|�����Y<��x�N�Ǆ��?�"ai��sq�X��?���RG��	b�5�S�u�u�)����8 �Z	v�.I��qHf�W����a8T�(E�	x���
O�c����uX� �
_TRJ��_F�b$�~�yĶ�	 �
�]Ϲ�<��Q܏�o��ނ�w��t���1Q�����˚|�䠰ٷ�Kj��%�F�]����H�XjK׆��P�Ĵ�r]wx1<mN�iv�e�������evk7j׊�ि�dԿ{;6��,�3�]�\�|s��uT��q<;??�YR����	��{L8\~@�,���J�q�Fd�v�崦��FFD������C�&���&%������Y�$�*�����yGk��5~���H�����Ibhfb�r����K�\=��Tл��e�!4S���[VbTl)7��i�e��Xr�B�8B ��Y"J�-� i<�JaH���'i�������� ���	�kfE<N�M�)YXFyF��N���'�o)<�cN*߻({0������sġU6:n�|7�!B��Ь0B�%ː,�yJkO�LE�!@D�=I��>�E$7����|4l���n|BnQ	��ƶ ���ڱ�����L*P��݆���$�mė�+��,gn��V
�Ő�y,J�iy׏��
���_�X7�~�jn��P���5�<)�g������[L��K0�]vGU4<p¶�#_v��tn)��I)rъ�T�f��+5���pT����w�R*���bO��c��cMF6��zy��wt�\G��lˡ�KP$�Iv�DC�2/�u�p��	����\��1���Z�Z�!8f�4�B!��Ӑ*o�E��X�8N�g���͸�7�>1~���VU���=$�#�����9'��g����f}��m_q~C*�;�3�j�k��OJ�#�0DFlK�5�ٓ�����9�+)�#�'�ˏ�kf��b(��&%cQT�w	�WA\~�Xt݇���32��I ��H���D�oo©���`��+����m��+���LT"�289����KcG��F�/����U[�αm�����p��!�\�@{D5�/s�q#d������ª,*|����W�D�V�m�V�+�����F�8���c*�A�b�&j#-��G�C������>4ti4.z-�_̦OϮYꄴ����o�;�BU�<MD���XN���Ƿ?M�J'T�������؅�����!��	7�ҋ�[?*�T���;l�h�ME-FN�sg1bU[1o �4�#��H�s��͒� ���*��n��R��EӐ��k�����H��L�)��"���������z��}��_B=����V�
&E�k\��QH�^#�G5(��XK$lz�M��D�,z178���熽өNRP�ѐc����9[���[�#�����c8�������|��u��D9��t��3�y���i�9�O.�h���͆�P m9�OS����`������D{��/�ש�T�X�EX�-��~��e
�,�v�Uv��i��?ʈ��mӲ����Q�(��P+� �]�5�k��:���	�:�BL�RLj.�h`�.�_7�B��x{%�~�e���.\��ҖZ�c�h�}1��?I!ڰK%Ń%KϓՈ͘���bјe�ڮi�xug�g��j! ���<��EK���:��ћ*��Y��Y	KȎ�nw�䨾F���kR]�o�	� 2�5��,�����h9�oF�PEn Ę�P�ݬ���ĳ��;#����fd��Vu�$�r�_sv}LP�~��]Ԯ7��twF�Ɂ-_����<�3oK^���r���6��V&h�έ8��Z�!p�=��Yh��q�5��n%;8C�q����;M�ǩ��~��ZDWA��{r��$EH�$NG����Ϥ���a�.Mx�����|����6���\o{}�3"��W:�b̴a���g��������k��݈����sr�`?��{k��A���@�UG��Q�
��V�2;�0��c��c�����	��B��}Uh�n� _B�"�p|�`���v)����]TMN<*�Q_ �jR�����+W���� ~?G�������uĬ�|�lbg��aP�m�Ν,�o=x���z���Pm��7<r��L�ɈA�����~Tq�HAHKX�J�ĺ����_�c�_�*k<���g���͢����!��`����6�(�M
�����_HE��ٿkQlR�/���$��%�NM:��ۼ������l3��A��6?OUb����a|�{�`����'��u�E!����=�K�t��F� ��~Ե�W�`#�hf�CyI�ɓ�h�l�I��B)!p��j�8q���[���R�<1[��tV�,3 ����*�Y	݇��&)�g㠋]�¨�c�� �s\�%9��ol՛k��2Y�©���ƈ�,>��Y���υ��+���>$��5���pH�/�}��V�,QV��^_1�n��f����l���(�{D����,boe&$��ZJ�`���yd܏2�0�q�_�T��_�e��q�A\7��}��~���hU�;y$�r�j?!�hR��nE
���}g~����n{���
r�X�`2T��a
t�xm0#�%�0g�_�U��e�n\��b����|��AbM�1�	�t��\p2�{��iO��������)�Bv2<�f���sCez��CS+Te*>�I����~�Vt�3�m�,�7Ԣӻ� N���2���(*��n���ێEO���o�KD�vjeZ>����2�D�"��� ����s�+����<�~&���g���G]f�RL���
/��;#\�A,��q��K��3���e��[�b�"�y�����W~ꕿP"yc�L�ͳG��=�u�M������H���U��h�#+2z)F�e�j͚b��k+_0�j+����sfF��}�C�9q ��:��+�n nUBl���휔�mﳃ�$��u)�A-��iCB;Ot���F�֖�����a���}�fIadu`�V�b��ܓ�����+�E5]��� sB��N�ȏ��μxJ��⚣�e������R$O�avF�u駍6Z��H����85�줈��@70�UIW�m�����{4�GC�#��boѡW~�]>�Ϋ.��C�!s�T]!����A�\8�Go���������[
O��iDӟ-W�\���&�� [�$V��:ƿؾ�������D\��t��l���QI����hRn��]��|?X�Yd<��<<a��L��!y�h��@�@���^�xf�6�ɜ_�����Ť;��E]����]I8�H�ץ%�S�meC�o���d�!����l�w�-��Z�5����c b/��%�V����^6;�T9���h��1������bx�R�ay� �y<��'8P#^��&;�:taO�a$kE�S���%>�ܮ��;�ݿ�?.�z��*2�,�Ah�����y\�Z� ��=�4��- ʄ�jqe)�& �'�_�=oG-�t_q�p��ku��D�Xa��x,�aho��cv��}�|�J���.�֤���(_T���0L*��,��wJ��k��a�JР�=Ӄ�n;��#�hTXtp����3�Y��}�繹D2q�f3Q�}2�gc5/Qt�%��i�;�=O���+��O׾�4�#9n��;c�T��d��3�R�t�f}n��@�]K)�a_]��b���9`����%6��љA�ȥ6)�[�������W�W񸷵"r�<aFv(�oz���-�Mo}����"����aIc��7�C	�(b���>
�ā�'֨мڙ̂د������R�aof<�T��5����+��w'��xh�ڜZ�c������ț�I�>��I�mwf͕(��Q�_�LI���_�X��(L��nC�FQ
._r~/�-��ԅz�@=D�:4|�Ck3,�Q�v�:Saf��Tz{w(B��JfP���!M��p�|/%�wY�if�:�T�f=����tz��b�xk%�k9�|�[�s�Z�+*�3�L�"��CPIқ����nO�N�Et�����d,�����0��}�V l$/���6��)Uن��o���~���Z�������=\�� \5��6#jB
IG{�f>���C�9oBa�aW�1f�~�꟧3�=�w�k�#�������n_�d?g0�^�9)�[�\��C> ���QR4<������{�k���o��|��r���ߛ�߫�ܟd�}�>#r
S�ׁ�� �k�J��{�~�}��18�Y�]���naۉ��;��5�^2.G5,Mam��u��_�c?V�zo�&K�p��b�E�mWNm�#4���
� D�Ox�4���t�?��O�!� )ߺc�P$G����n��WN���c	5%�!IS���2��f7�(z@0���A���}qk��^����ժA��Q��XO~�5	o��4��󦎺�M�@����T��:�o���A���R��\��<�4�_�M�\�U�'��y{���/������
]r賁Q�F�Q��ε���'��#�&��2��T��z0g��a�%J@�\j�@�n���	�v7�&5�h�6�Y�[GO �Λ���ّ����&r�"�T��V]�J� r;{b̓��
.���'@V�Dh(�D�GQ;k�ׁ��~�x3�M�m�Q����2zX��!.#8�4l�ӶF�{�e����q��h���H���Z�?���XE!����� ��MS���0�m[�e1[�Lo?��Q�<��4��Q/�X�&��Z��2%�Q��T&s}�����L�dg{��"a���8w) ��C�@�;\MϏ��ωR:S�ONM�,�����U'���n�N`��T��f�׊�K�n��,OX��4��O�뀾sr0������c��}��j[��ɹ�3�e��C8�P(,�(E��,�V�����i�T^"D(�V -8��t����Tn~� %=jQ�=�>mF���I:�B�U㒢f�����< ϰ4�`�TvH��M�.�2T�ۑ�=g���mk���p�X.�I&�n�~J6��@,~��j�]/��[kw���GY2Z����_Sk�,����������(|X�W-��~Op��Nz�����C[��0PW� ��;��kV��L�����*��{׌`��?�)q�[���)�f)4/6�O;F�G�mu�!��e�c�����p���G�͝y��	�p�#��**����lIx,w~ڈ��Q �9���k�bx������uòB�����a_���'�Po
�Z����R9Nyb&�ai���hG�+��_�]5;��:[�ni?�2� կ��j�ڮ[�ΣYs��ر����Q)Ҋ7#�1���N��cL�6_������:�����9b������B�A�v�@��͒�֒�P��U���#V�W��ϐ݆�����<S�)�CH����}� D�W��t��k��?j��m)��3A�&B���nh��.dk�������Ymq��A�`&�d@ϝ����η���7"��&ء
����i�r&�P@2L��f��&/�x>��_(���_���G^�>P�De1[�	Y)�������}��s��g���z�K�R�Y6|����.����}��y>@Id{��G\�9��Z!)��^��!����E�6���ЖP���+�E�~�}ww���[6Z�W��@�M�Z�Io���]GL���^��D����g��+�h̜���U�<��=?�3�����#�/g�܈܇�j���#�e2I�-*�v�_�233l��YX�y�N�|ļ�v���4W[!���&��m�yH�oX%��&茍�z��z�4�E�/�S�("cZ5��l|�]rE���K
b}�h��]�^��l��K���<� ��?����<�~����� L���yg��=��k�\rB�'�^Gϴ�\� O���d9˖��Q��2iҀ�Ep�gt֩�~���_�)�n�3Ƒ���L���sZ�G�'���;��{^���B3���8O��N�[=E����3?{e�D6}J�2	�o�����uB����Z3�	�\�⤫!2l�ߧv��vYs����k��h4;�f�}xټ��D�蒵�8*-����Gz�wT�PSb�ml�HD�bI4O%�6Z�U?�J��s�ɕ�[�W��⁍��k2��r|ůթ*!V�=p� �
���mě�̰j��&���+�ỻ���e`�����|�ț�t$��{�}M�	^H�j���V!���X���s������;7Z��'��QE�<����/�&
M�lc�."aq4f��D�mks�n�M���G��Ȥ��m�.�*�ҋ��X��n��Wn�{�ndR���%+h��{N��������AT�n8�ϫ |��1^f�0��/���N��ļ8�ɦ1剱�}P��C5��nuK�=�PA�t���Sp�Ō�.�0�
��ү��٣��u {���l�׭�ޅG��IG��;V�Q�4���Y��t�y�A��/��!�R���3�N�����>�V��H�����y��t�~)���A����� ���C(s�NL�z���^��Pʆ<T��@x��S�l��U$u�'�k�e�����/��ieIV�b�U�bX���v��ڷ��i�9m��s��}=8'����O�|a*N���Q���H��Nn�7c<�(�1�Y����=D�Hɶo|��u���1� ,��~Qe�G���AK���%��v d������.=�&���g"�7/J�ݶ9E�d�ԩ 5���9��|W�H�����ɠz3c���sw�i�Y��]l��u/߄�s�c/����'۶�b���w�}�5�om F��Ֆ�;n���-��%�>�6�<pb���(JV�,4�I�>|^L�7������exA�"�
!D0��U�p$D�	�����l�6�^H�,��[�����^�pMi�`�l�q�׿v�&y�J����G�m���(ji���!���,����ϛ�~��H�Q�L\ډ\jJ�H�b��M8��{L���h-:�3|������dǎ��L���r�9mx�f��g����Ƌ��-ԯ?ђ�w;}�8��t�09} !�@�U��1&�{����͕���=N�8m���"d�hxc�[�#f�����e/b�WL���EQ���(��g�T]���\C���\ �k�İ9H3U��b7d�u$ ��C��4j�m��-V�p�T��\�k�i(	��`��X���_�Sٯ���k�}�c�'���OO�&�5����G��ztb	�z�|	�xb��-�l���������a|���;�.D��&N�&�+`6/'q�Y7�{B�@�U�(��#��r�r��[��s���y�X�i�ἡ�����啧ɦPd���n�apGw��P�E�9���t�k����_%]pL=���P�i�+5���L:Y�A:G��@j���KQ�֙l��j�d�>�ڵ�e�z..��A��v�*�)Imł%�0�?1I�N��u:Bp8~͛��(���ƃ�LF"a�=e�����u�;F4fWm;8���v݆�j�.�cM�&ր�'�1>h��B�o홞��s��6K�Tm�cN1��rk�v�G��.z����/X� .b\pnb=�֤�_��V$c�O�牼� �@�S�Hݦ����~յ�pK��Q)B�4[�Q"q�A�<���*��C����i։���.,"-"��HK%�*�\�eW��ݹg�A{Z~�ʹ�s�f���M��^U��J��H 9�=e=�-��5�� �
���hm��Uw����aT�XM���}���`�B��mT7�D>�M`gP�;��$( s�N�cl��v��/�����tn�q)�����uUQ�ƃ���2�fZ6z�m�z���\�'��kvHNk^lI�h\.x��l)I�W��o�j_`SW�]wH�=;�u�a$����G��`������4)l��f�O�hb�ɷ,��=�<��+��O3|�����Q�œ���RUO����.�HWSVP]z�y�o�_%����<2������3��9+���'��DvP�F妀�[Bdaz�=@A�Y�9^�kױP�L�'�]t�N����4-�*��!����벞���0�/�C��V�_�([�=[>\����~����!jP��ӯ����Ȏ�I�s�Jf��d��ctƓ76�הLH�������r��-N��~�f2m�T�P[Ȳ�����>����Շ�Їd|&J��ɺ�a�P���~#�P>0y�+r�m�O�&�LOH���t�Z�?tFBJz�9��{+��R}["%�%Z�f"�n/v���,;je����:��z��[�'Bd�BFW�!@r�1����ض7�Bt���-�䚷�/��۰�f����4��vߐ���`�z�q�	��7%V��,�o'2��W�����0_�7�i����`I-(��گu�$�j��?�(�rX���a���ro���$��.%�v���ĜN�Nyb�%yd1�Y�U\>+J<Z�'�#n��
%2�Ӏ�pk�ՔӰ�-7k��%Ձ�����H9$�]�+�4��>c��o 	1U�m��u7������Z!h]I �p�-���jYW���b��2侙��O��b�T�ȏ��xe���g�#EB�Z��Ý=���U6k��ښ�.�oWuK1u����P	����`�sR���%�8sR��B�p`����ӭ�q�qӞ��P��R@��}4<h� L7������9��5���oZXx��k�ToƆ^�?��m�ܝq"�VEu&L�eI��!��������'�l]�i����T�O��:YB�	*UHa�F35�i�ZTJ�J!���8O�Q�:���{{��j��l�Z8e�h'��t�5͠<ώ����b��u��[\��������!P"��`�oR� |�l?%�}5�O�oOeh��
'i���W&���TL2�y�o�	�i�f���L�ZP_"�6�,�b2�/>�
���S�p(�~(�o�����Y�@�Ѱ�USM�(���̲�5�
�Z�s0���rv`Ák�T�mWc�ޚ-.4��SIk�CIFu�������\kf_���(�PG5�4k���ڻ�;��E���a�ib��E),I�Lp$+E5Y@���չױ�M�}d���N�x�uX��Jk{��/���5����gi&�ʇ�.��~cyѴ�G��6|���La�i(|`l�����s�K�u�<�[�[2�7]������i���e��7Ko��&E���y&k"y�2̱Nx�µ?.�>G�t�_k�-m�'�~�� �*Ǘ����[���݅YO����Z��}��͌�������z�-�3�i-�U��]`�d�?6�ؘ�u�CV�X��Ԃ:�s��鹎�h�Xkqhk����O�U��$Wm�s��f�o�g�m�u��j�|�~���0��0�YN�?=t�3��o�_�-aWr�֪�vC�>�:@Pq0�}"<#<{��z���������u�\�@7�L{����{ˁ~����>v�I���&}�ݪ�>��J��_�L��[�����ɰ�E�nk�/?�w*�{�E�-�P�J��5X����_6�w\��du�r�U�/쎆\�����.�� ��9�~j<;������?l�� wD^�2�5C�1�2M�>�;N�~�涽D����5�;�cL�m�G��dcQ�`e��� ��t�	�[Z�=�w:�S{&v�|||�y5�Y���9�	��l3#]�˨Ӿ���g�pǾ �Xٗz�GF쿿�=>���.���z5y��?͞2>GnZv�a��-��.�L��!�Am�:1
p�����~��^�[&r)\���X��!/ND2��	�:�_����3��>�m�]�]i�h�O�AX\��{��%���N��n�{U���f��O�+0y�Up?��<I�%G2j
CD��w�������
�l�`W��
�YD/�It}��yg�iqd�����,xw/��Y�
k�'���"���
}�V�� �z���ºc����I��
���PK   �i;Y����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   �i;YF@vw'� � /   images/36b3ed9c-16ef-4839-89fb-9e068aa5b597.png�|�W[M�7V�����w��ݵw�Hqwwww�Cq)��G�}����?ܬu��L��̜��gNB�%����!  ��$Ŕ! �5�G �[OT��[�,!Q>Np�v"f�)e*'A�� b��-oğt&$�����eB��*�F&�����o�U
!!%&��
y�g�m����#��\b�x�.�ۅ���k��U�_�\lu�4��#9*=�i�Ѕ*�l�����!��A}���t�)�~+��c�Pj�p�qY���i��M��̃|��ߞ���K�^���KVq�/�/ ��5�����҄�v?���v6i�jnk�s�y			=��sii����f>3?�jvv6+��ܕ��ҷz,22r�a�elÞF��,&9�b}����dUUQubh�)�����r�~���9�N�=�[�o �Xp�j��Ш�qE�x������e��s%Nwi�Ku���e���0�hSh]��q�pҊ�j G3uu�����g�PK��̯��Owwwu��E��?�R<�3�/>0i�ί�7@(~X�P٘ܮ���r�"�Px�d�CU��9l&m�d���҈�OAb�o� %O�^�FZ�A�ypp@�Q��y�į*gee�������=��G�f�����E�a��;Fl�:�>]���[ĔTW�N�s&E�g��D<����$�J����B�M���/ӛ3
�5f�B��Lz�i��:/Q�c�s�D3��I@iWZt��c�y���L��IQ�#a_�k75$�u�͉� ��_�
X�2��#�}��/6�6���4L���;Ε�ϼ�\!�?��˦��[D��}�����8�6��fv������B7Kå#�v�x��K]	�����+����&O{y)���M4g��&t���zNp��o���Z�GTvE�h���˵| t9�=_��=��}:_���p��R�M�!}��@I lr_����N���7/�W�g�������ҏ��nn�����ז�χFr���������x��C�	��8����\y�ЄYJ���Z��H�="���$p��q00��T KX9'�|������.���,9�[��:�_��O�n�ƶ���f�
Þ��o�_y�o|I�`� �D�2y�z2;{���6�������r��YV���hBA�/O���rΨv����$�����<i���Bu9 9��:]�)]���C�r�r���&�-�ѷa�q�{��h%"GL�I� �0WJV�逴�Rx�w

i\�G	�*7�^�����<��n��*��s�1И���uZO>�
�D���'yz ��j���BL+�[ M�D����_9Q(������^	���W�$oJ��=<�k�6��968=���NЭ_D��^�p�~����+'����#Tj��,h�i�<������zfYh��=_�a�Q�f�=j�JBIvZ�.@G��2���k�|�l]�r����eR1�ŵy�
T����>����E4�_KON������I�3�؋k�A�*���}�"Q-ÙĕZ`+�( cج�՜��~�V�{]T1Q>-�퓎�$��T'Ť`v�)z�G�:�>\����\�I���W�+��f���/�c4:Ι�����MInhRU/���7�G&�k<[�I�����Ig�*+�9������;�p,�?����j���(ǋ����ų��K>?���hg�������C���U�7g������N�?�ǔW��nU^~�6�3ZLgs9Y!l���/v���F���7�t���[ŔϘ��AK1�'+�e�G�>K>vS7Ǽ�#�Î;!pzd�+"�
��И�	��4��㝕�ǘJʚ� $�0	�̂0!݈̃&Z=U1s��=G�h0��Խ�;��'�$*E��r���9��	L"��)�{���?'0_���F��p>�u�ܛ���qs�ѣf����������EH��kt
G���L�<@�xzq��2;���=q)A�A��{dB����Ҙ�bc�J�4�\�3B�v�p��.���w����TA��2|�,�I4��ȟ���J�t+K��9=���]8�0&F��; "$�L�Ԝ&�QV|`�[a�Yb #{;gw�L0���Z��������i��"������;���rȞ���{�Z��|�u��/��Mm
�Z�a��f�&phl��Y�$[��
?�8F<����ez�QD�#Z�*H�G���*2�i�t/�T
c$�J'U.;�_*�7�h K����l�C����ZΪ3M*�a�N�'��=�T-�5D#i|��(�������J�9�2$�h$������G���G�ۻ�/8t�ޓ�]�N�պ[�M����J!��j��q-���ϸĄ����t��&ʽ�5����RÆG&�ʵ��m1ƽ�ff!7�%rn����dgU���uX7����,��� x���x�#��{$s����a$6|�b���U�'�8^'�����x;a;묅��2�u�����+�L�?�$+�4ዣ%�bʕ�J���]�҈Կ�!�XYZr��)��!�͊9�����`�=�E�*%w�x�=
�$�2�Www�/zzZq�����<��l?:G����mϐ�3�C���� ��������|F��x��3��=K*D�nk� ���)=�� ���f�˩�B��;�,��r��B�"��a�ן���t��q��
Ŕ��LM����d`FE��SHi���#[���1��gd���&pC��3���M|,�x��y�������h0i��9����JrL�:�����=���8�*�r�+9���r�8�Q.٩p+��^"H����7�r��iB�x���o�����������G�y��Pi!�1r1������k���_Yv�q� 1��m����l5/����1���,�W�7�I����1.���0tl�*�49,�$sip�w4Je���i0&��Vhoռ������J�S/8{i(���Y�����W�6`��A
�;zd7�0�42�f��F����+�z������������P����Av�"�ԥ���x�o��4ڊY�+-��A������'�Sn�ƭ�plF��q@&ff��DB���S�	�AU�\��v�C.�R����7�Q��в�Q��a��J�.�m~���R`�Y��"��&zl�>:_��E�.4]�bb&�Hr?�3�(0��T��
��`���n����Z����ːcqBx��"�<��^�P��ğ?gT,�|���8�e��J�f�vl���F���˕�k��o�:zz��F/�4b�3�*Nc֞�M��|}���W�"����R��B�X{�W:�0m��;��O& �����Y\�`���1 �ĳ;ΌT�9���T4Xۄ�Om`Q�Lj��Wp����{��_�so�O!bໄxW�"������&��K3B;/�2�"��H9
,&T���vw.��&,��ц�3 �BFGf�-O�g�D�u$��*�<#��EI�^�Y�/�4�߻}��?��ƖXL��+���.��lܚA��p�Y��#��
-�:@��A�
RN3�t��@�����+~�`��������V+l}�Hq	��N��-�5���4WĴ\��	�H�rؤ�Sn�6u@�F�v=��-�e@{Gg������ZhH P7 �v���x��s�����o�qn�Y�0.
QqT����|�חgP�/��Mj����"�[������K�)�q�^J��HM���ckl�g�(���{o"�����[�M�x�b�=��>7�@�]]��S���PW��A��O�N�n�!&]�4�&j0^�0V2H��E�b'��#r w�7�/��M�[��%P�5�����f0�E�+�]9I�l�嫂���Xr	ulLL_㲴���N4:�Շ8�,���A���M����[9���|	��6��z/C(w��[��:���K�Q�Ⱦ0�Ŋt�^�$u������@�8�PW�0d8�jjj������k�v�c��ކ8�� yN'ׇ��"��޿:!w�CkCiM2+w�\rM�����2:�b���E�]T|���Y$A��. +�ɾ	�X:rz7
G�� ����j�j�7��WT�����`N�������F��Lw����j��|��9�:���1�k��P�R��俞����}��p�/��"�� �����=���|�--�� �n*f	���f�e����	]�-Hr����n�3��TM�z#d)[ڞ����i�=ԣE�%�;�Q���t���f����#��a���D�$��N6����2ծ=y��]H���$s���<��8Z]L��E����ʖ�'�~v��Ѧ	4�tBo�`��i�W�mIx��Am5u1�J�@l���`kBjy�P7�������az�����26)R��*�|�ߡ�p����ޔ�����Β����*����|��9�����f�^bb��H���\�ڄ�'G%�Aΰb�^�H��8Ԏ>��o���u�uY\����k��w 2(����L�;oT����p�zY7���,�F9�g箤�$���h�h ���io\���P�,���펷M͙�%@O�R��W1�����y-���ꀾ-�_Co��!ˏK8`Q����m��DFYM�J�_(�O�$m�#�(�H�p@HH�H�i��������τ�C]��˨[�jE�|��.�6�  +�D�w��,��n�N�P�
}�5�c��9������u�o�HF��+�T��rPT��d���FV������gi6Y�H���s��e���O�]o1U�iV:lAg9��o��.$aW�`���D����� թy>Y����^\|N۱�V��o�py@��؛�`|_&����YҴ���2��H<��������)��m�.������`�O�>r^��.�s�7!�Ó� e�,+2V
��8��˅�n]��opH7��u�.%��K^���Ņ�⓻e�*],�A���J'0�H絇q?}�k����t�a�\��H��\��4�3��xM�?;���V�h;���װ�F
�i	�=>���Ç�×�U�uF��U��>�+��Y�Y|r2�@_��\�:��P0صr��7�L��xh�e�Zp��n��P5���趓���z]��y�����%H�c]U���O}$��^�c�|]�Y�<L�f�гޣ�s;R�c�d��S�jh�HYcpct���M�q�(ؿFF;2�����:���:���-e��"�f��
I�M�j.*��!���G-95h#��aʃ�D���!���!�<��7CwB�n��|�����[��|��_�z#,j�c�1�7��S@�E5*=Y�2�an�ی'�����R%�9��?�1��������Vă�d��|?]]>Ëm��?�t�?��rȥr3��SX��npxfG/4�1sy?�Mi���z]�,tԬ]I.~ĩ��{s���RQ��y�stt�`>�p���f&R���h�"y�aF���l���ݎ�6$�6sf3�����K�Dǉ1���9�ς̱�D� ��~����Q��(:�뿎J`�Q������$���p�'�;<<<�A�����op�0^px�/T�%�DA��Wם~2� _IE$���o���qF����d����߉	Om
º���iG�D�
�%��Ĵ�ܿ] ԖϟO}^� X�hǂ�/��6=�Hm���<��Y2�wg-��(���v򴮽��Y�|�o8i|nP��X�;���(+�ۛ����$WѾG4��bȩ��`d��Ȥ�?�%RH��,inS�l����;�c�Kj������X�sU�U�K�$��u����|9�{����TJ�Jo_�����%TI%HX�n���;�.�Gݏ�^�N[�hQD��Vo�h�Snk��ɸ4T�R�l�붓��i��e
�5t��OG��]�Z�0��뤿�E~G�R�>������������Y�����j��S��F���e��r�Mj��m�P�kd ���)�4�fԎ���*�s
�iX�o<y���I#�kSaH��L[���ӵ�0,ȡ�S�A�6^W��JA�\?�Ɉ��fL���U���)�v��O��VS�8n�s"���f���Fx1�����2��r�Z��}�?����
���S�~�d� g
9c�g���4ꮦ/(5�g;V��ZO��m��9����e=C2�ojSP)4A򱌹������e����&U铸�^���.^!S��"���D=�F�{^ǅ��b�:ɠ�2����~ٶO�
-�zD��qٮ�z+�xz>y_*&���fߌ|h��]���_靃��y��]�tu�d��Bu�!��D`�-��?����jpJ3�߹J!ÿz��h�5���0���jW��RBR�
J�������w��yymJ���?1Dc����{��AM����b�����s;���冥!�_���-9`�L4���;�f� ��{���s� 9�Rɀ&c/�aJ�!|lW� p�ſ��m�o|�g�mʷ�_l Tu���6��9涏!%�������!��+Xg�f���yE��4BW�b7����������n�W``b�6��J��"����©��C&�]m{l���!�����T�řf̀�6����2���1,T)���G�㞱b�)�Gˆ'F�S3?�?��^1��+VXr�)���K<�Z<?ޚ1�y����y��{v�z�
y炁da���0�abᅋo���F�D�x�_OOCrm����ˍ�4�F�p�E�f��V�PR���"x�	������5�`�#Y.�y�̨�,������<�`��E/���I������gN�%�~q��C��ϙ����D�Ap" 2�|��A3:����AO�H��D���������bo������r����VBt�\)��aoq���G؛rQ�*��HtǠf�2������{E#���'�����:�����$���d�!+X�ˮ�?�g���WT7���y?Þ���jc��}�w�9]�B��)`�^����0�9�?|mlȞ� �z�c=��9�S��0�~�ƻ�?wF���c�?9*��h�T�s<Ϋ�}�.���@C��ť�B~7�V���� ]ˍ��׵@?&���5q�
�-�^��Hɗb�J��������R�5L��u���M� X��\��α����U(o���7�x��<-�A	����~/c]�F�FJJj�Lr0	)�j��A�*��r��u����P��:bo�O�
#����9˛�c.��P��+�[U��{�������8���P	Y5-����|Xd�Vӫ�l������7���F��E�]Z���y����yFxS�% �p!�܏Z<X)���h�ʮ�_/$^��t���1m:�
�ˀw��J�#
|
���L�P�7{��7���%I�S���9�6�E���8;��ld�+婗�Y�E�*?j�_����ѫ@sJ(�ҞByhR(�p�2�B�z�r�C�f��Ta�����.&�wUhf,>�g-Ğg]�3'O?ڝ����:K�V�����ª��Ʃ�,�A�RYhC�g�i��K�������K����sё5�V���:1଩�8��̋���0�y����=��r2�������n���K�����@��ul�?�����v�&6f�])�ʭǻ 7��}��^R�puL� ���ɏ\�L,[����	����lS���gr싍�p�{�E��%�4�8����Z�wU��Ϫd���o�'9@(^>��^O)xנ�6P�Q*֐%JJ�4�]������q���F�Xb��OMJ:�/3^=)���B��'����n�x]NGT2�H��P�ѕ��Hk+�D4u"& A`X��a��԰/67V���ƹ�bӀ�p$��˹R�/{	�*�mg�u�5������>�K��������wZ¾�rK`M��e��[6���1���ϟ���4W:��\�����Q?��_�8:P�LO^�k]Yh���keQ�u-H���_�O���1�#����r�n�k��Ŗ�M�K"� ���D24�P���~�ZET�(�$U7L���V8=��u�y,����M���W3$����#��/��ϫ:/��}���$z������fl�1�0¨��s}���F̅_�Vh��إ��ӕ��g	�]C�nO~���Y���x5����*�nD���(-k�R��(�Daac�=���<�a�M��8��&: bEv�!���Ύ�ƨ➭{37��bD��XڧFS��(�(/p)ߗ�r��y���E��f�]/Z�e�����A�"��-�f�����'��;�wt@pu����p�`����T�t&`Q@���eZ
�k�� �<�|���(������E�F𱦇a���h����x���N l��pʮqe>�Š{Y�ڎ�D��֝�F�K��o��B���dڌ��ܣ�⇗��9��ob_��~/8.-�������M�j�JLLrF>��0�+����b��� T4�0����Q�1����l���`KpM�(L$�E�l]W�E�^,�\��*T�N�0G|�%�~�1A����^�B������X0i���
FؐX۱���Ȇ�~��"iw�Z{��Lh=��M2��ZeA K��>A��R�б+�VXt��a�!��l����PY�9�A?��{�%-���
��A�4�ܬJ��)sְP,ic9mrO`w"���5��v���d��SҁB����ȅA8�Et��	�0��p�+��{�4�0�#��l���� _��F	"���H��n^5oI45�W�o�C���b�Vi��-ؙ���=f�3L �|��覠���-)^��?����ߴ/�ǋ�UT�	�����uCq�b���C�� o�j�e�c�����ӻig�:4ú��m�mւv�&m�!v�]�����+�E�<t��l(�jH��M����p�Ľ0��W�{$�eD
�8F<�|�w�*��<F��:���}{P��i�/�Ǳ��t�DV����X�=RN�ߣC��3c��E/�&t:'�~��+�@OĎ�������\u� �e�.��.��ӄmjd��x�B=3O����py���-�/>��� ��C@-,d,�p�������9�M}֬c����yEq�2���WIJ_�u�:���
DC%NG�f��0�������j���]���f~d�ɀ4�`خ�7W.~���>�^�,����x�s�s�5����^e@��J>)�&"Jǔ,��v��,E��~�D���<�hpD�m����, �)�����D\eqa$�L`�T*H� ��6�c�կZ �Yͻd<�.M�� �q�)�Kd�>Wॢ���e��\��Y�Qqv��w=\�~�fʅ`���^���KD!o�LĹ#�/��@L��n��5��`�Kg<�舑���"�\Gà�$�\fܘ��Lc9��͕?��l\6LDv���@M�iK��8R��ɷ&&��y�:�������\88�f^Z���_ST�^]��$0���<�7���^�{�6K��1��W�*�v���i l-PK��� ���w�]h��%d�7h�]q�I�l��?#H��Dc�_�+J��4�o�\s���s�kBbFEP闲�~�����\��A�CZ������Q�B��k� ��C?]c;~%���42(��U��g��	��C?��Rh�N ���OI>�IdE�6'$ƤH����{M��4�4��٦�M���Y�b�2c���7��>c�m��L�KX��1�=�s8,Os�N�Ol�s& u~n1�2RJ"!^�̊%��n�<dK�ȫ�+�[!pұe�侩 �w2߼G�QRN�6z?/&�[L��']X�㢖:�����H�ᕔ�D�|��b�A~V�੅�x���v����n����..�c	߾���	������+wif��>u�	u�����jr'$ ��{=�{��Г<K233��y���u<ߜ
�>L�l�f�f)r���h���pPr�qH%i�Q;\u���1��>f��W��og�Vu�jVر���z�v^V/n(fy�w�]��$�I>���>�~f�����+�7m2g�Pi�3T]=f��aEp�����9w�@�����C`O��?�I���WA��? ��@�n�������$��}���6�P`UM*�3t�ݲ\��B<��.���-����̺�O�S��ڇ���c�Z�(���k�£������/=Y�t?�R V�&F<�٧r=cj�z<�Ȫ���l���&��� ��O��J�q��Mzzx���b^
D�;Ào������XMѥۜ�ǐ>G�:��v趹�eh�����,���#>�B˅�N�xX��/�Zc=����{�c�NE~��Z��l������8�t��_�jI�fE4Ŭ��x2]^�@�c�hQԻ�YL C��R�C_x����E�L�Ooz��������皌g��vmu8&�?7�u�hs
�Ԏ�S��c�Ϫ;��#6�L:fA�{��]��Ar���㓜���je�?/ּ�0�hD@����Q�'Lءg|�$GG��D��S]��[�S+���O�dh׸'��de�l]�]�~�ØrT��'s8���%���%�G�{����O��D9����s���I�)2%�>��-�X��lִF�C&7lJ���'𘉠���Ӏ��Î��E�z��r_���@��;�R"��&�l+�*2��!c�:�j��.7����B$��xj�b�I=��z�����n_�� _8�4q7�i��{CE�0�1N���r����U;/u�34��Vљ$���h�^�_�<��z0�rt�����=o@�C!����D��U��*����.2�߂߸��ۧ+�C����A5[vm%5�,��R�m�n�!se���@H���� �U�X^�}�֋az6]����A�L��B=&���i(bCLdeR����t�{s��z��?:\�#���]������D�Fy灥,_{�`K�D
9�M�i�$�d{`�Vo��;%�鵠`�巜4?�=j$V|j+�������/�����e�e\��Mp����+���K���.b���fsۀZHȄ�R���m�3����T��x�+�.?�� ���v4]�7B���
2~�Vs.���gӘrӨ���Y L@�F[����c����>p�Èfe������_��?��Y�V�O�����W�yKK��Y|BY�f�%�p%�=��d�ôþd��+\��Z�	A�u�]u!������u�TS4p�����(���o��z�NؘCV��ӿ�ǝ�oW��upE�IR����5��nEԗhw�H�a��	��O�0t0�1WI67E,7��:�L�l�{�A(u:����c����J��ci�ӡFG�/�@�`���&��	����u#k�E0�r�::6���ֶ--������:.�B��q��Ai�;�,�b�+S�t�x�z�$�W:�����ݾ�u*�����"�
��$�)�N_��$&�Ĩ�`�Ve�P�[��c��	Z񯽈E;������h�m��2$1r��ͧ�(B^2VԢ�=,�~�o�d�E}���X����M�$�a���4��b��mm1�L@*jN�H8O��=�Ͻ*,BQv@-@;�NW(�,�:hei�I�We��to��y��&�$oՐ%���U-qN��f�>�.R-D9TY��Æ�A��n%�E�S�S���hI)G«!{sZ����J�d���'�aA�����b��D<|�����q Mk���&�����H�mRWۅJ�,}e0C]��O�O�V: ��(F�q��1��/W|��l#T
�+L�Έ@q��'	������R�ӵ6��X��	�&��A��Q���u��}u��-K�������ߡ�5�C�_�[ͷ�E�TBv}ý T*1����	Xoc�a�,�8J}�c����l�8����S���ŋg���"�����q����m#֙H�J�F����Өp�!�_�=�,Tt�վ'��!3��E���y�;���I�p,��v��˥�/���<��܏譽n�3�8[XX��b�mIڤ��U��*�	�@q 
�O��dr�2�>�*����戣�����{SM�n���Qpb2B�*��  �y�r�[��!4,2���yv]�W.ko�{����n�<2-B֙���;��J���MI����.�!�4+�}��$&���H �ߓ�j�J�uT
T�����^�B���η&�
�8Z�ۜ���h�e>L��EV�6L�k��Z�M�~��J~�jj�������������uĨ? Wz+�1���.�c\��+����W�4c����v���v���`�jN9o�A��d���T6��α�a��xm����_Ih�G�,^��Bو�9�/�y��f��\��$��eM�7ŀ�+��C��6��Ξ��cWs�j���vO`��y�F��>Kl�E���w#%-N� �]j�O�$I����kL��^��4n���sYW7P��
��Y�GR�p�O`s����Q�ð����8�+��ù%��s%��l(��J>#|���^��l0Z�������`@>;KП��]8+_�n!Ւ��>ة)(ʡ��_q9��k/��6~��1˗��/���拋��G���e��,�ЭU�~< �Lw�g=����#_˹�v�{Kz��̞WU&���H���B���ur"�&�u�*R���ҟ�+ƈ�ߕ��[wQ}y��Ą���}o �m!�����4ܹ.�zDj��
����) N
�w�{1��5w���m\�A8��@�>��@^�1{u*Ѩ���F�K��G�=�ڝ[�;�\�w�Н�	�:X=��m�mK��k�U��|X����(���`�����033jJ7W�L���A�����i�bI:?��)!j�.C�����(֝/��|m����tZ��H�I�H�L��j�?%�l<+I���tU��J�6n���}~N#�u2���"�>X��2@O��?�Є.�1�L�!�e�7�{���.��v����u�t$rC50C)㐨���*�sa����5�]��6AR��'�mvtϗ���m]~dX�)IbҪ���2�	F���G>�8��|�H�x���!&n��Ъ���pd��e0ܰKh���A�*���w��]~�<R�`�i��߲9x�WS�ʡ����g@�t�����BA�h����8�O��*πU ��+����EʜM8#$r��KJ�M�_c��K��{?G3������J�N�	�/���]��au �ˀq�����~�P��b��?�����ha�6�)�E��x�ت6E�܃�6��r�����.�Tf^3v�5+q��3�d�Q�:?b3{_��?�=H�D�%V*K��9�OHL�9����g��V���g/4O<GO"8\9�K�o^��b���� .�*�k����+���_dvE)@	�(�����!~�d:>�^0Q��@!\����bﻍ���e�:�N�����(W�,#��B;s�u�*���䎦�q^�p���	c��k�2ͪ��������
�{���Ҷk���EJ/H3�R���ԝ;(�_�@��a�wf�.-�jʋ\+��|n�
�R�`Ńany2N)(���4v�w<V$K����b�s(��^,q7s�@>��lM�+T'�������+������.�$x��}�=ZX�h檜d.W��MuUɦ��<�U�/1��+��k�����@����#}Q�bºaK�ĭ"��༔d�����;���T=��y�Z��	���GN��Y�(΅�j��:l�Xy��$�"�-UM�OO�!��|���j�qo� [.�j6��S�����K?'����zʮW�H!�h�D_�]����!������$Y�&_�d+M�����	��`
-J.�+�*U�k����Ij��bA��B��B���z�׌��A�O�7t��6�!Z�Lp#�:'�AuM�������ֻXv��.�������U�fk<��^���a��	a4���_�rU�yG6XFo9�F�`��4
��E�9Ѱ�f�r1J���44�z�S��kݟ�[�o!�y�pu�O�x���@+/*j��-RQ�]�v6�1�b�6�����W"��³��ǖA����Tb:����bvH��jZ�
��������92��rԘ� -�YD�Z�&6k�e�$��B�
{
�Kb�3+�~�6�GזD� ��x�~j���.G�)Y6��6�,2�w����n�E\����v��y7ܲ�*f	v�Oe4_a�W<Y.��7���!e���H�P��r����VPGכ���3���.�ņ\q�jq8�J�h��/��(��LL�N���7���\��n
�QE	dq(��bH�p� �r��O��k�u؞�O���U8���=��1��Εt�
ei�ȅM<tB=ô�@��}��p�\�b�gIe�+*��5�=~R{i,o�)����9�Kf�n���!Ӯ����|Ax�J	ଊ��%��İ��	/pU&>�C%���FcV�Li��Z����T��F����������#����m0��֔�'�����0ᗕ��t�b������l�w+NG�U�R�7V��y?}ֺ��Qq���'�ZƢwE&r�����6z�xP��FOA��m�^�?w �j����1�<���as���}����2%�*��1:����V��I$φ��kx�$�-� ���.P�e�Uķь�瓖��`�l$��^�f��>�ܖ�=���	����D=�R?ሲ�I��#�:�+%U)(;��������,.?�2J�.Te��T�*��@�Xy�������Y@�H�/q������<;�WYMg�m7�.�f��vٲ���YMo����%���ق!6!0�~�	���p	�(��cDi԰�����7J.x�\6C�̺˿h>~8H�fN��y���I�D+����볊|�*α�H���B%�N�:�E!�\�Ɔyx8��M5�����8h�v�7�~����A����E2rp��tw�bF̱s��ȴ
�'�߼T<d"�����ڊ1��������6�S���0Y�߮b:���SdwG��|y��|D�����=��f@p������*��Ce�4�E m�6���m�F_w]VJ�z���g"�PK�/Or��:���{(�-rq��-YMf��;^�"1x�����w�0_��~#*��
ޭ)V��B�����c�B4�(�����e�p�?���X#w��v��3m���/|�`~�X>�mC�('ȭE�� O���C�9�{�? �G�kXm����/A�
����M1l���|��|Ɵ�R�<q--%�<ñ�ɥ�ݗ���}�ϙS�%���-.(�u�jĀ���*!�xĺ�w�yr
�a�t ����%8tꓸ�ǻsъ��U[e���<�����<,���E��1�� '�� tjy����	�|ِ!$�wWxt{�$9E*�	�X���u;_i��$�������ReP����	`l_2\�f���TZ8��b��ͣ]s�����_�M�uJB逵�?wր9@���Mr!X\Χm��,���� ��_&�� ��l��\Ƕ���5�8�_,7�<1-&�xP��������f�@S�5� RR�����MN���8[���9g���>�|k` ��)X��^G��4;�ZMog�njr�5IWSI ӆ�{��"��p��c|���=		����^g5�u��R�3*��a��H��^&�ݷ�����i�����a���A��k+Z�^B+��H�U�m�̝��V�9=��]�:"�Ï����߰��PG?�5NOO 6�p�,�sLk��c�s%̹4ы?��^�D�W�ViRy&U'g��f��Py�E�'x�I6:jq���)�0���2�oE�- ���S���A�c�!U�7'�����AM���$?3?T�O�44���jn֝�u^�z�Y�K���4V?��i �'��h�L;P�ZI�
�	eۍ!�+hu3���fE�9+���J�R�j��@�\[��2���[%W<W�ԭ�h��C)�E��?���wg���>N7�8a��ҡ�Ib��C��5�?5�T��^���ǆ�q�����g��"��m=�_$�pΠ��::f=e���7�C�"����o]ZY�����|�4����l���O��o��0½ذD!Y�`��Pd$�BD
*4q�Dpf� �h�O�.'�H3
�F���\Nq�E�bMt�O�A�h�\Na�D�
 ���OT�I��7��nx��c�/����j)�͌u�I�1_��[$R3T�a_�W�C$�����q{�Mk�7}=�y�|��w#l�ě(I�!�%�����ͣcVi�\��5�i�Ma��(�1d���S祡�/����9h��do���~��f�4&$G��q����m8˫V���R��m�pbl�����]�f�6���);���c�+�⊖f�08�w� �����% ������n��3Xp	���{�&��,Cs����M�l��@��H�1J7)jh�$(�"��Z]��ۗ���Ә���Y�Q$꺥ȏ��*Ĩ�@f33AdȒ��`l���lHS�+����D#ҷn�?���@(a���YV����H:O%���_	�4�n�fު2�i��H����\Yw_���uv�8�c�}�3�R)|�M ���	�T.�[�]-�E����țn[���@A�����d���X#��fl���Kb�|BP$�E
y#S@G���	����?/������j�֟|���?��.�q��00 E}���4�(��]F�������ɨ�a~U&7��V�TS�T�LR����D���㼥����].�x��͚+��<_v���.��ݺo���wX��X�Α�gU�EI��}�Ƴ�t�hQT��.%��UR-�"���R`�t�@ 1%�%]CI#�A��Y b�R�<�:�_c=r�P�x�Cw	�&J[5������܋Vmę�1bÿ���w�^�u7�4(���/��n؝=�z�_["�p��ʢT�[�<�܄��x9Ij�����A����_x��}�	n�b�l��Rɨ����K�"�A���^h�n���(�u�/?t�)P5ڜ@�k��'s�"��Fr!���{��o������k�-�f����G>�E��*I7��	�Uޡm�J^哣���S[�he�9G���$�㼭�ǔ6r*b�q�hB~�%���Puxƀ+��Z���@_�j���r�
]�2>�Վ�uH"���8e���`507\�~�L+i���W;Rf���j\���a�%�p0�h��g(�/�q ����������C��o�`�����il�D�-�}4��k9���`@���p�x� �6�ɋ�c����X`�M�~��`� V�P>�&�q�|��J�V�=v�	�h�BU�f��q��pG���ч���j2��v�43PبU9 t��`���:����%+��-���"�=y:�����G�%"��6<tn����i"��~
�%o΅+{K�j����L������/���HH�~��&�\�����_�/����G�J=7��Z����:�v��}�'��w0?��:^�I�KR�v�@�8���2I34�J��p�CP�%����%XJB�\�ϭ��(���bPەE�#�T���I�; 5H�b,4����g,����1��N�N��	�J��Q��y���8k��È�D@�ٰ�]"���K�pH����)ĿO\|c�� �����"L��!OE�D���qB�
9A�dt�R5�hM���j���v�X��bEL�Yh^k�JɩJ�\��ш�QT<���f�֚�������<�Y� �Xj$��\CIp�,xĶ6',�q���}�?�@TT4��+s��tz$��\ ���aV�c>{W9P��>i6
������KQTe�eʬ��w�<O�S�!A����b�ݩA"���2���Z�⤁8!�\���$�oI��㰄��e�_��*�-#�F��t�	H���cİ{��ؗ\��0ߺXГ�o�]|���C���J�e��H\�A�e��9��	�� �M�!+����py=�?gгY�Jؾ��o�0ɨ��i���j'�����,A����1��wk!]h��9��A��$l:ʯ�e*t�'B��3�S����<˨̰�?j��&�6a��겋���b�Q_Ez�P\9�@)�����@Q`X���9�F�+���;([ew� �FԌ 3�d3UA���0�ajUzkY7����-���~���F��KR�#K�'�o�6�W�`��y��ok`~s�!�+(�l���8�	"÷8���B�`k5�f��kZ%^�˄� �t��OE�Y��I��==�����eE��J�:��$��J�L�Bz[�m�?p(g&�<�-o�Erǫ��pIf��lp� �8���|-�7F��x�Rے'�D��yCoD���N�O>����>�ls��<�Z-��u�_Ǣw���|rei��ԍ�M��2 j�"C��C�|�%I�u�"d��D޹�oցA#����eS�^�\��1��e��Pߕ�ބ���@��|;|����!�ϸ����8�/�un�����~f����П���ػ�F+��A�6�K?�t�+H��`��K�k>O�^q�V��Y�y{sW4���r<��MX��	˶�̯5��y�s�R��D�Cq�ϲ�?�H�j�,��О�#	ԟ�:|�6����UO�
�ou>Q	Cq��u�Has���:�:�h�!���b l��J��Iiv:ph��X�Q�Chf���&��-�4HV�3�s���(���t�9���w<i"��Z�5���f�0�
}b"�L9/���cQ-l��R��=�(�עCw^�7�D�S2� �O�ǐD|��qt���?���hu���:Dˆ0��x]fe�a-q#/�8W�5L�ʜJ�(%+�	��������V+�yZzH8ܯ���&����`H4EV;�gE�8��-T����1�)��D
��$�DpI�%,%-�a���,���o��\^�$�>���1q��Jbzt�*������M̳Gt5��B�}��W�٭���c��?L��1�,	��,L�V��O����Va��s~#������T�5�q�\ �����\d�"�� ��¼��Ԉ�z�@
���^l��o���^������ȉ�a��~N��Uz�I�����y�$���DU��]���1\�5(�N�}.S���w��7Yr�Ѵ=��G��Ӎ�0�Dk�tB�6�oj#D�pw�؎󞟹�D1��WB%p�a���@B�Y�$pf�@�/#�D�G5
��"��������q;�Q��*��k��JQQ*q}B�e�Z�u���~Fb��Mq�7���f�$(t礳�3�W��51Ɏ��΁Kx$�-��s���=}C����+R�ҟ�V�H?3���i0WW�ϵ��}Y�S#2�	�c�+c_Y!>��8��J����Հ�S������8�D1�lGc�H�W^k��U�塝wT61:e�(�MV����C�^�p�]�D�A�t�L�]������9&�����ˋ�zhJ-��/�5g��Ĝ�s¿$NK�4	U �����5h�n9��+��K�j����G��Z�[��.����\`���{n�tc/ĸ!i���?�~����/������͑��3~|{:�^(~?_"�˘��Y�7�~�� N�hE�g���@cy��з��[��(�t#��v"R��Z�ev��J�B7�|�k��C��T�]����[W�ڍO=�E�,�$�p�*��]26{L3�P�U�r���7V�i\���݉F��ىXM�:��lu�$�X�Fb9���@��Jϐ���h��尛�쿻~���-�ؗ�yǅ �ʙ�L^�M�He7�j�8�Xt��nJ��16v-�^%F��ө�烄X�=��	tc� 	Lg����ڃxZ��m��$u<,ĭ��լ-�ah�(�ѧCේ�a����Z/�x��J@$gG���pT<7�~�P���#T����GY \��ƽ�Uv��g�Q!�`����~N�/�1o� ���b����^�����5�`%�	��鹄���Yz�W��#\��� 2'�?R�FF�b�KKK�Pʻ�zx�o�U�nE&ʉ� ���0w��v`> �}M���ᓅ(����*8.�m����R����H�E����9�3{E���"��8Ƒ× ߷L|���h�4�M�GT��|hE�W!D_��,���R�"�[ة��L�){A��i�}�?�7",��"Ci �k ���_ʡY����"\�B>.�N~��=�T`�@����Ka��G�d�G��z�'A�6�ݨХ�����Z����"U�n�����+n(9�MіZY>`V�� ��6�=��"��~�_�N˔�B��Įv��5��b�9٫ڋ�HC�q#�_9R�|��f�`�Ž}�G/�t �����od��Ȗ S	��P�n�3xkQ�	4�PV5*��������Tg1��� o�_�лt!��oV̰ܒ^�q���(ұ�f�㬣�;�����W���j��R�0ypW��S��ogO�Ӛ�y<~��㽕v������@KK�yq�B���6�&�9�u]�.Z?9T3��t��ͳ��.�r�C\\�||����m�>�3�h�i�xC1�`#Cs��HqL�p	��s��+�(��EKS���8�r�x���8�R��TJeɤJS�<� @,�b��؁{����ƶ>�?hq�ߏT���4Dp:�Od4�X@�k�2K��þ��X:�@�b�(�_Ghz^��!)���dL���&ځ�����.���p5�&�BB]�	�����·��.�|���T���+`�s	����P	r��B-X"��x��2�*��6֟�O�X���R.�>G�X~BN�H�ʔPA^�*Ƞ��?u��l���;��^�!�8����W��*�{�:��ɍ��@~m�`D/đ���Mdp�����Z0YQ*�0��he4���{�0e}������7�+���r>N����H�D�V�[�+]`�&����&]�1*V�>S�W�V$�J7Ks�J0��r�� nTA%40&�"�x'��@� Z�!�r5��J>[-�*�N���G��	��D��5�X=�P�U���GkH��7��yCD;�o��~�B� 2�Y��sP�|���l/("啣�,j[$��F�8+nd����/5'u�/O������w��2}Պ�W��eI���H�(�ҍ�V&}v�z	qeA�Y``"�!f<�����v��-01�п��$r��Z�O��l���]us�����J+l����ۑ��x��AYC��E������H{i��/\y��?4.ݩ3��Fo����L��U��S�'r�	E��u]� ͟{��:O��/�ûpX����7"�w�E���PR�6b�Vt3 >ƴ�$j�b���JY��S0;�*��V�yb=��-��_n8��	5tI�J�[4H��FH=΄�tN�Av^���_�`B��zZ&s��r=kcd"_�Q%�(�q���K�q������kkk�\Nܿ�:mE��-���w���K�*����ryݞ���7�,D��A��;!p{B���x�>"Jp�	����PB�6��`+#-T5���l�`�/K"��C�D��P�|R���6�4�j��b���Q��%k��h��BHF-��Ta-"ӂ3�Es�D@9�NT��]��_ק����������3qCϙ��*�ܣtW������iHew^xd}6�FS՗���8 N�� V�Ӻ� ����/ ��9d�>3�8��z�,�qD$����F��R������@����ФC̚Q�,c*uUȓ��<��!�#�W|��m��n��?�Fk6�Ay��4�ɍ0�����ϼo���A���#\_����<l��0�%�$j�G�@�T�����]�@N9l`��p<e����t��c��5���G�.�=�ʞ�C�u+D��L��±���{67c;��'wI����&�����3PV���I�C$X~�.Ci��'��;�QuH��2�E�y�s�w{i�
��Ad�wĢF
�����I�����H�Z䀘��It-3zF�k�)���y1�5�`��zBT�k���kp{�a;aW��z)���I�Z��P���YO{�������(��i������'��0����6N~ar��?^���y[�T��ԋ~�z�F6�uH����s�/,�~ '!�*|�HH/�g�C��4�Yg(H�1���\&����gC�3�O���dD�M½���-��c�ћ�v|�D�ȑXM%��h` �H��$3T4���B��Q3{��?$j@��3�Yg��î��f{��?3m^�L�y���|Rn����^�A�J���r=K�
e���18G''��[�B�m�J�Z��������\�NG�����unnn�ڵ� ��,
J�\C���#�i�K���Ĩ���c"���(<)�Ͱ�P�0خ����^xL:��?մY$ٓ7]��=ޜD�y��P����� G$�Y��aN����}��zӢ�E�b���<^ 
&{�Tc�<��/��sy�������~`9f�D�y
��_l0C0'�DJ�R�2<���+י�?4�͗��>�_f��F��0ā�+U�����,{�J����j"s��v��wx>Tfx욙��R|�F ���)8�'�ԈĮǅ���X
7�q��q�+�a�) r�h��s��u�_k%�ϠϢ0�f)S���i���I����%r،�|J���9�@��=ˇOE�kC|7��6H<���Ȉ�ؠ�<(VK%���ZoCV.�
����T7�I���?i��Q��dǼir?�k|n��T*_�a�c��5�O����Z���q��J��E�V��[ �b�fm蒆�j�E�#�x��z���0*-%E�rIkhW�z��{3��O���I�Z6�m�3��㦂N��Z�f�%l<���ec�a�\�2�K�_�O��6.��S�[Q"��r"ޡ�LϺI��n�<�k����El�կ/Ұ,��&�V���3�t�]s�ɕA�B�ݭ3�S.���1����,� ���۲#�~���O��t�F���b�UM��E��.�dE�͵�:��Y@���s����'9�5``���r���_4�<ܬ�OpWH�h��AUj����`�h����{���;V�Z��/���<y;"����Q��%�;�5�o)&,���獩|�	bf�?T.⪜�;]��';{������cN�!�")b�F��e?��5����<�V����j�ۃ1X����[�+�W�<\�-v#�L��r�]���B��煋l�]i�/����#	�#�C���s:�m���U]�?ۥ�n&�"�Ҷ��Li&�a� S&J@0d�)v��y�N�cK�2���R����*M@������^�{O� ������	 A���4	�nf��H}��'i�=���C}Q}4�W�/((pC	�(B'�k̏�����6(��T������ ��pO����2�/�X�p���!+;
�a
���m�I�We�_��O�v��1o�f�DҞ��6�������~�C*�3P�۵]�GE�Ƙ�F��ԙ8&I�o�g�g�Q��g$6K4W�]���ߥ�Jg<���2�A�P�I"��<�D�+�9��ɦ%� ,�s��3�$����S|1�v� � W��6+� �v)�����x��{�^�J��uϣ����a�mG�K"����e�>6�4H>��d@
"��c��Ӂ���m<�,��/BDg��
d��Ök��2��_Y��*�� Ky�j�Cԁ��h88g������N4���0j�7CmO��]������ �����/H�
ʐ 1�J�Z�+��:$.eSU�X��W�ӏT�ev��h-$?d|�:J�~�".����¬�{����
��1�Mܫeڪ��F�A�8��(Ǖȩ�Pꑸ^6�>����#3Ч�fH��Z��˲���o��b����x� �c�U&�aA45�B�}lY}�n(�8�R5�d�'�ߗ��m!�4�g���#�ӆ�R3k��m7~{EX Hd�}§x�h�e��:�z{D���_m��P1�9at]�"���� �pdq��"z@�_�0�%c�Ze�~��yN��GyV*K�لsf�.�ŧ��}��yt�9�b(+W~D%w���uHCB3������v�dM��tn��rc/��wV���Z9��������]��j����eu>�F�;v��\��L����Y*�OH���6_�r����s��ꫴ7���J_Xn^U�9EWܒQ]�륎M_	е\�:�w���%�1��(�w^�ҾΏ�1o(�bA�p��bs=]%��eza�`J�A��`d ۳b�q�u
�;���!�\�5� ���NҜ�8ȋ�{�x��DV~A3P���ǂ{�=����!U:-<�.ulM\�%	Me'��?������ �[5��0�_�g��:���������!�>$ �lVq�%҅P;?�9Ԡ�0�%��XZ�=��8�e�� 4�}i����y�8��(jt�
�5R��FJة����5ؼ��_
ӥ[�NV\�E��T� z�>))b�e�8F��Z�4�/�=o�x�گ�[�b������̻�I�B$�U������� [?h�P���M���u�I[zӁLOaj��5�}�a�@�j3��m!�E�b�\��_|F�v�)X�P��PDB�Ŕ��\́� ���au�Ι��d|�7��P�.lL�P	kRP����m�o��ٶ�tVޤ���w���ϧ����(QYv%&#&�% ��	|���Q#�ľj�u��p��2��е�AF^~PD���n�~����O�5B�F��,�K_A�f��H���sW����V�on5�L���{ܯ����9�5F��-{R��HbV�Xq����--�8t�%��#����f���2z��݌�l[m���:讇�*�F��Й��D�jk�̘h����O�L�����D���v��_�vu��@�g+�C՛�>��w���f�I ,��W$|.�~Io�V�-�	1��	_�a���ɫ0%/��g���䛀]SV�3ǯ�F���l������\=�:���r�y��;�wå�?P���VE��'�f�>�uV4�ޤ	JKK�Zۯ�ߔ'�M�=��Ւ��_� ��������1p&�\9���{7	��X�������@��I�.��+숉,�����hX�'a���əb�ƞ�2���'�^��ò̄$I1a��CU�^�_�IT�zH�m'��rR+�Vv�3�_�B!A��!S��������nrŉ[t~O�D���ރ�c#��	��q�zA����w�����<�Y{XԼ?e�7��4Of�tv�b�;[z�o�5�8Q\G�ĥ�6�go�'�̖�IG�O,��4�;�H0��% �S�o�}��)T����UF"(%s�8ƪ�f��0�c��"OaH��F��qA���h�U&���v�,�P���U{IN�!KZ�'��I��V̊y�7���eTgjSO'4?a~n�q�gaڭ� �W������u���+�x�ELFX������m�l���x>1��O�8,j����M�J���9�����M$��������������ٳ��ғ��3�_;|c��;;�ݯDwc��Jz�;9��c��H�N��XCLp����M�b��n�����M �j5���cS�����L}ʒޘ�窔�"�s�b�Ӟ�wFT�*>�y�=y ��dS�'�~�R�6ZGr����K�~2����1�+�\�6�gd�?g�`o�"�^M)ܠ��1���q3��W?�D�?ٹ��ɦ�}Υ_���Ȩ�t�~a=#,�O0鰋�U���3䰄ʧ5�S�)4�1C�V-��$�r����I�v�=���f36eg����p�|�_v/�Ic�WăH��6+��xhsE�Vk�;� ֫�A�.����y�>��Ro�mZ�܉O�x%C�5��-�P���_M���O��{�>��>��3o�(ՃV�#�\�6��\Q�?m^�h0%��a�[����dBZ��y�b���S&ꛚ.V�<0�w������ѹk+_��u�v8�z������g(Tİ	�X�s�Y;	���j K�j��A�K��1�_�*$R$h��a'd$!?M �!�:nz�I
���+�vS�������9���Ð$T�����>j�P�Y_��VG�꿜��?=���O��gEhT�w�0?�u:�u���[͗nZ_qSP�����J�������Х�i:^_?����'ۦ��Qj��� ���p�F�����3@*�n(���.S��$ ��#�e�T����f�{L����?���7�ze�f���ST3?�/���y��sM���_:��J!�g�\A^��oP�B���T�c�,��l	�7I1>[�\����� (5F��?��v�,���o�V,��������<�v9�s��8M�AJ�����"�hc�1V�/}��-�i�
Ee�_��9�A���p{���N3x}y���6�Bs�=f�����4<c����
��
R�S�5ʢ=�P�,�#_O&�9�=����>yyw�R�Q<���tzA��L�}��V�V�@c .�t
�fE���ʮ&��m��U�9�-ߺ1�Hm���\���醌_�.�P ���� �!��A�5�MQ:��aԞ���.ǋ'(e�������U/���]@��́�=< ��+T+1D2at>��N�d��Ĭ �lkbJ���%�).T޵���|�Lth�$w��R�D,�lJ�� 5��AU_��V��k��Cֻ�Y��#3�Ǒ�II߈�WX�?Jp=�P�0I������E���-$��t'=i#�l��}W����f�̦5�ͥE�<AF� �Y{[E�y�G�]�ص"�mBr��ro����细�yp��t��o��ȗ�mNX�VI~&��`#lx�1&UwB$����.&HAe4�A5�Ɓ�^UG-}'m7�5!����� ��W��������h�Xg.���]���:20���0���*1~ly�P��
r��:��P�s�/�«��Q��#��$5������Y�Ų|��.s�.6!ϓ��0�����H�,�ߜ٭!�%>���u��)oYR8b�k�z��!w�D?Q~@rǊ1�&��S��^�=�Ut�ʝ���!�s[��y{�s��٤W��K�=����<�w)�Đ�!��!d�>I2x� �u]6���Wǣ�&>��ay�����sOsp�2�w��\V�ANg���E�wF�4O���[mI�8����[PU�V�+�3�%�T�/��E��τ����z���}%���H���Z�����O�=������o���<|T�)R�cC'V&�J�fQl�ￖt"ga����w�}��ɸb�����K� j�d���Rv��&�:ܒ4�j��Y�]��4}S�Le�����J��Q�Zz��D�o��L��{�!Į�\���ġ�����z���ρOb����z��'���zZ�=]��a>T/�����������~��:[� ���O	bU�+N1�6���ym�I�i�@DkB��S���O�+�i����=`�]�I�C����\=j�����r���co�<�ǟE��)��3�,<�"% �W�"�gN��E��|��:��*O�<ó(0*H�����J�8�~z��@j"��#�Tȑ[8��"���#\�
J��^��A���P���J��h|��F���9�͓�"+]�?� �e�؀X�����Nf��֖�_w�(�m-��8�)<��F$LN�#�UV�a]�4EۊT>�z��__YUZgUŽ�Ũج#��^���o�M�	
�A�Cd
q��Yݬg��,f?P����k]�ך�����љH>�Y�ӕ!��K손ݫ�Z�t�Xb�7����� �s]aH���#Ž�B@���n��`T�-�y��m�$ٱ�2�6��qo�%�ؤ�2@sd%��	��9�K��uA�u�P<;�|�6!�|jR��È(��[�x~��	�f���Mn�'D#���#k�	��T7��~�$Q+�腭(�iq2f���P<�����2v�<g��g�����1�ߓ��Ԉ5p��e.�ME3����i}mR1���i)eR�4Y��</[W��5�!հO�-�ol�T��x�� T���[p��4�rC�V�{Ո��>����J]�ß�^08?��F#zx����z�{�B	��L�bs7˨2�ٗ�?M�����c�fQ��G��^�󄴾ЋA�y �j#Q~�|kMm����7���버�5��\U����m��aUc�������ex��	�U�,��\ɛ�v��t����f�ڰ/ST��mA��1��g�|y��0���M-�n����&���L'��ri���g
�-Ceeex���]+��:kj��!��2	ic�8�88��y���v��e���j0��\}b�����
����H䍁��b�B���Ҕ'��_��)�-�^n��^7`�-:.'�cV�e���g��tCb�7��5��������u\���Z�M �)�-`�L<��c1�paU��ӌx.�o:�a@O2�\�{~o������qUk��$bƆ�+�����朆�fb%�Xe�S���7���oN����M�����L}[�A8Ze�Z*&�x4�E�$���S��;MSy��p`"����)�� ��|�B)�R`�X�y@��.����w�(�unmg�߮g뺢;=�3����]�A't�U�ϽmU�4UQ" �?0j����haz��`�=��H3�N�h��p�߶"6����*��i|4��W��.6���b�n��\{����p���
|�X' ;�.'��/Rj�o-�Ca���Rܢ�֪^�%B(L��k��У���`�|�\�8�@gũ�-
�,�j����e%�&n�s�Ľ2-��}ێZy�Ql�>��12��8(�z�e]��B�m[�c&�ۼ@�'(4�Y�Nƾ���JX�ȗ��Dt2ө~[G|N���}������o���l�o:��J�O�] �� \o��ָN� i�dJ�VlUlRя���DYQ�hbQ�պ����^����+. ����]��?(��3��Cl��(�!�:����w�o��Q����u�w��s�y5�-��1�?�������м���E���U���o��%�lX �{*䉵����7�-l�@5�3���ٍa����;�:Z�h��c���n�:��A���������9 �t�|�C�-� �M6+�(Ա������T���T���
�J�#X��L�b�F��z��B���LI��t�.�[�YwM"	����t<��E���c����Y�N�#X M �T�`��z���;'K��zM�L}���yy���b�����7�dBX6��h�
[�f�����=��Po�uݮ��~(���.�qC�4���i K���	��g,��r�}����O���}��w�ƅ���=8��fzQ�n�<�@�C�.��bƉ�l@H�QãIm�1v�չNە�b2���!�z��$��Qa�B���y5���2���X9��D��<o� ��-�;Ziy�D>g����8�c��4�����5��f��Cs���Ej��V�.�7$�b�PU��`�Q����NR�2_�B߃E&B�z���y��w����?�\�M��]�g�G;�@��n��:�"wR)--��\���5L1���Q��O�S�TL�n��hw�V*i�K�t��#O���&������x�%��<|B����h^��J ��L{Ǳ^�*��'q�ЧQ�g����17�5�&EY%���m�x�\fa�|j��v������?���P�L]8+"V�손U-1 Z�
�p�/D��k�.vU�u��]o�t�\K�s'�H+˼�v�~d�����c��z&g��
fDaNH.�읙Ae��D��A��!z���-��[G�Q�%�vf�E���\��(���<���Yk:Z�!2�����͙e�\��9��E�%�6]|�,Jv�4��kƙ�9�V�q.�E:��o�5�r��f��y� �d�;Q5��d��/v�e�� �'}}�׉bżF�����7��m�]�I�����Å���#���NMO�r��s$T���du�$�N)Z�ڇ��k{��@CQQ7�$�Y19���r�H@F��C��2��j	dp�h�!)��w���ݬ�q@z��!�'��y�ޢ��by2�+������J�2�/�7��/���s��C���3��-��� #}�T��\]��~��C	s���)��b�r���KG�; w�t���q��t��z�����gvE4� 9>��|���o"��g�K�T.S@�&�4��b��1�=az��#�"I���RpK)�Ib8�ᒓ��*u%Y�*l�])�t�E���$��G�yP�p���dC�E,LE����p.���\��M��g����>��>�ӹN��5`�]�I��Ϙn�i��褁�Si�wF؅�x,�x"V��/�2HY-����B�<���w0��o���3q���?-�W(�n��eTG"��Ԥ�ϺX¡�P���"G�>�XH����h/�2ԽDo4��Ȇ���@[C�J䇬:��6�<�9!�PFl�]�3��	l��]�biR5Ґ�%�2��p�n�5:���1Ǯ�?�<�_�e���Vb��O]F��@$�4s�2��yƉ!��L `&34�܏�`Y?u���%`�*�������q�ӿَ�7,��Z��:��'��!��}ix��!�"���`eLk7^7{T�+Iy
��U�֬=�6��4�����,)�*��tH��H�{�}���|���Z$B������9���~	�<���Ф05��^�D�w�Zj���٭�:s��I�]�$v��?��ء+-�����a������*��Ҵ��'��
GV��r]�� j^��hZX�_�����~��|z��o:�������v����+@�zA*�0�h:��Z:�*ډ�i a��
���Z�#��m�A���u���y��T8(F�j5��ح�8 8��k�Px���݅x��3k���@�o�C96���7yQ9��:f�P1�j��(Ӛ�
r�H|pEN�1񸨒��T˵��pʆ��(e�Dvh�1D�����z��b���3x��
�1�]�C��19@�͇�*���ޟ�J^W���ϊ�����'�9|Ņr���/ϭc�R顔B�]�fДp1�(�S$��-]���2�H�?�"�#���W�(�;�ܒ�qm�����<j�+�?�+i�Q���/��/��������,��N��g?=6�:�Vr�6��n��@��]��>kW�#�$}7��6�BS�Ə,+&%� �'*�W��kv>R��8�ZO.�~Z8L�w&����@OVt��V�rD����w�W�}���p }�.!� "XV�X�"(�Ng��i������Џ����-V..ǒ����O̢�jEC���"�����_��N����d[�W�?_/4�U�+M�����X�D[��(JV)�'�Q2�
���r��O|8G~����5A~�f���$C�6��l�r�$2����%�w��ܮ�2�� �I�ő��3��������W9�`�Tc�ZF�U��HI�ź�瓃'��BM�A����_�$LR��C���d�d�/�����c��6q�Kv�,�ù6Lg�� .�^�߿���n��_�q�	��?�:M�$3�s����א�B1fԖ�����Hwh}�Xe+�2=N7�*�`zJ�C���/���|�|�\�/~�KԹu�_��wl�
}�����9a
�i���>���:�s��h���y�&���i��	W�T[�!�a��I�1 �h��uw��ʎ��d�#�8�<>N�M��5{���n��6��R<R/�����'��,���m.�T��r��X�����v�Ffsh$�|C��o%o��'#�e�<��]�)'�~���%Ek��̆��bP�H=�3aN	a���z>�g�#s`�}��'C���������*�;I6���;��D66<Q%���Yb�&�:-�Y$ 4���<���Nl+�Ģ#%q{}g�YS��2���������*�-�"��ϐ��v$���,S/���*k�[� �&Q�R�IP���HC=�h�&Lj`����RnVÐB�BQS�#�#Ed�� �[��]	�z��!��S�yR�|�D�Lh&]?��&sf���fD�B�.?/+�Z��|�©;�_�L�YBű��3�'�*[�B��1	��8qN(�V2����4	�I�!��IX�w*�����H�w�S^@_(�&K�qT�X�A(In�r�O$ @P{��a��u4|?Y�+�B���:]DRi�O8T��	MK1g�D i?��լ��ǆ���~��I&�>�vQ�� �U���=��`�2�E�yU	��\��Rm�ae&���jz�}��p:����N y =?�e�����q^o��-������n�&���@�c�]��ؖ��� %!W)�D��%t��f7�t9��t���b���Rf��I�W�0%_�,�D��d痴��0�ɹ%��Z[�f��Tt/����X��P'Wח���k� ��_����m�ş��ˇ���
}5�4��;�x�Y5�Rʺ�~�Ѽ�^�k�+��r}���wrp�O�M��ҏ�A��QqY��j�s��M�����$%���h�E���k��aV�ʚ�����9-���^�׈����t�$g�K,�Cd���i�3�+s�=--2r�)1<��a!Y@F:H,����s�Q�ΐ����c3�n��pS�� �!���Ԡpnv�Dba����".u��#���g�ͣ:�����b��I ��:a�܎�Y�f�
�D�on�r9����%��[�e��h%~`����꙳܃nZ}�;^r�u�F�y]���|<E��u �*�y��s������k�>~��/nb:
tO�%E�����
���/Z���S`�����BjhP�����C@e@�n������{�{�O8�|g����Z3�ٸEL����=���"���N \�^����l�R���'2w 2�	����R��zq�L�\r���%�*A<��������Y;2��J{��m��5���^6{�6�p�.���4Z�s���
t�;́��6`��1��(���p���ܚz�,\����+E	&i��(��/F.�����)^9U�������\?����Wݝ�������O���
+����̽��`�W�I5
���4�՘���������ӻ�k�3�������1��.��0P:�wԓ�;I��o���Iwx�4`��s`"�_�ap:y���],��Kj���.���1U��݊��?��-��2�����t�Q|����Ar��3�ӵ�`���"��=�R%X}*��̴�c���b�5�{��4��(��~죢Y���g����FV@�h��Byq6�?���C^�7��+M#�Pr��j�%#�������*����̑=��Vp��Ӑ��,�12%��ӣ����m���i�_��k���B�
/U�l�����~k�k?]|[�
����L��MΓD�r=�[��`{=F�\��]_�;(�C�jڐ�eD!U<5��|Ç�������ɖ�?k w�KQ�	���������h�2o|-z�x��GaR��v��lQ��MM��PR���`�f�ճZ���0Rҕ�fRz��Kq.�Θ�~t73<�O#��:���p�O ���p��r&�)��)U�G,�r���4�V�d�;�e��Zb�*-�}@jk�%�7�9����*�j�i{�:��������UKڢ��X{Jl�%`�|�������y�0�tK�[
����Ӯ)��.C�A�xZ2�ˆ��D/z�������O�q��)���b��B�d:i�5��3�<����D��~�E����_X���#N�G�0n*�CRʤ/~-'9>D���]��.�Dm�Bx^5;oS"���2a5#���,�����:6R�����8C�=��L����讞m®�0_��=��L_���ui�(�Oa�G�|*�;Vއ��lL"q�I����������3�(,�M?��D���]H�~��]p)Oȁ��������JyU�U[�.��o,�~ä3���S�@�<�9��sM2:��Hi���"����0�s�b��r./ʇ�I�����}9�� �)a?&�����z�0�P��8z�u�]�����&���5��Ԙ��5އyrBw7���������ᣥ��1q:h�?dE~�T� jL-,��o��G��{��m�Aj�Yn8i��a��, ��X�36d���h^��F�'���o��v�,�_��Rj�wX�tI�if�D�f?l��m�Xx�����$���2�7%��~���~hr.�i���O�Pއp��G�`�-�-�J���'���(�ڰͲ4�g3��[����a�0}��E�N�<�f��2j���JI����u�c�{&ȫH�8;nY@$�eX3=gP5;ӂ�Σ�bۯ���s}`�u�zR�����MX2نiAK�i�0����[�O��G�A���Ƣo�>Il��r�D���sK�������m��yB6�L;>���$��e���k���+�<�O
5v#QhS�㰲w-�B���~�{ ���j����O������p�=�-3p���dm۟�=EHM'��\G�tg���aym�61�Ϛo�ȼ�R�X��ǯ1E�U� A_�2��5��q�S���Aj\g3k!�1z �c�<�%2�oM�'�Ҁ ^ZmX�Xt�\]�UQU�R�k:�µ
`����]���(eS����BQg�6���`��>�}�Y_����bQ��0VҺ����s
�2�Z�z���r:,�.G��_�C
�q��5�b�������g��*m@�b�ۉ����M#����Gw� M�s&�Y������4?����/Sv�j�Ȗ�Q��5�ׅ�w��r��jd^�p~M7O2[572��lz|��26�Dz]0����!h�CV��xy}b�*1,5�_P�,�� \�͸a�-M��Ʌel���~?��D �N����
l����D���I)����{��l�	�u��-�C�T���1|}HR�I�3&&�D&'q��bG^V.7������D�3�)��[HeN����߁�Z��J�Ĵ�2��T4��K��p����-I�y&��`s����o�Ȯ����A~kGPNoX
�O7#���-��ϧW��B�e�¹F(��"@�7�VJ��S4��^!���2��f��C��s:ۄy=措�i+�B�8{?��+�7�wCDQ�q�o�?$��a'�V���4ĊO�&! �M��s��ø����'�>��.u\hh>�r��׸6��oa"�-��a��Fn���z;9yh�H�Q���J��I�}K�xƇZ':��a����c��dk>�� N�qz�4u,.Yb��91��K=Ai8,Us��/}}j*�����%��s�����Տ�1���M��w�R����~�t���'�Cy�V��;U`Iz�qm����r$qG�O��o^���6���iH�6M��MW����U���$X�#*'�A2_�0x�Y}M4��FrP,�s�����O���6�.�N�7�@�te��T��p��e>�Sկ�����G_nl�Wu�1rٟ�9^������,�M%�^��K݋�o8>8��w�����9n��F�$d[�gd� ,�St{�˞��Q5�t���pԞ��0�`+�0��h���6�I;v�����G�{F���Q�[��6X��~z��~�+�[ۿ/T��(��Z�2&��G����6�U*�4't������ݘL���Y"�41�B\N�����ք&�7u���D[e_�Qoŏ�Ƭ/��C� ��;��+\�߃D#�H���D����4���A�$�(�]w�	1j�S3�,qT��j+:�~��u��6}��l�,�5��k�\�>i�~_����D���o��Sȼ�u>�!IJ�<uK�Qy��l�Iuuu�(Yh�J��ߘ@��}ēh~�44��f�K��m�{[XVF&��]���)`����b6l�k|�J�A��G�폯G����W�&��X�`)��`|���L~�hC��T�W�g�}�E��8�F�|��h2r��0W���n��y�c`�>��
�-$�uܱ4���%#��р��ZJ��\\�'�>� 7vw��۟�
$��p8 �N���W�TL�o@�f�����h�?*׵�,Ae����vMP��V�>�T�$G@j ��"���m*Y�E��A��ӎ��M��6�fF�엀R��޲޼z��?��~g�!����K�W���զ��^6��H?����1$$��a��@,.�!n?0(���,չ.���P,񳼲����]dЅ�cMS�=�X$���ø��`��4��w���k;�o	|�ZK�og��"�7&�9�KZ/�dN	h���e��+2�h�������8�k�Qׄ�z���gD���	_�`��0�ĄŠ��X��/4��/�*��';S(���!�`��:k�jx���nX�YN~g�I�Bs�hnMc���^�b*����y�ﭕY����B�U�DIǁ��9̯EC�a#Az�>�R�ؾ_\��w�&��.U�?J��!�(�[Նx��A���O��=�L!�,xw�D/K988�u~����>�_ymz}Y(�Sy��K������{�z<�}lĮ��A0.�kC%�	Y+��q^P����!!y~�J
�w~�nĴ�ޙ�6�_|}�֖��&�¼nȋ�<�����<	y�����~H�����J�b�]�{����Fq�����󋞽�3lXN��O�0`+8Ynű�S�p�{��7��,iب͚Cu�)R�g�ls��e�ʱ\%i�s��+��a��k�$F7J�c�r�	����� ^���	s*˚A���.�a��p#6�\4&�P�ТL%�MaM`���OF�kd�N�}��K�$��x�2`�l}����䱂�%�7k[��o��C5���15~l[jIH�m�`i�k�&�L���PL���G��b�Q"g�ɜ��k���@�e/�S[��6 ܴ��ё*�qS���aйSJ�����'�E-�п�	/�o�(x�(���^VT=�ҧ$I�? �.���`���֩"&�e:y��2[a�h�sj"7l��NB�G乑������k���;�NK3_�Wʆ/x�e BH"#̅�J�~1(B����L_BQ1]1�]Yu��.�p�}�����CZ+
��rv)o�a� �f�������^��/�Z����qU;վ�?,B���w�R��Й�T�ڒr]��0�������"��g���g�p�3�mj�
z�����~:�\�O��.�׾��,��Fl�c�T�㠩G�@v/��~�B�D^�G~�Oָ S?��[�|)�qKTxÑ�g��h�� ��؁�+����_˅p	��U���N{@tA:� [j�x��:�x�y�2~O	��W8�s�^�+��^��Մ�W`��n��j*��<ZqȐ�Z��Cz6�e�#��~~~smz�v����X���l|�]Řj��,㦭m~�t<h�u��o�M�G���/)�p�$&!k�Gj.�h��<�ɤ 8|���Y8��5���΋h��i������\�\�� �'�^���rd�?��~�XbD��0�X�!?�ڲ�38��Әt�f�"�S`�}���L��*���?D���i��Ul�!k��_7�D�wf�2� ����'����QjA���t�\��-[�<�|w<7hF4|����~v�H���$�Us&�jB��4��'_i��Wˈ��NvL�c	��^�n��J�jg�Z��������m`rl1!�y|�A����3���%jH��$i���M�+������7��W^��O/5ۿF�s]<��~uc��_��RBa�Ͳއ�v�]�䶻TZ1lxf���s�O|~����.��j�f:�g�Vd'�ij��È;� �N?`�f�gD@_�ֺb2?����!qA,�ȍFP7q�E0U�Ї+�\&����*���EH��ቩi�Tk85C�Fd;�H���>9�<��b7�]���Zm��Н�Cܐ
�C� ��O����`�+�+��(<�4(Ci�NVV4���\�5-Oi| ���N���5����)ܖ��G��EokN���V���R\���):w�<!��T�idm;?�E���jp���B��d����aH��]��zlk��k�tI�eA�B�g�r�I���kj!�R^���C�FQ���r�8y���k�z��_�! %A�-/���L�,�sL5?����**$�mY\`�$��Q�5ԞT�є���b�˨0Mq7ɇ�D�`��=�w]DX�������,�l�!��2lw<�s\u��ӁԀ�+V�:C��.�L5Aԣ͢�L �xě[�U�?��mH�	�����}���Y�dާt�I.�$�W��Z�����,1�����u�`�p;Jf���f��a�"c
��W8鐼�y3jy��K�g����E
���n���X��R�×Ӿ,��ɦv+Sc�Ɲ��y+�����U��f�'F#�Uv-���%aF�N�y֜P�B���
|�:�X��V����Ȗ�}?|pص�)e �4wIj6j
u���;�<}4a'm�� Rz����9!�[�(R��d��/3�i��ok���	�F ����m����ꏩ�bX�h��U�r+/ 3�Ԥ�`�0���9�\v� ��9��昖�9��7��5ƏI!������1nlћ`>l�3Va
�������:����%����|Y8B�X�jB��HH-��ǏV6�]�M!�NX<Cw�1�J����E��v �a����[ު�bLW�c]�=w�ftQ�'���ش��(�w�Ӎ1��VT����F!��|�hH%ӗ��LͱAgSU�����vo.5�E�_� Z�j�]���>y�V����0,�X����c	�3���i��c2�z�D]N&r�`".�F?��F�����Թ��a�kE�a4Vî�?�W�̅�����$���}��$ɡ�P��U����N�
WB�*�|x^�M[�s7�9�dQ(�	�٩�E��7����ZB��'�W�q�D}&�90F�3{����!cHF>�H;���Q��D�4�pI��	�Q��r�a���gح�Xu�c8T� 4�X�7k��pȇ}�猪͡�Τ'��~Y�Cb�BL���XI�V�F0�ϳ�b��lÚ�~[�A�%�؝�,m^�_!�����
�5��)�Y����{�/��&#����U�y��V2��k�@	�\�'��=�BӔ��&��zi@���W~٦���I�9N�^��oR�a�JۗJ�l��"
r�����_(�	����`M��&�.����?\F|���)6�ja�s�y��"���S�ZO��䜫�&�n�Ȉ�}�/�y��Sr�:��߽��[��w�K����$� ���+'A��Qy3� M�E���}�mZ�K���Q�,:��gO��[�T��|D����(l0�<w�~]#�K�9>4&m1vY��1=�.qNz�H��*V�����ګJ�ð\��_2^US�W�^]�"���?L��z�I)X�-�-���ө�`}D��3~G�x�_z�v\M�*L����ձ�MS��A���.��QGE�s��%�v*������rEc��Qh���1�������P�~Ԉ%G>���6*��"4��%.�ᆀ�{D;��/�pB�]�� �|س{ɚ�\TT�\o��v ��zdN��b�1�or�����;Qz���Y���6}��ە�5?#��vK�9��lX4y��šMu!�ڶt���p��4��R�ž�����Q�-���)U�~3�:q/��[D+��P�U�Zt_b�dQ:u�f��dD�kd�����֫T�K��F�m�>lo��q:�Bv�b���Ty��}?�Yu����c��Ь�|��}S�ώ>�N�Z*����P�1;w��,l��ґ�ns��x2[�g�����Z��2�-�)"�|�:3u���٫W��&���&5���1�M\�� �9}j�.N�&�XOlܴ�6Ѣ�t�����
�b���}.iA6��m����QWd���{�'�V�t�>2��M.
�#J2&��\+�}���_�k�,O4�\�<�U�8�x�H��Kiu����fi��g���Nk|����m��o�k�
�#�t��n�� �cҾ�P\TFAM�E�Q�̳��!�ϋ����b�y1v�����J���:&�=Lt\�����5 �J�y���g�����ș�8��O����9������1�4: ��Q}�V�f"�xL�V!ڜ�	��NF[E.i��/��[X�fJ�b����v^��B����4߸$5�u/�ı߃�����a�$_8L���z~d[m�0M�iQ���| ew�����s�!�[��8��e'��?Ɏ��ɏ\��}�_���Md3<"���p$��@Y���>�� -l��APE,Q�>ch���8���e�s=��.4�୬�5�v�i3�v��|L!�JK�Qz�f�TmXc�w��ى�h�����mYO�����;���
V:x�jS6�j1zlћ�SA1�;#-� v�RmJ��%���ᶃ� ӌ�����T�?E���W����b���K�ſ
��(L�ϓeH��Za�?����{��h�M�)<�5����mo��,U�gԢb���bx-�Y��K]Zۧ�yF�2��Q�+c��-L�q���f����<Y����9>��˱�<��H2���l�x�(�M���ζV��JeT��vj ���S�}á�U�;�h*� �����K��h��� �e��lq��0�D�p�OT|����r�t��"�[�B�V������!UiSg�eޥ-�LR���||�܅x�Z/�f)�j�q�W��P�FX�ʠdRp�8�����BE.$�6��E��mb��D��ЕXf_Ȉw�gjP�� ��t�>�:�:]^:V��z/x���@���h1�BB�fBv^�����d�q�
��$��`��ا�2
���W�����r�w�Ŝ�7��<���ˮYk��G�ۢqY�4>��i�Y�E�A�A1I����F�ZU�{�^�˫�����
b��7;���=��͒&3��	�Zv�o]-�7����q��i6Y�� � �	�S�>���-C�}`h�37�g'#��yߙ�RaC_���F����1D�e7����#�u��A�dp�	e��/(}3��^�?4&�����~��δ�,iwϟ����K���&�8�b8���`k�UT��2!J��u��ةG�ժ}kPv��J�sE)�	�[�^�+%�O=�:�1�L��i�Ch�|���P�$�g%ђ��I�+�4RJ 3}�D���O�OQ�_�g�辵�����'��Eu_��2�a��5�f�[�����h�5�p$��ŷ�ꇞ��,������%�&���Gw/�@Q#:W�q�?#�N�Uz�(/�S�Δ(w"��rѰ��	�������P7ψ7�D:�pE����'ԁ�T���=�n�Kh�f��ȳ����X�!l���FT�����f�ᕊ�-�?�"�'��P}�~o�p8:@�e�/5s���t��%i��o&���I[lrbH��o��
o_�O~����8r��<�묐��Qמ`����ook�[���U��P��w@S{IrK�x��j�᱖��5ꑩ�{�ZLvL��K����nc?Ky~
�D��M���Aȯ��!�
Y���������e��U�,=b���0 K�r{�{�z'ܰn����QK��c-Hl��=m{(�EY��@�Z�$	��=�R�cT�#`�m��a����yBo��I)�M��
���?ۊ��|�F���0L�TQ�7�1P'���1����2G�����z�Na����,�C���d���,�����}�J�㰫���&��,Ɋ9o߁%os��Q"Xb��`t1�����+�v�M������L�R)`協���!��K5���Λ����@Uz�q�9�CG��ɸ�ҁq4���yZ �Y�A/'��������	j%Ώ\&������Zi�ϊ��Uǭ���9��W=�jW��<$����n])Id2�%����3E!�1Q}�W�"
M
J]��ss�?�@�\���Es-/�����������W8)�������aCl���=�H�3�S����z��(�C�k�?�U�V��O˖p�Њ���z�k������I� v�W�z���%��+1ʞ:� ���v�᫆��V)p���D;�{ݼO�,�M����#���Q�(XCC���E=���e��,Aӈ�m��;h\��7�Gk�[ʹ����Sf�}'	�����ݽ3�R�7�!�3�^�]kЇdEl]�J�:e�6Vݪ6�Z�
	���d�B`
�����Wwܸ�u4�D!V�Œ�m�n�tnfo�N������|\��E �-���)tU�̤0<�`��'j(����:�0��!g�2;X�����wԵ:T�6��5�^���҉��I믮�%���#�:V��3�(0��_��Y/�.�r
;��Ⲩ����B��q���5�f6���ñ�Y(F�j+�M�7�>Ӧpa�no�^z���sM���@h��~pi�Y �n�-	x^�N%��SS��JJ�L���߹�7��{�@�`1�Ԃ?�D��M7L�8���A�9o�E�j
�0�Tܗ$�UˤxN���8�ݟ<�g1q�nZ��rL�_�G�C2��dvy�TY��R�7�`s��hv���Џ�>TΒ2f#Ǚ�Ŋ��&�H������/��t�Ɉ�2�p�����6���z�DE��s���a`��^�x�n���a��#���P�<��}~�9����0����O�pK�1oJ��F%E;gK��f�e�SO�/;ף_}>�\y�����<=���l�؂�X���u�6�����t�rɿ��㍓"x_��/{9����>��"���]h��˸���uJm�"U��Ta�^&b��\��0���۾�-���$>^�7XD�� d����-�R��	��ǂ��4@���Wq|O"4�%v"�^�skm}��i�R!���y[�!,4b�l��{P6��W)����U�񞣺�:��t���훺D��ieGtMF`�.q}[�P 3+ά��dh�P]S�wX#Q��a<%o��\��U��B��^J�7�]ߡ��hm��F��T�/Ɋ�ŉ���-�,6X	2����ip=Sɳ;T�UUi���g/Y9v��H����H�9��W���~-`jI�{�ݭ?��a�)VB��g`�Aڱf/|���L�׊��(#I��T$�_"�؟cj�z��y�\��m�^u�,K��`�Ċ"�tY_h�#�c�oR]�S[w�.2���wx+r�fu��;?&��_°K���R���Nw�آ��	��� �O��|@8+b���Ƥfi/0�ֲ;���>��𝸌��_=�����p�Ҵ�U�.`��{6e���|��t:.�NSx�Z ö��z�M��%�\��r���f_���K2P�I��}Kʶz�S�k@��R�ķT*��g��"�V,��"�$9�E+��و3����mߣH����zA�ҒP�n��GǙ!	�+��>��뉈Ph�8��,h�������"T���ĝ4w��,���0�`�=��S.�h&�毊~l�� #I1�95�sq�
��\�m4���/��b�	Dʺ�åa��*Wm�4�+�4�ؘ³�sY$?W�YV;m=��;� �>"Q�Ũ�����7i�F:�b�O��,�7���D�xj�r;P3�F�􈖄
��Kp4"�3鲰���ݥ���k{v�ې��(��W�S�,�u�c��k:J�������a���-) �Kțj]�Lb��,�	N�P�e�$�����~�\�����Q���9Mg?�2e��H#@q#��,�Ӛl
���	N2]A50�TX��W�L8E �B�<��׽/�19��n��s ���^���H*/���a��t"��P9�ݟk]�����`4y�7���#�#Zٻ�8"_�l�-�:M6IƯ?���[����d����y�.����R��3'�BY)�L7���|T�ӈj渍��`@-U�cJ�UJ�[2�j2u��؆/�.��Y~�����Af�;��j1\f؊iׯ���l̢`.�D\��ӡ.w������/�{���<lp�ΙU��j�����
.�b����0���3D/S(cd�&'[6V�Mie]�,p%��M�E<]��k����fR"�c�!�.�d�rZo�Ѵ�s��N�o�[��}L���2��e@�6dP��G���f�e�� �����G_X��?%.e�x@�v7�a!��x���߄J�J��|����xpz��q�K?�Bz��cs��y�X�@��YO���	�aIQb�Qȓ��� 	��͆Bf<�`? �N�����u�Yc�Yp���*�������3�\d�kcX	��)YZj{�-��+�!��I��e�{h�'q�@��֒�q�g*䂧�I���ڎP �{sP@W?:�yx�����!��[��W�/���Y<�yྴP3�ߪ��
��J�x�����j���?���m�P�n�v_C�x����/l��i@}{��Z�o�IZ�Gj�+룐^��z+�]�bRn��7.�q3(�!�ĕ��@ܱB��7�\����>���eV-��7(�O�`R�wy�H��� )>��&f��t��#Ӣ'���p.�/]��4�pΏ/t߶M�V��L�7��R+��(7	+�IU`�}Y����I�^W]����J��C0U+�n�
��؄�2�c�r!9N�k��&�����1�W�_�:�~���'�+&Ҕ���%�z�"V
)~�2�c��QS�6;�]��y$�j�Zfv��4�,�x*nS����'���Q~�N̲�ߠ=�������;dfu4篖^����AaH�>�_B�����9q�'�2�R�1�/|3��K�˰��'����b+|g�ЪWr����`���WY��L	���~�ʾ��~IT^J�	�,���l&:(���}od�Ԭ��c����n��u1|މ�T�q�M���I�zO��F�GD��?�H7��FIs��;�dw����c�N��RG���@ՠ`QF�v��̏p^'�x{3$
Ʌ�/*�A2��AH&�^��?�@�svJx*a��(�Qs��,��;ˏV3_,rؕ����$Ǡ�DEk��=�������v�m��h�=��3(�3GW6pɮ�w�\O�����ׯE�y*"ږj����)W�`�c6��K'L��@��C�ގ���}�y�\��Xd����+��(9_T��-���먬�`�\w�N
|�{�)�����}?�I,��Ԅ^������rR��wAȠh�ी���K������G�.��!���ian3eh���*�)���s7��H��^���1���{<��<4Kgͷ��7�S�!�ys
PX�n䁡oh��Ѳ� �)iff�έ[9�0�D�؍Xr�tȓŧ�G���Q�j�_�ˋ��Z��]nR�Z�~������иE!�$�mjD�B��p'�W4#C��N��#���|m��8��@ƒv*��n�����_Fv��?O�=���n�U��g3�ó��/�:�P�%Щ�K
P�1��4��Zo~�g`1B��ݡ�`EK2��F*�1W	��{�����51M-?�\����]�vȹ4E�)F&�w؍�t�5�O��=@�y���S.�T�����MIg���3��,�N����J��G��T�g��^U�{'P
�J�����7�b�^�\eS�m{�7�g��S`���%#nuJ��q��Q�C%�d����gZ�ԑ����8�x�4�o�F^���rW��
OQ�=�n���(�U��HE�۰�o(NA��R��;)���E袀���x,��%e��Q��y���vOr��pL��V�QY'��g�Ԅ��dL�Y��ST��	|h��n�t�s(� z�+"�n�G��A�� �V�f��r�W��=�V�/���?�=F^�d�"���QL���v��QƐ?�b�pw�q.!Qd���:On��zt>UK�Ƽ��;�+�����:G}&�`��d;G��+RW��>j��* 4�Lc����,)���c�׌�HW��#Vte-�j��~.�<�Zy��{��|�q3꽻�Ti�#�_�d`Ji��d��ҮY8������k�R�e�e�& �ܫ�;��i�u�L`+���ڥ�Eܵ�����~8'D�A	7O�C���1���o��I���RcsU�wn�/��Ϥ��PS���j��i%����~����̓�I&e�M`�Oq��
u%�������d���t^��H=k}����<˅�o:�bC�<r�*��8e �8��"Ɍ<�ߍt�]+̈́�����]:^(W�HW�j�R�P��wl��� ���A$7V!�h2TMe0�ڊ������kM�-���x���5$LO_&�%d�N<0�L+a��)_3M-�2)��"�}��A^���Hq��شr�dkj���l��\gz(���k�$��� �������4��_��ii�Ƹ��v���YX�����,�Ldu��h[�0�����>/�@�cT�[+(�2@�����B$tT����ɇ�8Պ�>9%H�Z�|u���k�e@ڏ�ТrM+1�a�!�ƥ�X�)�P�X���IlN���_�,�(Tɩjp����,aI�609�`� h)��J'}�t���җn�ʋ/� �úp�g���-�@�X��a�T,$���E1�v����M�z!ђD�UB}�������i{�������$�ʆ�/��ڨ�đr,�i++�ة���
�X~� �͓>-�x���o�6��Ot_�mҲOP�h�*�d�D����'��'�e����*�ā��0S�{X`�ɂ 4X�<����g"W��5��'~��1���XX����X�Ì6N���cE��}�)cS��٬�%n{�	x*j�l`N��1e«Ke�-�驪�B#����\�� ����aN��+��6~��`[�9�P��0!�C����X��>���^�@[E�b����3;G�~�ːJ+\�J땁��9}���������Y!C�%���j!2j��m��^�ׄ�+�L����X�GE;G4���h��O$��}�eWb�Kѻ��S������N��ќ�!�e���[�2���pj�~��"(�Qm���8#s#�h��7��}1=�.��X�������g�=25�(����$�Rr@YN<"݈����B1ڱ�#4�ձD�c$)M�m(���~r����_�v�B�����j$j��7�N�u��%�Kr�gz#��]�M �B+*�]��B��VQ�\ú�B��{Ը��+��qT���������ٱ�,b�f"�ܧw-5/u,m��m�������qc���T
�*���+Ra�&DT��3
)=���#lS��t2�f�Ӯ@�1:"�|���������O�Ku�'��$G�NL;��f����_[�I�
uD�h9,��XpN��6~�U�H]4M���ꕨ`�j�Xܧrqb�$j�:���h>�E����כ��`D;ϧ���0�l_���l�n�L$�E���'*���6cm���P�G����S
_b=l��ջњ\�L��`\x�Sn����"�������p,z���)��>ݭ^����V�,S�bO�'�]^�#�~����3FS��:nO��Ã,����k|K�'��|"��D��z�l�^l~Y�C�~��}�dV��XF�J�V=d �&�����$-q�!g��dBU�B�9R����;z*ɀ����8&���`�-i�Mw�����|���k^N�l{|p����5*�T�o��O��=DM˵]�۸�͇��nTd�cM�E*�d��
�zg]�**���*��;�l��o�^������z��*��u��t���:�(x����b�Up#[�K���^�y-�#�F���\x��HF��8|��Db����ːo�-��{��j����G8%��g�$݄Gr�B�4�vBz�2�#)��OY�S@�-S1��L����D�=��*�/����]�����;��FQ��%�Z=sWח�[CE�vQq��3va`H�x�9��n��p{Dm�I����Vܹ�h�A�|���g5e�ܼ*�4W>(�YC��F�@�6K�șr3���3�C%$�����:��9WN����J��SwF��Gr�+(eA�R�'^�1����,tT�{�㤪z�UюCR�b��z��[��<�Lw���K��:��K�#>���H`�0�d41z
VЖԹ2(%�^%�	�~�X�׺Q%�����@M��+�y���c	L���{dh�5SX#db�f�:2 �3���2�\>�>�ϵ�V���^|;�@���ͧ�\pht��
�����-
�|��H=��N'SSb̦Kb��J��A>���H�R(�.�};6dѤۜZ��O�}��+���N9��Yq�tT�oN�oY�A×��GӖ,�H��2�
1y� ձ�63�SQQ�ړ���6�1�tS^l�����2v>��f�/��o�g��蝽��~}zA�Y�Z�O�2w˶��[1G������%�G�#�|�s �ρ��������;�53L�B�<�&�U00�q-?��I�ʀ���D�e�fR(7���R�h��^G�Y�߆&�h� �}�x��

�)8���8�uHd �;I/j+Ў_>����/{�C4����O&=Uw�5�,���?��j�z��4K��?p�.�����dG=M��BIJS@s�`&f*Nq.K,����Yk��7�c��Lh�U�b�&���&u���O�)|3��8�bXm�5=��E�M�s]���TS��`�| I��jb�-����&[p��P^/�뷈�&<�j��>)��Y뒪�toxLn���y��s~}�g
��c��o��<X*xT�u.io�s$$o'��D!T�S`�Gd�ΌWާ;U��k��C#c��7�-+n�9K`��yUr�<��W�Ǝڥ�{s��_���*1�1�^���: ����n`�<��n�4(�>l"U���-�ҚtF�M\�b�8 �	�m5<�"�e�ϗ��k�M��l3G�������=g�����o@�p��:��{d�M��[yX�\�M,t�Pv[���;�t����J{�OS����Y�Η��,7�%�76Ȧ:�������퀦���,lp���^���**�hY��A��m�����	��	��5���6�k���1o��5J����*a��G�����]ᘯR��?��a*�EU��!��UC{ �$����1�P)�����q~��q�~�t8�yȀ�h��й�m��7�����;wm���7�t�5R��ݎ���?�Y�[�G�M��ʁe���e����Wi�t6X��D�)^̃\��q)o��*���2�&�������9Z�,��6� Zk<������N��MHpz|0T:S�&߭�U̜�.�q,gF5֤`?�i 6p�l��dF����)@�%I���RK�4\K�)"���L!H�Z`M�(�:"2/ip���=�!�b(�o`R�X�d>2j^� ��V���fZ\�����ǁ?����$꾰lt��%�����p� eXn(��Z׭� �2@U��W.���RI��j1�'@x��/˄0��u�BR�:�$�V�'V��,��J�RC&���[���rOz�L��.D�}�3G]���7�0�ת�����ۗ��\|wt�?�]ًA���6��X������D�E�y�4����^Ņ檇l�
���d%���f����h,�1��9�.VY��,{R
,�mBxҹlQ��eA�<�#�-A/Eeڰ&E��4�o�A�?�ɣ����h:����8mWxW��!���ӧ�$��D��WF��J�h%X�����f�#4�R,z&�8;��B�����cX�;�.�PB�\e'`�F��tŞ;�2 ����ő���{ݑ�.>:���h�Ewj��t��e^'�Нrl�6KJ{F���,AR��ͼZ�'[�>ύh��Ap(��F�Wg�|��^+^���XM�1���CQ����WŢ�m�U%���8���w��%Uf��@>�
0"�ΔY)�Fx7��<jW�����ʉ�=
�� gp��@h_��y����YI�g���Ùq�����j�_�I��IU�3 :n֜'���>kux�9x��.zsh`�X�G����h��q�ʘ<(,1GH�W�����x)NC>�E97q����(��
�r���F!E�Oi�l�#yC���E'(��9�;u����0x	y��>�;�q����3s�x#��T'-��'����S�Q}�O��Iޢ�Z�:h0�:�9���NZP.:Ɋ��}SЌ����X|�3��K�WA���1ip�(L$Z��t��@n��"�A}r��@'q4��;�s2)��e�x�,�ל�ex�o�اk��h�'�A�e(&�6oY� �Lr��(7�S\��G�VVȬ�{�"i-�^|Z��v�ʌ�����w��Ա�
�5��k=Aꪻ��$��G��y����lW[S#�EH] �S�N?��1��?b��eǰ#jpb�v`����¦�3�M�E)Rd/aY�և�4�R��/R��Q|�\铡`����%~B؈ד6�p��;���v�V���#���ߊ�}�И/q�� �4��9O�/�dV�� '썉��m` ��`������p D���a�7�-D4�$=�67Z%�Lo&A,�G|
$u#i9�Hw]]��f�p�)M	�`�p��[څ\6JI�)�,�+I�Ƶ��h��dȱn��;� i-(`t`0@�xwUXu�	0�V��b�`�d�?�=q��=�=��q�u�v��>����~�/�dĝj0~l�P���YO�/j�*���;�Q,�)
G���N5g�[�:�y	p�p�����G��K)��PSkv�����c�&᦭|`u��*�5K��pj�6|,�Xh�ָ� 2|�h>�ƾ����uC�M>yywj���g�#�ԧ� �n] �R��6���J �����f�ʤo�t^���W���6ƞ[tm9�+�!Q"u݉���5D 	�Ή��7_����M���4S�!��weuue��Xm�$����O��<[Ynyze�^=r��!�?�(4���30r�傿 w�6ˠ�5������ �Li���U���NNB�ڭN��9~o���&0y�À���f�L���B��t�*������.i$̢O?�UU=J�U"�� ��6��!d$���K#��5��X[��<��*�Y2��g�l����Ak	�<��V4Z�_G�� y�5�v�kyiiͩ.�|]�O��[�
ޥ�`S�M
ᦣ�3���n?�ڭ���E�-�6�u�!��䘀4����/��+��t�:#����4e�	����E4S[B���J�|���ʖkj��a�����p[h׌��"�9M�D#-�k
��5���n�r�B�+:{�9�)b&�V���m�i��U�
6b��m�D�|FCf��强���u��uu����f�{m�*���@�K ��V|.;��(z�o4=b��̯:�4�-���R�e�Z���S_��t�����3��럒�z�Jca3{ߋ���t�JB�|��eV��@K��v���i��B#���Vg��&�+��
z���!SD�T+W�XF-�_L|ڎ8fT���~�NOX!�y��a"y�Y!�"$���nY�����~�� ��-�X����q@�V��@����'(ܼzH��-�OQ�C��II%��ݢ86U�~��Q;a�˘�%I�;hJ7Ӗ���Ʊ7X[��O�
)����K�Fȡ�B@!��
� )3#$_~Ϗ��^�&�|�{5P�o�,JV�r1���u�o�i,	�jl��<�V�.��)�X���{��K��w�i��U�UNYU��uv�j�W�4�|�k%$�0�6'�f�;K��M:$ioKz��Կ2�e��,�l�e�T������4��"���Pެ��V����ร���``�|-��}{t���`vS�eS"^�1!P�Y���ܻ�&�%���A�.�`�%�-ia&}+T��D�]��� 0k��v�pGL� ���{��RKO�Qh�=&C,~Ū��U�\����44CY̭iy)r�oL��Rh��#_鈷�*~?��H��ƈ��o�Y����KtR�4�P���mdR��E�S�C�k����ahlW�;��t�A�vs���Ba�A#�����y���*fz�~����$�;6����?FV
��L�X�q�X�1G�S�j��5 �2��z.�ꌂO�1����<:���28��䰴2$��}=���U�D.�V���`h���-<|�l�l���W��'��Y�F����D��1xz��_�Fi!J��(f�'����20e��`F*K��З6� �x�&�0��B,)�4�L�j�С�ܗ�q_�p�[��$2'�]��费V��=�0Im��ԙ��=�:�FJw�!]�77/UzB?�<o��Q(�8��v{�������#7�ˣ��x��2�P��/��U��� .#4|��v�Nӎ,�c�k0�Pk'	�.���Ğ1&PN��z�~ ��8�8{�:8`���@Q�����ϟ= �O��"Us�Yp^�U���%M�,��Mj�Su�,9�3���YVd�Z���S�R�_ϩ]�܈�OLV���x@Qc!F!���[�No��L�7j��A봮Ŗ��
_+�e��0ܹ�j�$Y5M�y5��7'�.ڟNʹJ�W��ќ��a�`B�a(ং��j����w8�&;4>S�YC�������S��S���`dܪ��$�JR$��D�A����k��P����߄F�H��sڭY���i�i38�vZN��S��k�$�ц�:�7)�$9�+f�o�������Q"�uN��k@']�;^��x[�0#+/�X
z�ߖ=y�wL�����-�*+�m��v��� 1��Zb�$�ׂ�[�DK�u�Ԁ��R�a�.�r�vl>jQh�Ѽ���H�nWS�A�@��'����N�ϢJ�Q�g��9������]�d&l<N2H�+5��������������4��c�k�<7O��������f����t(��fG����1v�h���j�v.\Ie�!(���mu����/.L9���r�Cjw5����Ǌ~���ċ�jd):�o�XJ%�Y���!�c�S��@�2RP�C;JC�'j�.���2��V`;��Ӹ�2�R�"x��ݛfm���X�5�v�v��d�3^#�p��6���s쫽�󝔎a�xgJ���P�괴*:�ӃP������(�(����.|ۓB<��)>����/�]��M����d��=8��k��/�k��z�?IvӪ�H��&`
οl�)	��W��l��>|/�t����'��YBz�� j��'p�V�k��e�u�����
�M��� �����U������p�_ڡ�i4x���A�@�|nA�G'm�u�i+�|���[�����0�,�ε{� � tᏲ�7"���. ������}�z��6S�a��|�-�r ��X�p2�Xޮ�u�ўsO�G,�|�2�\��|�՜r��H�d���91�_��;(���<�4V���4�O�8a-���zˮ_�㺲�%J&+=k���� _�6 ,������� }5��!�ϻe�ӌ���Ep��.�h�P~�()�ŵ��-�.W���{>d��(yg,��'>�)E�(��'m��}q��Z������G_nw��y�UIT����S#�����Ɠ�[N��o��1d�&Ќ���mQc��N��lN����Qk�m@���zןVq����[s�������[�ߙ�_����9�!���[��!ε:�����L_�F�KM
{Q�	�{R;�aD�G���k�7b��"B�W�P���ڴ%���s�և ����'Qֆ��	��T ��y=��"��
1��օ�R��ir�t�\/�7G|���ej?���O/6%�
���7�3a�9�Iw�\A:���z��ux*�|Sb���(	Jh�%���ժ!zT��w���m�;B�?͘P��~��tX��JM��<D�,���:�B��b��ߠcyٳB�Q��_U�[�j���$`�E��&��ߚ�ew�f�.��,oT~�*D����F������d��D9��o�N����Ō݂�4��~�H�l劌&5�; ^��S�b��k�˪<��Q_��+��\�BZ�w[:��#��al	��ä��J���{KU��v#.�7�<����!Me��Q��Dᢂ�AD!���ƥ�y$%`�����q|��x`�\ĿDe���qS��Z���j�&�� �7������d�/�.���'k7}�0A�~�xlؔH<H
�T&V:����Oû������rq͂�Riӆ|@�K�rl�K��Kʙ���|�����]x��n�)=j�D̏�OB�P�gY�F�:���`�R�Ўf�W.D�&��+�믢����y���?�)�"e��oJ��o��9��|���y�WBx J�z��"B�}�K��XZ�p�#}0z���I�rp$"��a&R���[����f��r>��o�G�&�|v�oT� {c�����_�����*xhA�R=�$��J����N�`��4R���F�U0I��H�v]�҅Q�')��?'�T�müW��R7���kl%)C��wn{#��3L�Z$v�,"T��0(,K�0U�	���'�]����W�c��T׮�����$�_1
H���a���sĪC��S�J�f	�/�I4�Dք�8�*W��!���O��8��(��⮕{���w�'?�e��y�"x����:����-��cn\b9a�3d���G+q�`�l
��˲P$] Y"c�W�`xn��	 ����%?{i��c�֘CI!A�L湖U�C%����䮛�m�V��o����jr�I�C��l���'z�P�}V;�v����R2A�BƼ�����
��-Fd&	����!d�椡fG�[���$��v^��'r��?I0�����WmӰ��^�N�߶��l��m�y�g�?��o���gu�Zc��0J(�P��/����C o������K-�T���Ec-�r���U��Z��>;�L�Z9!�w��E�����E���m2�[�G`����������_w�7G@�D�0���������Ys�[� Sg�?�9�=��,�WQ�˃�Y�+'Y��d�v���m=d�c'��gX��-kf=eM֠���5��fs�a�����d@|ZY�l"e_������h�<@*ey�;Mu��Ӑ��-�e1R���������m�7S�Q�%R�G̽8�nJ(9G4� H�q4 i�o;�l:(�8�>$}���|$����Q��m���`۠�E��V��ۄޘ}<�ۄI%����1e
����.2���쒻��\FV��L��+��j��3�P���㍐i�s$t	Y�-D�ut+�ű��`#� �Оxp����ط�yV�M�p�P'/9������4�1l����U�8������2��M��E-D�&���t��A��v/AKE0�1�n�9$�/�����X�׏�MF��,<@觚�SٽXM��򫻪�7�v��:Aj^%�(��1��׃�k.�L����'�l0��������V���
���,-����ϚB�5�����H���v�9��'�QmD�o;R�%C���'��t��(��C�A<�'<p�r��q��)*�Io������XGf!���sS��.$�lS�
|i�,���k�0`�S.��Z�Ƚ^��=ځ��uq{�����g�$Eش����NBe�9L�� ��ret���itJ	D�Ѵ�d�IN�2��ߑT4Ւt��[Far�nOD��,���Vh3�����%|��|��{�"[VM:�c���8�Rpq�ջn��W�$�Ľ��@#ǧ.�0��4D^���5��C<B�n�i���f����-�g0i)��1ޫ�.����L�X�U���G�:	!��H�`i�������(;]6B�Ud]�z@Ln����t�_�7E���z��H�����k�݁�+�0����d�6���>R��)
��6Z��=>U��ݭ�&TTʹY�f������ic�_O(�P�!�M�6)7��f���?���R�5�z`2����#�I�\� �eW�5���
��K�U�)J�)a8�	��z�?�5�q������~5٤��<�:gE<��,�������c��~ �ʋ��V=�+�7x}��1h̼+21%*��QIU�8r�5Pu��6���e�A�5��Cݔ�_ԸT;YdN����ƃ���Y4�Ѐ�{��Y=��3v��J"7��|�	��Zށ����M)�<z��}��mg#�Ò�U
P*�k�(��K��O�Jh�69��5�zs=D\͡l�(���� ����~�#Q��_���b�rE �H��Ɇ����xO��7-J>�{Yͧ�kX�r+D�;m��S�@�\(�0U$��;G�U{�\oY�,$QݧÜ��Y�g�b�ҊE��YU����"���\��
2�zĽ���	U8m����|}�yX4��Q��T:7�J𝡦M�z]�}�M,������唨DB������AnE�8�NY:�ّO����D��F�,�{,v��r�e�",I�:��,�J&{��.tz���%���ߪ�
x�\�m��O��I�lL���3�~�Ϩk�g�Ge���ʚ���+~�bba�eV��ſ%�~�s���h��iV�j�Fk�B��kFx�¶��8���FTY�A"i����v���̬�5�T2��YK���P>	9���.qB�~Ѣ�K���SS)C��9@Oq��U�1�Q�^��	Ԉ���Xw�g�S���}r��Z��c�4������+"���sG&rP��������I�iu�盻�=g�W�k���0S�@LC�!P��\Bń�Z�Q�O��ߥ�܏�Rx�ow^1@��� -e6Xѽ �4c�Z7�r�G(j��|�</��*�s6qܶ��2��޼��J�[�����
���Q��w���v��"��[�|�$�󟣂�>9�|��x������:�� ;��Ʃ�f3���eEu8�0/O}�)
�s����$E;�R�$S2!�:�N_���D�q��=лRB��x���ab����F��>��p��r�q�:�㙢�L�Ԋ��o�ĭ��o�m��V�%���Aa�QC��:�j���Rf�s��y�n��r���̽V]�ӈ'�����ͦ��X�b�~1�<��&�,���A�P���n�<�1�o9䬌�����2��WX)���^\�"���E�tш��ɬV��"P���rkAn�k�������z���o���
k;.}.��������@����
�C�FU`D��=�Jn�l�ս\wY�׏�ϊ�LY�/w�ܡ\�A�&t̽\�ǽ�,���t����l��|�ز�Morڎ8�jc�&6Y�� pm�ʳB��i#0<FEr�z��H]�a����7E���qd����{v��s4W��*ZΞ70&���NF�9�{�il5�x��������?��.�	�����)��g���o$v[CA���x��������h!fp�^�?�G���q�AUy�NKV�`��aI~>�?�3A^	�e�s�������h/���z}�0���Ak��_�F���[4�w�����~�����<oZ�X���Lf6��~� .��p"�_��vs\�W�b<��ޕ�{]��Y�jF�����P*&V���J,ϠDӒ1E��������"2���(H��0��SR�`5�A�w�e��Ǳl|�����bRM��Y +�Վ�8�Fsr��N�p�*N�?بH����^�����(�|�=�D<�"�������T�~�9Fu\Y<������P*����D����P{k�:�d�L��#�'Գ�tZ"��4�]�mxX�>��&��EaJXC���4h[�Y�������B�a1��$��C@��)�wn� -L���D\��|����Q�uy�⹠=��Ժ����4_-��c�ɧ]�Fw(��RBC5�BAϔ��~��|���s�K2��c*�D#�7<����#5��f��e.�B�!ǉ�P]x	vR����A��tHRՄ��Y��%���G͞���?�^ 3Py��p4xD����bN�pZ���X�_f_��̟�������:|������V���tL:��a��\�ݞR���'�-�Ө'�у�]LE'�Y���Wanъr	 +���Bu����J��2s������2��ϗ�4讃�O,B�y���R�=&�"fIW�Z���)�ȴJI��I4��i��N��.ݭFo/�����u�|7Ӑ���F�w=̤t��U]���;݅��n�k���BPbv��<�]�}ޜ|:������/�ڨ��M5K���sX4��^h/d���+��5Ն,N/�A�-��
1H.����,�c�Ԉ.����]�d`O�'&�E�?RZ6��wX�䴇��'>�'�����;����e��(#qEI�i��5WVw=P�=�+ϛ�*�I��^*���ψ��hL!%�0C���ʭ�כ�aTM&�����a�����cWxۼ��ge�̾��I嘳T)��ޤ 4g�i�]�ewCR��控�r}M��s5i4��k�2��ڭ�	5)��"�x��E���u2#�Tgqɐ_iH�Y��PiT�jM��~�����/��%��ͫk=��� �Z�k�ʹ
ʈ$�s��l�d7����#�:+8�r���m@d�K�X��C@��˰)�f9�&Q��Ƙ8<Ye	)���&��n�n�RŁ��rg��T|*�-h?�t����brʟ��^����}B�m�ޒ~�0�����2,`����s*��͠�@tذ�A"����I�swq�i�Q����{R�� `fl#����-�'�v�.�����z��.%�]¢�r!z����Q�V"_�5S������F �4,2�7Ej��k 'Bx6��D��f�t��k�x	"Vm��=Ls�2*XÓd�q|-� �z�"��t��V0��݄�-�����;.�W��g��U0r8����1[ĹK�<��.�h�NZ��6V����D'��_����N���-��	���1�JB�u�{��b'��NG���[*�6����	"?�� ܩ�c��<�
��
P�!S�J�g
c�aBY�2�ZmRF�I�;]/��@���<�Z��@6\�_?<����jC����Õ�ܸF�R^Q#�ٟ��J��!�(��I�7U�����[���ձ�|���ԷA|��_��.��â�n�	=�k�0D���սk�5@�l�4���r�2ʢ�e q��M��TVL{)>7�ͷ��R���?��^���ڍe�*:��e��y�]��A��z�W}��p�����&��]��ƌL+�\�p�SC�|l�a�f�T4xLF���eڼk8IZ�_����ڳ�Qo�l�[�\��Y\��:��k/#������;�	H`e��w�_T�yW+��?�gR�Ƽ7��͕�k)t?W��~npm%Ģh�đ���a�8��#��f)��V:w,��q�y>ل[�]a��`�p(��o���$�J*����ȹ7��g�)�q��|��p��X�E�𜸥�_zݡL�?-!�\���2����vt�ۥ���9V�q���g:r�:4b�ĭ�[��o��m�>�XW��X�D%iN���8WC���O��W��0-͛Γ�	.� j㴽��|�f�Ԑ)l1J��@Y8���!t�����v;�f�eH�XS�8~�0�	y��$���{�A�&��x�ZZ��^�¹ѹ���ݒjD+�aM�	z\�� X	6�#D�	"�=t�h��	*�TCHjm|��n"�h8be31x���8����9�qN�����11�J��A��P��آ`p0�%'R��)zl+�:dS0��3�1��Ru9LH�d��Oq�:<c*_�q�2w����u؛��Lx]q�9UhE�1�/W^.�<="���k.g�I߫�U;_��y��H�-ӟ�� �y���+g�z��fX<�:�o;u�.��ó�C�)�^ӻ&�"�|��	��9�J�F"��fKm b���q5��I���]�R�[i�;eO�$xU�s�6�H�X�٧�\5�y�_�h׎,Ѳ�m�e�O�cy?�N
Li?�-��ԢGe��r���x���y|E�F���$�����
�+6��(�[��_G�%�7n\��K��ק�&�����iɤw�@rjA�:�;��$av��i7�{�:ܪ=��sL�|���mS2���5�<)�����s2�%�g�+$���hp�9��[���p?����u�M�q�x.�i���[��۔V�~�B۹q���a�}2U�ș=dB�INit[���Z�e��>���H?L�	.��hu@���trU��HrJ�+���4�Y*����Y B�B�(+��	ymQ�d��|����w���f�q#K��_�;K>1���S����<���Z���{`�,M#2K'�}��,9+���฿pk�&��c�G�}4���|?�HmېlŃU7���`��wu�&��K�4�x�8���̄�2ST�,�y٣Ʊ,�ER��@�~��y0��F��#X@X���1nѼLhû�IR�c}PPI��mگ&����s�C_���^��Tl`�l��x������{w������'<��kTҙz(e��]>�V㦍���q]M9��/�E�v���;�$�E�W�0k��F�X�� ���qS�[��0�)���RѼ�B�8�����*�*��%ͻ�uo)jvtn6�Zư� �~����T�G�t�4��}������İ�h�4�g`�jϠ���q�94n�*1�W���?�ذ[ۯ�~�0�a�.LQ�R}w��� s``�it����l۴�ꇫ�Ģ��~�#���{Gn�[B�0�Y���3�j%�|�cpW�S�A�r��j���S�¬�7�H��c=�C�Y�F�����+�֤riI���e���uE�n�|�h�E@����PB��Z���L�l�Ė�P�����i# 9FD%���T����]�Hq��ZW�>��5�%P	t����@�k-�B#3(:y�}������N-Jg�@6ɹV�m8ʄ`�\_������@� ��D�rT�
�=m�hZOG�po"��yԈ����^��4/X�f�;q�Z:,���������8�V\�� �Ό�)�|��5grkg���L��M �mU�	e-o�!	zL��mTaA�H�ŏ��0/���t̺b�&���W���6p�����{�^��\��Cg��v�?���1=v�֤2�����z����3'�q$���'Y��Y�~���¨�DN��1)���>���wc� �yZ��jԒ���񸟢)�s�uՋ�����ВnBJ�ɡ�Q�{F�5F��.}S���0�_ A�~&E3�	>$��`BZU:�7�l[&=KB�9;���^�NM~|��Z�M�qҹjf�~LP���k��My"�ؓ�&�I]t��`�4�(��L1M)P=u�a��i6���l!�PtXT��9�jp�A����e�_�wgO�>
�h��c����i���$�B ������y��N����IɺU�_�ܮ��׊��{$E��t���v����<���+<e!�zq�y�4eo���yPǚ��x�:}������#��ܩ�є4�no�*+#����_Aی�H�&�F�w��MRy�Zn�@�㢔��<������� �M�$0���k݇}|0y[�d���Tն� ,0��"�5܆I6�	�,M�Zɴ�,���S�/REz���̸{k�y���x�J�g )E�7�T�Fܻ�14�oZ��X/V�rٯ�y3)�4|aoRMYY��=_
�<��i�>��GQF0���J����Uo�i(�ƌ�7�X���
�-�e.zCi8G5i;���[ĸڈ�G�Ӿ!.\�`)���hH��؋A�OCdn�6�x��|���f_����g���#��-<�-
�܂���,��V1���}�<)������!���B��`��YM\�6�� �0>.�&��U�S��=A�������(����{JF��7�x��f�G�"}t�Թ�X��f�CvX�DT��q��-�aBD!��>"
��4�@Ԓ��x����@���
�[ʫ�.�M�n��x�\N9��n�q-ݕ?������Mfd��T���駓�ld�b�"�(g0�N4�u�o�[̇�M��f�)�6��(^Z���!j[��킗Nޅ��8T� ?'�Oe�2�{�n�Q�����>PG��v�vxz$�Ј�NM���"0�Nu+5k�X��߽�76 -��봲���I���W���/d �Lr�@������i(H���Y �2Q-07�®r�"�V�d�i᭲�in�� 2*/5��ֈW��Χ�y�����9���uqo��xo���ҮD�H�D������KL$̵ߏز�����L�M?63ƅ����\N�s����=�QG�\�;+!�%���Կ-,4a���-�,�\4�x3u�s����	ͱ�T\�����50!�+��aU&l��hG�w����m��B�B:ۻqZ%(��c8okL�L�bf1Ѧ���3��U����|�g6�� �KA�A�U�F�|W���=em��q���ms�ۯ���������l���U�� u�#������<��n�B\}Zn�6���!{:~Y;kk�Va��/"Qn�Ⱥ���*��!r-\��'-��g	d1iw:-d���@<ϖ���|��Z�f���}j��T�Nx���z��/��8�
b��-�PڤiƇ�X���<�ݬb���)�2����4$rS�D��w��8��j	�]ӕj�"b�Uʔ��}���Nd��h��b�Ľ'x՜|���=��xz��ݬI˻ZI~6U�c�<��������{�EQ�����>�І�O9n���9��c�0p��2ߌ��
�;��O����5����|���ɢz'��H���w���(,�V>\z�e���N��l��[戳}d,�h� E)�ʩ�) �N&�N7ݬ�����4b�*x(�V������h,����W��=Y����F]G�z�oy��k�S|�ި�!�u!g�G�+	��6�
����D���I�^G�����������H���Rԃ��b�#jDL�D`�!&+B���Y9�D���w�����sf�����Q�Z�viL$�"���[ٖ��<�D���>䁗-r�lW�mي��M�D�2l���(F�G�]����[e��������a�n�J`���y ��Nd�ެJjcw�>�ɋ�u.������[�����[ë�/w��]�7ރ=���w}��<����M`vc��'Ss��%!XG�i�d��^���#�p��貿�i,���KTBFH.>R@���h������2rA6�����в�0�џ��{t�Z�k3�~/_\\��������I������?�WG,2.�Q�M�O*�I%#0z'׼M<{�z�� c|��e�M����Z8I�Y*�I��3��[[���l�ce��c~�)48�iw���>�t$�hsmz;{��� b��j]wC��-�\�{�WW�.�*�ѳQ��+:�E@��M��N�e��d���$)�2�_.uZ�P�Eűk��T�<��SΉ\��cqt��rP����!��<��6�'�\�ܯ0>���l{J����u��5�0ί~,���Z�>W�D�����=��a>��;Y�4}\���82�3��$zL5��Q4��Gb_Ԉ&�o�w�� �ݍQR��Q�}Yç����$zj�h��m]�7/~���������2��~}��=�[�F5�s�
�C#X	/�3�%P)��a��z���/�7�ߌ�$I��j����3�յ� B:@ccĹ��)����۵�7�����'����)Q	�2X��ZL�6��f[���s����i"�;�J�We�qv��쟆WT�8��]�\Q\��"�	�4	�~�p��7�Y~M��/�#^���q#G�V�-V.�vY$��P���ܼ%N�n�n#߻�d*��j�����q$B�ϳ����� *G�(-�e���Q�wh� 4xAd�?�о쵑Xщ�����q#����Ɖ�
��6�.m�o��<�=�-�aO�\�a���?-x�pH鷺5�Ͳ���S�Tn��n�M��#�XԠ�f�K�AO���ލ@�/�P�����@Х4���̰��|R�f�>꫐���Aj�ά*�4���]�9�C?��	N��f0�3���r"a��1-���a��L,��V&t�@9�j�2BE9��Pm	g���v�<J���~0�n�#�F�IS�c\�H��g�p.�FD4����eON�%�3t� ��'G��BGk�C<�U"+រ^�:�	Ϲ��k�ZLXn?Jq��+���-d��Ѹ��6'H�bW6��bWs(��s��<��)"�G�m�<>y����(���`��������x�o���ٲT�TG�F�ye��z��h�)&L\����e��ؙ1I��nu�F`��l+�z�b���{̸�WU�:��m���"1��F�ӟ��Z��a��"%��D�ah#�+��i�r�?�:p�P*�Mm7��1�����Z���Nݵ(�ɴf�|��O��4�������o�w�ռV��+�*
�q��P�E0���ׅ�
�K�� �����5V���k��!_+��Y$y&$��>U��F�[��1��^��A����W����Ȁ/�ت_{�k��yg��9�ZV�T�/1����lpK�}������;����������Ll��*sɏMCZ�7�9��"��0��e����&4CS�|SF��m ��,�&�������L������f���H�ӂ ۄ�v������~D{q�l2�E�;�a�L��d�EF�!�I��\T1px��h=)>��Dg�qp�(1�y�����Thm��� 2��3A� �A]��:�.��5Bb���������FZr�N��<��?�.ҨR��`�����K���fV�U��]�s���b����j�#k�qA�Sf%A>{Q��@t���F�'@"����n*�H���î['iVE9=*��ٶ,ĵ+����_����y��n��ǧ�ɾg�̗��KH��vD�3U��(�KA`G�tGpvoɱ��.�)�vX��6&$���1.�gT�r�G����3)-��{�*�c2-���&�䊘1�_�>�$/��ns���J��n�<wr�՗�x6*S� ֝-�WvL��|����'t�=�,�"#<pe���m��ș_����j'j�[�z��j�i�=N���ܘ6�_[ F�� ��L�\^��]VO�̑���s�����يg��Y�t��0U�z�0��跌�a��ǵ�Zc_9S���<z~��j�1P��?��*,�.�.!��h��5����K��{pwwwww��q�߳�O�a��7k�1�F�z�0� =���'�Δm2�Wa�X�Ԙ��S���J?���aE?u�QG!~lcƘ�z��#�`E�U`TT�/)�$���/w/O9�����X�c�"6B5<"TA:�[݂'u�R������>����{�(W�0���j���y�.��AD��)0�L��;�`/�����Rp����������.�1�uQu��9�N�dF�.�|���g�w���v�y����6�$�C+�/�k�P޸2y�s�%H�Gq)��b7�����y,Fm,���wFhWk2B��E��Hq_Oo�D�>��5�ğJ��x��A�M_NC���Y�Z�mՔ�(���|�+7� F!�3�Q��BYe�����K�ǟ������C��cG��΢v�Z�x�2����AmDX��0D)�[ *���^��ʙ�, QK�1�г��[£�R��=�=�D#�I;����k'�$z	�5p�Gf������񭂮�F��p�!I*��hq��}�sQo��X��T�l��T��,:�9��y9J�c����~�xV�c��n��Wg��������i1o��s�����l�e��p=:��h-: �� ���[*�!�~��n �2N� )#=��fj&�]+���z�Ne�q�a�a��hy�%��L�Vzي�e�E�� Z�"���l���n7��z��![@Q�Rw�cy�0�۹�E��q<�g׎��{��s�0�A�����sws����)g[]Cڣ���A�X�p\���׷?���\i��ܦ��j�R��CV|����ԅ�(+0^N��� ��NZD+8���TV��@�F���<D�.��������s�#Z?U�Z/L�+�^�Ջ���QS8��"ǅ�5�f���B���>].��%����Ҩ1��H�#�_�¦�
0�ǎ��Pi�?���C�[��B{$���%��.�{"N�WF��/�����R�o�9lVj4"T)��V�C��׊N����$��T�V��F��r8PB�V�C���nbj��)�݂�"{���z���C�V��9���c�f��3R���+�ěKڞ3wN��]���]�����1��ƻ�y���,���+�EI�01m�ź%��>��/IX%a��~���r8Ś��o�;�q���G�x�Ű����]7rQ�9+�FBI���W�<Ȇw���Å�[�^wv���UR�3@u��[����S�p�lI����LER��'R2o���j�j�:�3�s��B���
��5�"�I��gEn�
������Ą+��|����F��dF8���${&�_k%����t-�2x��_e���������µ�}N/:A����\��0������(ƢT��-˗�BT��5�UÖ���>)��]��Us>;�^��#����1���u�d_�Ɫ$f:Q���-�o�ޝ�����+�n�C�Vm���#�,͡���3�?�E+��&��8���)����آ�i����{�
΍�����k��Mx4tX;�.�:��50����Ř��وW��:�>(�{pT��1�E����u�o��ר�����Bn�Z>�޴���d�N�yQ*X���ؠ������]�rU�Hw"����>Q) B�a�.7k d�:�:�a|���cQ�<���p�y��O���Xw��t�!$��:<���Aۑ��}����π������L�#z�1�F��C_dj7�����7iUda�-�U�|�vuс��;��9����x�ե�T�v�xk��� 8�&��	oF��t��?�w���TM%<��������?{d��g��X��/5��4�kE��O)Ѳ��=��(��֬#���nɩ�q\�ϙ��#����<.p>0~�_���mѤ�k6�SF2)��Φ�-
���(�ҁ���~~�F�ǤL���bI��<���m���װ�x�CMf��Rf���ͨ�~%A���j	�����
���,,΃�ݡF���S� ?���_(R�Z�k�����E����B~�E��4)0�W�\�Ws��z���Voe�[*��&�������vɢ��t�@45#�;"L��]lR{��/M�>��OT��F4o��41pY�13��b���^D~���Y��(K�v�;x�3W��7;x�.��J)ȇȈ�.ɼ0�塤$6����\l�"����%�+��l��c�X͉^��^���]�{"�
}�7Od��%����$�cTO��K����kVY�A���GF�F���#�H��;�H������NQf!��2��v�������f�D[�,�#�gr����3Q|n�:�ۚ��"���v����q������b{\g*��Q,-���KHn-��؝�T��7D��y�d��=ڥ����,."��`	����q��~@��IxP�0� D����m/�+[H����$���9m1����w�vF܌�T0#к��ڬ�)J��7:���3�s��������@u��H���yY���m�l �(3���/zJ�S�es�RT��MN���˴(E��X+��,o2Q&���&��J���^/���o�������Oa��W�Y~�������ޅ�&��W�w�'�����Y D6�����0�s�~^�4װ��� ���A�,l�S��-���S�s+��<�T78��&��s|�7!�#͙"'%�"�� 6����ú}�	�ƏXb�Z��#x��O]_��e^���f>F��:z�������%��kH=*
�2i�\�T5
fԇ*�\q|_S�����a�;:X��)���f�R�oeFў�.�}R��qŊ+`^�(��&�Ȥ�d��k�Jթ[�dh�W��(�v�Jќ�j7!���zU������
31t(w�]b�ڱG�L`�0�ù:����¨b4�8�|�J������v�v@5nA�	��� �#N0�H�t���U�bB�B��j���(Z�@�J1���`gH\P�}���ݣئ�u�ϔ����Qz��������E__ρ�C6;�������4-b�a5hfz��q��Ӫ���Q'�(�-3)��B`�M�K<��s�B_������Q@�8���}۷7�����&p��2"jӿ:����=��z"n��JaM�O$��E����cz1��~��������5���h 	�=��&����I�!�܍2������G�NM����M�;��q]�v���$�4�����R�x3�"Eh�����fv����..�J�B(�ʿigk<�>��cI�k�4��:�z�6�~��J�L�j��Y��Q����!o��T�[�C��ԑ<j��m�~G�Q��
+�F>��X8S��'����Tb�j8���S�<�����}>� �ժ�~�7������ڶu�޼�Z��g�LRpp��kS8��+z)(`��ZiU��j��R���&3����Y�`U���H^�7�'~R�k��2������B��k�7��#g4	������p��W�
 aX���S�\m�ǧ�wS6ē�. b��X�#����@&p"G~���@��"����?#��gGE�o���\����T��������w��~]�wqL�T�	�m�P�$�c�v�c��=Q��������ܴ���������#�8g��V<O��V����⢂j"C���ZV��#�ʴo�.uu�w�:WF�J��Hn����"[��`۸�T�k�>�r��+�m�+����e��U]��;��)�Ko}���� hf>�ʠ"���a��t�>�HR7N�`ž<@��dNj�g>�*1���쀯_��B)e0�8�C0�g�W��4��1R������U���h|����؛�=�M�}ٺ�6��H"@G�W"ߝSv8@%W������''�roҹ1�)Lf�j�jQ�:1xa�:�/��l �����B!�b�I`�mk��H<�-��@����/�F�qR��ˍ�)�Brb��?�Pdz���mG8���Y�	��Hch����7�B�C0+���_���ҏ;��{��b���Tʃr4{CNG�%7�>��'��͕�T�w�<]z>7bs�c�c�;®��Y��|�1%���1G����6F
�q5/��sr���?@ڱ|+�N�[�B�?B����"B��@�rE)̈́�O@�"�<����pދ�W�+���15�٬7U��E�\*�,��Z#"���h��`�y���%��6��ٴ��ݕ���K�)�3�zJ�y�_���z�di�fz��U�DZP���~�rI�Y��pr�P�ۖIFl�ȋ���J7̘�=ݭE��`�"%ؕ_��)���ޱ��4f|�gg����R;�I��7x�ƻb��q$g �V�pQ��C���d�Y��Py��럔��T�@�B��̯	�h���oXf�#Z �]2������o���XqȂm��=������o��Z행ݔQ�*\Ȥ*�w��:��Ҵ$}�F�qi_��
�-xb6��~�H���o��S�K����}E��\�puSR�:6�C���DiC	e1J�%� 00A�<jX<�+�A�oh�A�g'�Jx�h��=K>Q���9e&������:��;=��v��Eٞ<n�S�`�R����-7"�m�J�m�⩟Q����ǲ��7cL�Y�g	U�c}�ڋ���*��|J��S�bP9HB)WumB�@��ս�?yH��!�h�%���BK����4 ٽ%��CT�J����H�W�ĩ#�ڀ���������%Qw��+�e�!|K��-�ݘ�J�Y��`'w�S���(?#	i�@�j�uNS]�-3�^�[EeC7��`���M��d"���^Y�� �\س}CŊՑ4l��v����w�9@�}��fo����f�˛E��w3̙Î���6�G�M8�5JFIUF�DjsP�@_'68�/�K뉓��F"T�������R��ژr��=���(�Zz��;��+
�����K�G%���8�ި_J�-�+ţ�,����.G�W���}����lb�QWw�"��� <�?�1'�EG��� ��n�<��of�t�_���t޲T�ɪc�*	�C��oKn���a\�	h� �H�P<2Y��-�c���,��#Xd�ǯ0RS��v��=e�z����v�ޤP�M��}x�����5�(��#�W(O��� R��j �q������ܵ��4ߗ5��@���/��aK�2��C˵�ew#���\}�޾9S�m����]����������)@�@��KΣ�3G��EY��b�*��%wM}`��d�T�P�� �v��u��k?�$X���x4z����X��.�Qh� �aL���Tn���uy0	�����P���*�௶��wA�2�6�@��KKj�s�Ei��F�Zn'$��?P��u��Z��Qs�E
�D�*��]��Ε���gyb�SY<��D�O�/��Kv稽f����!3_�KC2�߮�j��xe�6���n�����r(�e/�ɳ���Wmsս	S���S�0fUmTʽ���*X�a�(��$�s���	 ����;+m�HÝXG�j[��w1,.V�h��듆��Ȕ��D~ζ$�{Hb?�]'�$ȳ��߲���Ɍ|a���~��.~�������zl)���QCZ�%]�Ԥ���l��,	���������>rUR���'�o�1��n�����T:^Q�}�����0	�FIQ��$��MXl{ ;�Q<�Z�#=E>d��Y���3L_��)W�@|=����VY�톓�l���k�0
dd�ya��G���+��������v�?9���ľ�%~�ס�nsZΑ�Hu���Mp�s��-Yթ�Ue ��ޅ왤��WAX8NQ.x/v�� �_{Y�_����!��[H�n�[�	n�D�"[J��< ��G�бu�W�'D	����n�H�pAv#�6z7s�hD����f��	�}�[��B�թ��`�����z��Q)�/��C����q��?.B2�67G�B�Y�ϰ���D�����
�.W+*>WSCH�|����E�7�s�SU����]7ݷ��~�LvS�7*4�H��թO<qa>�mD��j�5#�G<+@m.h!��O�YG�v,b�6=}�0ӭ���20,ζEk �f������)�^��˩��x��m��IN��k?=&yҺ$�˞̞b�\Nn�W�Ȁ�X���y��Z6k�
D-]�����9]������^[s���c��w���?zx@n���h얢�������~���3�>Z��{���IG�V ��<�8��0%���K�b`�|ېY�e(֔�w�p��{��p�BR��]Mnu�xSل��YZ� g\o��ڝ��a^8~T뀁G�J+Q�y��Q?1�C��W���g�K�03�%��J*��_���^�9"���� T��΄�*	%ac��rv��ȹ�ࣚz���"x��19<;��lf��"9Z��=�t�����+�൪�`�!�Y g�uB���C�U�ؐy*�p��Zs�;R1��@�55��I�ɰw�ՠb�34�7�a"Y�0�a"q�G��=!�T�i�X�]���q�ɾj��jν��z��|S��n�_|'�g��ؔqF��� ���m[�FG8��^��8�E4�h����젽�GS��-1�zG��Zc����RX�D�������j����^o�� �@��94�	ܧ�񸙙�//�O��|��e�!U6P y�'��z��5[��db����j��g�X�/�S�b� Q��&^�#�("�~��������)�ۍN�fl�ڀ0�י.i�Ľuġ��J��&�'�_���b�K��7G�k8&��j����MAh9u�
/��K��g+����^!D ���iY�g4������p�W7N_?(eҜ��(�'�8�g�_��/zcE��qjX'yzou4���p���;��e(r�Im����x�)��^��HW��|�	�TpN���,�2���h#����"���|�>��aܠ��>ME����OF�M�EN7�ȹF(���QةL�Y�3����L��<{f�h�E-pQ<�̣ܪ������ʾyy|X�=\p����6ٽW�li�삎�t�В��#��T�h���v*�<���w�Y	f�4��wl�>.5����@�X-��H�tJBN���d�ʦ�:w�za�'�Q�����>��?��&Bm����z��=1��L���)�|���Β�Bez�)h�����ʰ�'��V��'�C�w�,?�f�zT溹!�5�9)"��Ν6�x*���w9Դ��42g��_NIM
���VwxsZ��>q�x���n�uV�����PvH���{t�αy����k��VXu� ����0	G�%~T�
��Y��.�+*��Bv�ޅ�W�S�<�{w��Y0�Q�4<\`�Fs4EL����(�c�R���w�Ө�����4����?�O�T���D�E�4č2g5�s�;�K�4Om*�
�^^,|2�����6IdPϝ���gm\k��[.c�HmeU�B��q�Ƴ[h��_�����tZ�\����aU�œ!���E��Ö;`��|��g��}���v���tyjy��6j�T��q��ܾ�&�1��Wŧ��d�����������$c͛�-w:����S6��h^�{	��
2
*��/��ј�T�H/�Z��q[��Z#����[�n��Y^Qu��:�R��;g�Q����;"��S�Cq�#s�[�
�Zn���*�C�iH��F��? ����I����
�k�D�_�eh�o��ў
6v�Q��APS
a`��;;�p��>���xK/M�:F����߳�蜕���y�X��f��b���ֶJhx��w�S�\���C��9'f���ݡ���(=2���x����>$�1l������:�`�Y��вw�t�������S��?��S���u��S��k�/�i��:����霐�_�S>.�^��;n�`�T?�\W	��r =���R�elµ���:�7�φ/aqb�}qޕ_)���8�G�.���*h��T.��|Mmws��� �'�Zyׁ�p���W��m.��?�R8�}/�x�7���'��Y�K�r�?��VL��5������k6؟_�q\l/w{.�ĸ�o+t������L}�1=|U�Š��~ ��:1`k[R��r�ryi�ﬣ����^�!�� �7����6�Ld��_����R�x��>��;��o>U�\,�L���Qصה5�����w$C��n>��g�y*�js����i��3�4�b�㒗U@�=<�!M�B}������^��gK�w��ڤ~�0�4(̨�K� ���e�\JǤ��� .mqu,��Om"�x?e��?�4�uz /�k�dR#'7���s�*Դ�	�7#Sdķ�i��m�����:�?a���&?C�]+�/Cވ�v��`���t����=��ހ�ۦ˃[���7T�V7�6�ⵑG.1�}N�&!�6C� �K�{���)�S+�J#aQXi.�qœ�I����^j}"A;�&5�;Ր�D!�]h��i�*�2�v5F	&K�Fe��>:}���;RF��`�	eˀ�$��;FO��<n�D7m��#L��bwP�����Z'h����K�Y�&.9vƳ�^������4g˷�ar�+��ݧ�4�&ԧM��o��\�x��K�≈��S��~�2z����\\�B2-Q̏�E�> .�R_�f����J�a�h�k��6,kE0j�vt�w�Ue]��f�_&{�bӖf1�Wj���{����� �=#L�a~%��ˊH(�gKόM�����{ˑ�s�e��px�s4�ݑJ��Ҡ$�s
���4p��9W��|v��U,j�~�z���Y* ʾ�.���{1ǲ����.ǉ�i�,�|��[����8�G�rQ���2	'�&k�h�\�ٹh�Vm\r�<�|h	�Q����[��*Pҡq�w��(��h�v��b[����P��r���!\Ǚ�-�������|��}6���C8է097$E,/��:�oG�Z�mR��3�_nU_!�SQn���qa�*#��{p�"�}�qj	�M!�Y^JCѶ(�pr#}�lt��T�/�Y�u΅���<O�6��-���(ɬ�?Q@j���;q�i�µ�_��S�'XM�%^��Mo�Ѣ����?
R)LKDP�Q�W7��J��{����#�m�lV�\�Ψ(�bh�dsT'�X�9ͅ�k�Z�4���?������m黋s��m�����G*Vr��:��Л�����	�b���K�.�
t̂�<7��o�lm��4�=���	/�W�L�*?�Y5�W�@r}C}�d���\(]��ܰ����v=�k��Z�n/�/iX1?EA�iOL�G����o��08�i�?�W�����ȫ�`9�I��Q*�lh=���n(x\b&�J`��d���K�B�=�j��ӊ16��9�s��B�Feι�Tu|�iC�7�[9{�c�#�Եǧaپ���Qh��oir���l���cY����e����62�󷵡�P�b�zN�g�pgW�#�u��R��ߵQ^NҳbY�óy%�e�d̯���@~����#�� D(�Qc�4Lڭ���Q��4i�q7=3Q\��E&�:�΅��$f�����n�T%���W�X�� ��x�[P��j*��t/(�ֶq�Jua��cn!��m�p�5�|��������3��,��V��c��e@��C���@�4W�`$��D��پZ�l���Y���iR�o��=>�X�HS�錙S���=^t��M�^�U��j
d��tJ��8?�n<�0���=ؕW��h��XJV�ac]�&K����
����h�6��M�A�����C��b�̇`W:��j�A�[☐�ƙ4����3dջ9�2��a\}ntf���<���X�c����^(᝴�E�&�~4ꎜ��-AM�u$��z0��ؼO9��QW��#E�va�/�7y%;��M�P�rna�i�P�/ ~ljD�䐏8�}�"�̂ϱ�[�)#_�d�?�M�!Q9L����)�ˢ��ݯYi�Joe�=hrh�|&��7��(��x���2�V��]��md�ͦ�0zo^�!*c{��o�C�c��I_��)��-��h<ȿG�fIBڨ���!/���Ο00ј;U@/RȤ��TH>3�R��'{�z4��öj��)i�%L���R�W?�f��F����4�yE��QT���gf�X��j���Ī� �]��`ҾKK�w�.<�}�A6U�G_%O�f����8�=1��R����-d����]�[�G+��8b�x81k�6�eZ��d�Ŏ���x�\~h-/�l��ٚZT�}��2��t>N<��U�h����k�;,�!f�Ҁx1]_ԏ�'�Ge1�Y��-�p��sk\�k!��_}Y��\Q4� �\�݂9��&+�%��Y��x��~2��"�s���	��C�Z�������<�����Df���T�**�vr���F׾�l|67��aOÒ���f篕��M;ʡzwt����`��F�VX(�G" Dd8RL/�/%(��i��F�8ė�&�.���3I	<���`���Ĺv�;X���ks�>A�ߝ⹓d�S���[y�Z�'>�(���`��k�G/1��;�h�F�a؃�XbEhm�4��VA����Ȳ���m��.j�l��V��y!���w�q����$�M�.���9����w� �S�Q�-ox7�n���@�8�z�HFuM�d���S��:��Z���ߚ��A8?,�T���D�������Jk�N��j0۾�IZh�`k(W��K�Y�����޲����~Q=EIT�p#����i���V�@�j��͏¯��5aeEL�᝝X1>~m/j$��Rr_{EC�5z� ����%!xA=jn����qXCͿP��_䆭��i<���2��;Ѳsa��ָX��G��� U{�y98w�<�'9�\��q���r����`�\{o^���)��@���ؑ:�ם������Iv0  F�JV�2�X�=Lj3M���a������]�>�t�e����lwiT����@��$0�������`|Ze��o�hn#yr��4ȫ�_���gBE���I�D�s�(ۤ��}��se�5��Pf%j3�Z�X��~i����e��#g�x���s��if~{'�S����`H���9�H�w�1n�^�d��@Bo�|�0�֟t��Dzx)��������`�/��%��گ��*�w���>�>tɑ�
��yH�E�#;�|�֟ڙ�ϔP�03����{��Y�C�z]gn6�.���!�G�8��_�5�lV�W�l��b���o�����~��K�y�C���i=��G%�T��<�P�p,�J�JDl9��/FvJ��rX��&��p���L��hPG!e8ƍ0×^�j��鬖�����Ф��r�y�=�R��W$a�	���v�}���y�O��p;��(ۄo�7�L&�4P���v����`�������!�u�{�".�uu4�}�_Ţ���jn�/@첸�h���D6S+fv�I:%���E�q���`ձ^���m��|r�`Z�έ�4uU*{g��ܝ�pv 8<���m�JSB ��4��9"\��P���r]���:��['J՛Ж0D�{�����*$��&�+07�X	�a��aH+�;Ic1�J
J}�ھ6{�ޱ��o�$�	�i��R�i�Cib�s0�����e�~ϓĠ���w~�����J��5��Ny�n�X���ϱ��9&�YA�j̙d����S	�$��QC�YIk �y�$�tR����c�3���D ��G��Xި"(ԗm�~�W�����4}-�ƈ@#�J{��HQz��w>#��	P�`�1T8�ػi8��P���J�Y���� ��zo�T�lI9g�i�w���-r��˛�vH}��_���ܗ���|��N�6AFaA��;1it�]5Ϣ5��Υ�_Azv�IV6�����86B�����:&��}èB����wQR��st����:y8��H�Yw�����@L��R}1��|.o��\!7+��Ѓ�L��z|��,��F�6�n�ip>_��_[ύ-�ۙ1����g�� ��Y�Xk���/���Ը _�0j�s�~Ub_<Ɵ�� �S��~��b��f6�g:\�9��5y*MO/�qoU�|X���}�֖����6e2I�=�������|<Ƒ�W�ܮ�얩;����e�U�im4���V�s�2�v_r}(_Ϯw�K�4HL�6d_���3S�!~�p���:���!s9��>6H�w�N�a�pk��N��~�$�T|#�35�C��'13��5#D���;��㦷�vUU�V{ �wm�����-�HR;��?��\r��l��G8pn��>3��}ca�54�a�߁+�=�R�S@��g���\i�Sȟ������ͯ���C�BpI8i����h4���,��R��c�dk~5�|c[V藃I~��|�N����\Z�%&�;X&��=Wh�TX�g���@?���R���w$^�J}�l�(Q�g����#oj��?�\>?%�}j�+���Td���l�7$���_�UB��p%T���}Gb+x7.w�W >�f�}��miUF��)9F�L�i�j'w����HӮ/��gq�ʙ�	�gKTP��$V|R��S��p��1�e�
�TS�3�0$%�S�s��$\�7r�Av�Ԋu$�#���F6K(�t�S+>�C�& ��𲡈r�4�Z�XA;蒿�cw�]�I��e�2���C�x��7�ZK���+�u����]�	��h�<�0״��D�mvZ�U*�Y�Hmβ�-�'�gn�؍��	�!S'W��-� 5�z�t�ü���I֣�cֲ�fE�B�h��7����A��PYCF��1��} �#�͔��f�U\Z=64d\]���-�=����^�(R��Z�D����B�Ћ܁��14~��	pG7�T��֢���J�4��{ֵ��B��P:>�"/Ѩ�.[�lK!pS� ��O�ͩ2��;�ʚ�g�s�[K��n�ިG��V*�~׋�9�2�^�Z&���=yn&�(��0�nN�7l9��{�3do>��B�M@Z�O�e(h�P��c{��T������2ɽ�^O�V�4]�of���^�_B���7���Y�
�������f��Rc=@N$��0���k�Bi�@٬�i�W1Y~����Ӿ�ڛҥ���n��sR�Wya`/�*�ؗ�7�
�p-��ך�8�f$�9��d����W���K���霆.�I�9�c��fX���x��A�d0�ΏK����*Kd�I4��\�M�'*P��P��@6���XrbmjK��C*,'��݊/��t� �߀�ӡ1:3q��^����hW��׻9E1�21c���1Y�$���U<��*�!m�6��g�XE�������׏�������45��E�6V:�9Ӣ!j�{�V�"�xr{pZ+ͤJR�L���3��^��r���d/5N���!uzxQz�p��8Ϛ�p�C!{o>{�����[��b�[���K�۲EEț����X�GO<變����K5�5Zy�ݗs�V�;ڋ/�[��E��㊼�Q�_Z9�S%pkBe���*�$��_�*���_˪h��)|�:�U�dh����!�xe�hx����4]%�꺺�q�;/!����p�p&���32���s������-��^� 6���^�����[G2���s��;��/�/o��~TŖ2H�E=�(��<*�s$�ql�!2Oi���p���CL?Cx'���Է*��~?�¡�j��U �S<�(��I/�?��"�[����$~N����n�%�O�/�����9�C!KQ�Y��mħ��G�W�~���[4��d��c��
�US*��5�]��N�c�y�K��S��Å�}��YEsR1��ϰɰ5hB
2c���:���yAb�s'<�L�f�ʸ�hvܤ|�b��Gh���ú^����T+Lm��l,=.j�\v�i2��&F�� �E��N��?Mp��O��8��I��� �/�������2g�:ϊ#�y�l�X��t!3s�e"?�J�f��}�ą��W�4�'�نE$��6C�D������ը#��&T:���,-�ե�u����z��&�Ыa� �L��X�E$B����oʦ<gǲcjf;j���6:�C@g3��n��_��S萔�]\,����(F� ���֠�г�6���U�i~Y�ά���~��e{�������&��'�V��C�]�G�=Sl��tŝE��e�U��vV�	�nźP9���,����>�ܷB�����O���<:���@y����-��P�P��6��;�wA�Ƨ�w���:Wh$�+`�j��^��=��A���߾緫�_�F�� ���og��鈣���r���CB�ˁ�'�#�����%�1�����!�{\.�ˢ8&O�7(Gů��$�0O�y>
�ǂl[i���r���qqb�v_��=v¿룐ǧ��G� j�~���/
����Nz�r�\x�c1��L#�	i�H�#Rp�:��'R���K�ۣqwexrD�I]O��ӌ_�25���E��T)2���M����p��}�RH�y����3)�TA2��}<����z�9�tIf��	w��]�,�#�y�E"����������6�T�Y �(sS\S�Y�������|�k��ܪ��Uq�V(k�l���.V�3�����al��Cv=���]Gl���F��Eml1��O���x��,��<����p�D���zI�3z�h~��lĂ�'8Jt�����S^yx1�d��wߐ��V�6l�\�;�^$n��0o�-IP�H���Y�r������.�����w��e���[o1�
M=0>԰������@:�a�i0U���{nR>'�� �N}g8?<ez���9)	�]�h�x~ŋ�K�vś�ʂu��qoe��
R#螽
h6���s��ٱ�j]6�N~{���V�i͸��lj�g�����F^�\�}����0�&D�%A���ꟁ4�k�k��s�$�n�s��ϯ�+�N�;���-S�/���B�����p.`�gݬ37�xQ���%%�A'>����vd� 1F�dd|�Ț��$ܴ�Q)<þT��7�Tj<9�Dfg�Z�o��i0�f��uJ���� ��>"-�&�1�2� �Ve�fb���Y����<ȁ�r�|���06�<��ʟTm�:d�>�nd����Z�Y�!�'��*H�N5����'���XK>(E#���?bWaA���4�G�IG���_�W��?�l�W �����T��=��@�z���k'��n��f&MԞ��E�� �"����RNg��$��NI��=�%���\��]M��Kk�6�br��K{Wq���ӡ3���?�߃Ym&[�Y�K���e����иq<���8Ʀ�˂l',����UlN���/�?�%Ck�:`X���;�.a�4��Z�T uČCϿ�˶D:
4#I�y���[����S����ۣ�D��δ��
�R�5�ϙ�D}-_��%��� MER�#�%��Ɣ|UE��@�y�~(�Yn��{?��ߍO�%pY<����A>��k�L�Tk_�c�Q�!o���a�A�C�WKf�K�By�.P�aN�!g�En�A���?)X�7�-^?�w/� �!�zfg�)�����V��	��掴�T�:^x博�+�Y�&�:�~�z��d�歗]5u�[�'Ld�������}��ɪp�pA�R���B�����K )��"�I���d�g8�Tv�x��|*�^Z?�b��坺̃�|Y���z/	S�{g����H�zQ����υ����%�})8e]�$�g�.+"���oQ/𗹑E�`���֟���Wq�)��E�Qv	��]}��+St�9��&�C4�[��&��&U&���|��t�55�T���)�+���jk'��7������<������G��<�y�+?��J�ߦСY��f���q��3t�
�?��D�t������hK��M�cb�ny���m�|N<far+5�����|�����ݚ�R(�*��ϟi�.m������ש)����2+sZ��`OhD�b��	�H�ģO�� �F|4 ��[�>�k�f$�&�ԡ�c@��_Zī8ī�����b3�V��H�
h4H��.e�2�`��ՃQ_`q��:Ey��䥂;�_	I��B����ɝ*����^���ʋ�DE<���Җ�K-��d��y�&�l��ZS�0�'M������I�W�N�?}9�=X��I	Z�oK���1���˖�[�Ku��L�"�����pc2�N�)������������o7X��4|�4)�1X��y�wh��Ϥ0�,_��m�2�U織�L]�:C�ԃνc��i~��W���O~�m-�[CcF�p��1G��i2��&l��a�(_�g$È�p0:d���ߎLVʎ-d)��� �b\?�җ��ݛo�����phE%1�\�#z9�t)��t��4��=�4/Ѩ�I�����g]	,ц��Q#�[��o��j���T411�gvT�]���3*4��sN9VkT�J�<�K��e���n�CTVǪ�U�RI0�U7�JKѣ�z�2�X@��MO��ZZZ>�hR��ӳ��(��^]�^�����k{ð����ae���}Ŷ����街�	��r|hh(�]�!:o��0Q,��FG�����R�.���)�ͥQpQ7[,E��7֠����\��a^�4s�H\�=�Ōҋ:��!���"��|����u_�N�Y_I_ѩ>�2���9��X�p�*�%3Z���y��xf�_5L�B5=���˛MaRL"���mo$*�bW���\����I�(yΙ>4�ɆYZ5�۠J�	�)|B?A�O�,�	�4��'��4���&^7��K��#�4�*��E�i�N�=��epY�����_�SM)�/K+p�n���)�:�'���>Iv0�%s���fae�e��D!3�/�7��[~�����n9<��Y~Q��4_���p�G�S����/���4�-y�u���7@Z7�/��ru�����c% �� E�s�޽x��[�x�-�T��42iLF��e�ѢE�X�T��i}����J����Pʤt�����=P
�S6��r��a��<bR����B$�����k���+���-)V���i�j4@���h�Ǚi�8	��*lPq�����s�}#��.�ѫ5B��r�X+�GvyZ3Vtv�C�fGs��3��F���SP��"�?���+��M��6��I�&\�6��6L��ƱCaB{�5u��y����ua��ƸsC4��K�3>����,^-^�mX�Ӵ��������#a�y��/
���F��x�؈*�LyagWn��G&Ô�\cSX�Q��'�0.%qZ�s���)���J������|��;�*��7E;�hg�׺����\�Kh8��ؤU;��"��2�l�����{Fn�a�$�#������v?wg�^�՚*��8֞T����-.|�	�4}��G��$�8�4��?���x�n�����i�p{|ҩ���fBSZ^5ig���X~����ˎ�������5��+����mx�`q�0Y�V�\�� /D��C.�+Z����L�!���m��ٰ����Bo��l~�����_ ���y�}IQO^�{����_�m���ۃ�]W�� g0u���S:�J�AB����������R���t5151�xh�};G��%��4�䊕xMe+L�H�\�b�H�3V��$��/�n+H�^9"�JؽWbR�s0ŋ���k�o���=��.:fY�-�Ƹ�I�YS�N�M�ƽ�]��a����h�"�m�X}M�\�F��;մ�DC�Ь{u����Qelo�l�|>=�<����iR-���넥�Q��: �1���Ag��h�ᴎy?x�fo�Bw߼0��Ѣ����K�C��ë���{����X�5Ea����.�/��?~�;�]o�G�\���!��Y/OI���SQ��gse�ɥ�8Wq����x\�)�:U>�+5�'F'�����]=�wvu�j-v5�f�#����~�	����O��{	� �7���U�2?����5A�¬�U���)���\��h�=,����0�í���N����p�C��O�َ˘FB���G����9q-���a���i�nl=)���F�8%I��� #�SL&���)�I��4� ��	�caɻ�	�q[�� ���F�g��d� e$h�R�R����d/ڽ{�ݑI}�� o����-�'�f�%�w���q���q{=H�p��MF�-+��@��g�}v������Mp�nN_u���eS9�J@�����V������|�e�DS�.+����:y/h�(�,�S�j��`^�1B��g�AT�P�p���-�.�!~2Z�5�N������&��o���[n�e��xϗ��Y��񩧞bϕ��4������*EpPx�������h�p�:�U��UWl�
Z3Yv�/Ǭ3ˊ�2M��f�T�̖��#�x���Y��u��2V)������� ah�Q�o���ɸ4E%-M�-q��;
͍���uj)`�����%}�����T����ŋ�2-���wq�3u$<��S��c��P���x��ptb8ݷ7ߦc��[�0f��ɡ02�+���IKuDG�/���1���:=UZ���ѡ����[�Hޭ�}�d��`��M��J@u��bת}�P��\�U��9���r@��P.�V�9�E�A�6�>$�	�v);�嶴�0Oו�h����.&���*e(M��e������Y�=M������3K[��x>�N���n=i��/�epd�r%1��pn����
��I������<,��^���V��G�����,�L1ܺO3��*�rŠq(�4��g�������m��Te(�8�7��A���A�0Xg���,C<pk%E��/�h����K��\�].u�s��z|����bu�:�nf��,a�0����oS�4s�a�1ƒ0��xqa�RV���Y�B,p�0?Y�-�V琌��iovʠ��R��jT�1�Ƕo���N�c?3e��c���0h�z� ]z`����]9�������4k��H����r:6կ��qڵ h�&ttvX�ңoj#�(�|g:jn���*�����W*4L}�LnLK��#��=I�	]�ڧ���9���#Ѱ����X����F
Vo���^z��0��k��y�q���ц�a�f�^~�@������ǆò����u��jM����33Z�K��M��ƨ9r�ʊ�\S���j�i�A�^��F�F��OL��j_���xV��� �sX�{�	\��K�ڔ��K��߫�w�^P�G��Q[�]h��=���9ڥ��s�Nc��d�Ӷ��G0�.X�2�M�n�� F�izxȸ���t�|���a��/�����T�-�1�$�GY��/��o^`@x&.�w�3�m�̚�4�pC�L�#q�x��-�}1���Ţ�n�ɶ�wUj��V�0X-*K����yϦ��CKZFI�B�\�QK��#���K�wzm�� ����4�Ъ��wGm�J��g%PW���.1�F	�����m:�b�fz��)I(5F�Qo���>+�B��۔
c�p� �� YF�aFʦT�R1���`F<r�nEg�����3{JK�۶m�>��$߳��׀0�tEF��Vd�atC4`��.-�iuob���O��]����&A�c�;�	��l{<����cf�*ߜ��b�_>+��E�w����cK�	&��$u�:iچ�M�	 �K�	݃�{�t��fru�D���H[�C�f}s��0<2ƥ��[y^��ϖ�C/�~z[x��]��Nm^�8,]0ZۖD�o	�����āw����[.����Ѵ�����r-Q������������UЅ�ͅ�CYK5{U>x��m���U�677�j��q卙�婲�A/uS/��J@u�Q���S���z��m�?�����Z[���s�����0�\27q��K�L��_�X[�m�e`S�^�G���!N�p���OUR���xF�'�7$I��^xW�T@'*�<�$<M?I�a�����U����l�����e��itH���JCB�+[�2L��h#M癞�����o�#+�����e��2��cǎ�Q��R����צ�'���郞4������}.�������&N�����֐Y������5�\��T祙�=���\��d���D	h�_�}��w�?��?sI�Eb,��#�Q���LO3���i|f���s1�I�,�c��F�5�iB���1$u�� �x�A[����p�;�qAN3]E1���~��菞�iB�����Qt�pY��%��P�`�0hhu��!ì%(�G��`>e[�Z�f���h���z�)�*Ƿ�]Ԓ$U��@�c�����~�N��=���g�t���VQ�1t�ų:B�*��G|�6���� p	�f��-�5�i��o,�x��x�4�u��dk�iX�6tFŉr��Ph˷^:V�����p�]�����K��hy�`ؼ���=4n�����������.���C^g{�w b��j錦�)����V�_�v���Y+�v�#��FG���CG�G�����-]ѷ���� ԯ۔����!�^���jK@��٦�����I� ��Rc��������h��B��3|��k8�H��)��J 81n�K�'M�!M��N����	K�'\�i��q����|e��p�+����I�	.-�=��4�$��$�9-�*��}��Ie,�������Y��a�>�;|�ō��e}��k����%-,�~�ϛ\,8�L�Rm��'sJ�嗖# YC��X�$��Iܖ0�O���'��5�K���)��Y�u��%PW��.���g�`HbX������;߹���^Z�>1<[r��#fk$)�,��� [#%�B1���[�8Q�P�`���L!C�I�	�����\��F~��paj������ֽ�KI�@wN!��I[�E	���Tc�"�h�]���Hl,��"m�[7�Z	�~�G��7��޽{Yj�`b�T��B�b���ST��@	]6��p3��@@������]٩��r�ҭ���*V���e�x�e�e+&0�*|�:����Nh3�619��6������jjn
-y-i����ѓQӘ��
qI���J��ɇ֕���dQ�օĻ��FGv��Y���r^�j�`��Ү����{���hXt�a��uqS����C�o�D���5����.K�1�����Ьˆ�5�ܣ����wt��R�F�G�E+�͛wes�� ��^I/�\~��N�,N��� �?��%�z��U��ޡ�P�m����N{����hS���q%��m��~��l�)n:�;���!�W{�V���e��h��U�������U�X�Mgq:,�	�TQ�_
�x�:�Y�����T��{q���SH��c�y�IxZn�
%�a{�X�	��7��n_O�|Mi"�a�ǿ��S����'����C��Mn��	��_�R�����W]u��K��ܹӔ/����A���1Z�����ЛМ�-�%������?�ݐ��ɲ����E��.�짒;�vغ}��+W�/�z�g��(4�Ӫ�k~����s�=�]
R�gxȖ�VY{��ܨ��2�H�^l��(N��p����'������a<�a�0)�KOk#�ŰP�:i�[o���뮻�	)V�]�f���wgHyDY��%҇�&&�t��v"{��ɽ���S�?�Pi� w�F����~u\,���J :�Hʳ����C�h�.���[�7��!�P�p�)��E���S�W����i�w�13�J�hp����(�`MUE,pmQ�Ѫ�Лb��N�Nj����j�G���V-�y��Q��]\�z����{	���7*N����W��_^vE���]��?=v�D8~���[��m���s<x��5�g6���T>J62ܬC>�ڴ)�\��u�FG[k<�Q���j���54���WI�}D�i��zý*.�@��S�2�d?�P]���=n������6H}�6D���0���MđI�/2���2@�	,�Σ�JA�9`�g�v���T�U��+�i�ŏxIK_�T��8���T@��Y��[:��k,-�f�J��$L��$�t�����4���M��ݮ��<�X���=]��iɝ����V&�[ͻ]�;ӌG3H{�WP����u�]1J=�1̥�� k��3P��,�t��,���-O)�[:	�����ޛ좴�V���w�%'�u��\p�����x%���J�L�L��a�8�K@k�N�Y�#׷=��3�����tQ�4r�g�&#�*J�Á�1z���/�.F����	�"��
��!�?�{��P|n7�PF��.���"�]|��o���x?e*fWs�V1Bf��v葙�������J@����|�ћ5SڧY"��
(4�/�
!Cu3bf��I��c���m6I��;D��Qg���	I��N���p�e�������X�h�,���-�	��.����CS�E��(���:�*��頾�|��5�c�K:RP�����0q�1tꤿ��ޛ��:��]����G	���pE���X��]���������]o��c�o	��G:�0=vD�e��%�B[k[|��	F3��Sӹ���\C[}�a���O�<<������-^�>�RhQ.U8��9�w�v��Մz�gI	th������ҁ2�R�����@�:�B���lBB��<�La�ݴS2�7�-�3����?s����0�8������vl����OY �" �{ʊ0=s�F�Ù#�a���S��'�����l܂Ki��������ݜ5t9-�G`�,�	�U�'�|`p� /�%va�����_����S�t2�e������>�[4�+sqc�s�$��I~��U�TV?���2���~�ƍ��ZY� @ݜ��[�i���8�K@�n=��k����ݨK���YSs2�&�̚g�Z�I�R�i>0/�`�ō��~N�WF�0���Fh^i����O	�ċ�@Q�^�]��z@��M�xw�a|�?JkV�q�J����{�H_�!�=1ig��Y��Z�?�H�fN�b������WH��Dɡ���>�(M�XsR��.��:<��|�
�R�L�!>u0���
#�S��TE�T::M�w��Rυ�P��EqR9$�T�����]}Ԭ:V.MN�qhno�u�o(�ES�I,(�O��E��><1'{���3�X�!Z�P����W~�D8��ናk��x��q~�ݳ{W���ODW]���b��0�����@UG�NG�)�*���r,z:x�p��֞SkPyEaϛ��C��-ց5--lW�i��	�U��
V�:���z{T�;O3	��4�ơ?�4��ib��C��Kyͺy�8o=]�&��bgL6��5�zJ�C� ��<^b+L+(�G)͔�8����/���hu8�4�����|ZN�>~2�+�9�vRS��fq>���$�eg�J�RM~HW����lX�M���ls{8ieL��#�7��4;�����m'@����3[���T�d�㡇�C��{mF��Ix24$O�	F�����~�2���td����Kq뱼�ghuLN��o����M�����VD&��3Su�*Su�g���x�>M�_+�����!!\���#�qb�B�Lm���c��Hе��	s1
EIxb1?ch���X���C�iegLS8���h�Վ�*��q]$�O7�x�+���Z�b�����q�l�!A\:_a)�H0N�ps����Z^�,�{�>h��x<r�:�u��W5:ɍ�����h��b��(���Q�������G}C��&������}c�Y�trQ��˼S/�D=.�Uwl6�i�e�M[P<�%��Q���NI�)�R��\V����X8>9g��m��څ%�J���ǚ񚘘�F�ji��T4�9
�/��-�/\^�����ݯD�#aӲ�hͲ�йtY������0~�D�溛�u�\-�}��hdS��Mk�P�̰�,��Z�B��t4:9;��X���]��)�Tf?Tq<��@X��^�u�3WMj3[4��M-\*��v���* ��P9��&�W[0>J[;��}��Nc\�u���~|�v����faN�Ļ
�ӑ�W�G���nO�=e��rq��،����ૼ$
���ɤm��?�ʿG����_�f]����IÔvV�ʆg�U�O#'�$�T�q:2�t\�׉�T�_{��^����~�#�=�SuųL�σ��R?�l{�?��w��������X��{�ڥӌw]z��A⧅�r���Pu��=R��/��.	^(���{�^k3� EAR��J���0
�=s�:�>�u���S'��І����q�a���KɈ��Ze�W�?��9��)�LH`~�/��/��!/
�ć-M᝕ruH�ޓb��$0/�B���3Xۈ-Xg�
.G�-�3���g|:.}��:��^q���J:Q}3S�Pb@I=E)@���L��v(H�)��LR։�B��K�d��`�Sz�����R်K<����R�1��SV�b� jX�Rq*
SEM��Ҭf���j�͡EI������'J"&G�bY{��V���:�o���0Ow˵-\�涻��'�'��k׆�˖��6���_����Ç�c��
+��:�/[Zs����%�-ZR���4hҩc޵>P�\�	KVR�v���c�tqV��r��a���W�Py�,+�s�G�;��Я%O7��o���OSb֊;	M V��ke�m���%dmoWs�$��N���?�z7�`�3Q<���]Z��i��MG�~�ڑ�o�G�G�#;�w:�Q�[��x�/�W��Q�G<��x�؞��Y�(����tR������8�6�	��P���IФ��a��$~�-?�=F�F��c�/��d����d��V0�����2R:i�zX-z7h�,y�I�m,Y\����b^���k_�j���=�����.��r��˨q���D$�����o߮,�	�=bƔ����+f�{$���V.L�h`^�X9#S��a6�0����!��I��ū
c		�
�F|8�� ���_��_�PL�9)Vٔ���:	�		ڗ��ȗ���E��a�N�H/ϥB�_���K@�ߠo�QK�)e��V�.��4F��c��6ӢJ���zˣ�i����F��')��dI�.&
���D L2G�(���[�ke6W
�)v�'m` �A�7�孱I�h�j�VS!45�D)-e԰B�Ռ��=��J����T��fJ:�"j	͚]�UU�0���6d���ə0\��1Q׼��{�U�Bwx��+<u�=���b��._�8lY�0��O=��豓G�k�#��84�%%jlB�5C���t�"B۬��Ҍ�����f�ݥ�LN�1�9�^��LO�����j���;��8��]�E�us�3�H��E��Kj�k5�i��*�d x��
֪U�25%��x�"�&�U�\	_*�:������K��3~��lX� �E|�k���*:�xC�q�Â��r���
o��<
��Hz����(	��[�f�A��{Ix������+M�wү�K��?&i[<�&c���xx�Nq{�zɛL
U|H5�N�C��~Mmk֬	Z�b�i�~�hϞ=�GN~��u����|%��o�g�~"�/����
��A4�?���k��f�f���� �eĈ�����+W���� gs	�9�$Ϳ��;����b5��ik�a�N����h���i�Fb��`n0Af�� �҉"�«.�3&���6r$���4����|��lQ��a�긟�]V;�o�~��?$�T��>��ܨ�nM��6�V�a��tp�c�b����-Av�I*gf��5[x�6�_�e��}�?gJ
WAu��f��{(�
3E�w�a����P��YFB'�:ju�gQf�%u8�5u�S�E���f�)���l�
�������WI����ʚ����Ma���렊)��765kX!*M�jFN��k��VU�i�S��j|gg[��moE)�q9�<>����eK��ؤK�w���5>w,L�ra-�	h�wo[G�Ů���n�-�^��n�)\p�f��ya|L3y�&��?9S�b�#6����!�R�F7�Î�e�W^�J��RYl�7a��)���NV�z�hH�KT׷ky.m�G틥�/nnڐ�`�UK�hSg0�sS!�4�)uMi�J��D���D?���K�9��z�nJ����8�#�����5���7ɇGK����O%�OU<��6�NK���<c�+~�w�	Ui���ɦY��⟁�xԙJ�y�w���S���w�O�oWKV����d��n�-��#�=�s���������>��<�&[������}�d�)b�y��?*��y������]W�~���9�W�[/���г]�/��_��}{�YՔo)��E�|yI�R�$X-^�̄�R�����������h=����`K�2Ƈ҂��I"�"l"t�,�p����``ú��!-�K�r��>�Qq�+k����͛�u"�ͬ�6Bt�xGe��˟Q��H�}�V}d�^&ͺ3)Չ�F����mR�7H��td83�y�&�Z�����g��`�*���gʱf��H�14I_f���ةc�W�3�����[��@���)_-����;�CaS���[):x��=�B�Bq�0��
8��7!���=�̇I�3�8MJ��Gu�TN{�P�f�F&��T=Ϯ%�¹��+4�LE�Zҧm�a�ء(?���u���������sqO���a=��Ļ�y9�p�.mi�}�í=�C��ᡟ�4�b��(��W]f��kdr:�I�!�%�J%�Lc-E	q�L��i�l�.B-�E���u�p���C����o��.�����?��ReQ�l��m��'���퉓'o:v����cvo��/��՚�q��E��Sې��
~RCä�fa��
�)`�CX8e-G�gps��ҫ�p�� �a͑!�
�^*JmY@��w�X���cno�����i:�]k��p�CNg��p�#-�8N��H?��J�����ɦ. �י��%��W�B\��e�������|>����<'|���<#9#Ҍ*{����;/��?�c[M��c�kJܬ�E	Ϸ��	��B��E����[)��B�x�b�-�R5|��׿�倿�!CR�y_%PW��WqՁϖ�1���g�������x��=}(8tz�N6�������K�����;o�c��!(J!�M�0*O�V�S�0!���00�>~�A�3��;�M���W^y対�o��ꫯ�b���8�����Xwy�`�Ќ�f,~d�6���$`sj�#U�H�n�#k��2OJ�6��_��TgXz�ON�U75��3S�"���|7�����)�t����O=S쩇��
�?��Im�2[n���4�p�
���>-�fЂ!=)`VwH�41�ZS�r�V);�x��IkɒT�`��L�P-ϳ6���n4�`��x��fyK�s���j��A�gx\��I(h՝U���+�����h���kO?fv�.R�K/</ܴq}�����E[%����KBw{G(�j<�aJwni/��v��txg���
q����D�eIn��N��W5���!�Nq��U~T���y��\��T������|nhhx���xe)��I}k��(��CE�QM:��������a*��شhq�,	�S�Ԯ�6GLlگ����e�:7jB��S��]Q�Y�I���3���x}`gU�	K?��� ����iʆ��(�Z㰵�����&<���;�s�������KܖO3��eb ��� ʹlՎg����`�[��d����} ����Z�ni)�)t�c}�p�Ϫ,�*�~����� ��?I����x�N��#�_��\���ß% ��m߾�k�����v�aN#�Y�a6Z�Q^��_��rP�كp�����Gp�Pk��F�7��A��b%��:E����51@[R�p&�e�ğ`�G��7۷o���ի_U;��(4���Qƙ�1h*F6�[;��j)�b�N$.��+W�Go���"��몧��nHG)��*�����kYJIňo�pU[;��:@:P��zG�ۄ�:�
p|s���O���z�b��Qޮ��i��Uku��Zfʚ��Q����J��6�R�ˀJ"iC�W�]d֌��kj��kvIC��H7`h{K<���ӒB�LI��X�"�t��0�|ex����o���k���Z���5�Ѷ5kü8?��/�G��o�6]�-,^>&sQR�Rۥp54[�.��q���Cr����ڧŬ���L��ĸHo���\��%�ͷ�T^S�ۇՖ��O�;v�=~��={���Soi�)�+�[�J�Mr�~Y���n���\Pw�6bB.i&4Xn=F�l��~��p�v�*�L\�--�	�c~���ś�gi6������׺=o����r�xU�s�z���'�bn���~��������Z���?���~�z5\Y?��~�Ϸ�1@�&�)^w��@�5�O\{����g�:��c�3�sY�g}<�� �cD��e��P�	F�����꓆�l�2�����-[�0u��J��\}�r����J F�i�^xe�w���|c���6���1+F����F^$(6����լ�	¥�z��T$�F>�;)B.�`��m�
o¨�6�?ű���E�'����ͨ?��W��}���1�
�X]'T��d�Ӂ��P^z�O����_�Y�Q�������)�g5Z�s���-��ZǭK�:Q�DtN�*�T�{Qu-��L���S�����u��?T��nT  @ IDAT�SĦ��w�0���B!,�'u���JJ�A���ni#��5{�2"[>H�p[��!��h?Щ|~��4�w�m�ɉbhk��{:u�`�F�c������h��`��D!Ņ��ݷ8n�
�z��˝���;?�Rt���z��p�UQ���y�����N�����7^z�����.͢���T�J�mTQ&lHӔwtIq���gF'Ƨ����_hnjֺFM��ξ)�����}�~��8��W���恃��MA O�� g41,�2�F������;o�K�3kӖ��E��N�ŷ���N`x���w�ۙ��Ќ�ܩ2�0s��bp�ݑ���m���v�V&�)�9ʙ�)�B��K�l�N�ap5n/��_��h���/w_�~����;C�Ӓ�v�Lv���u�����N�����}�V�X9�������&�0���!L4��m{I~������w�_��~��t[�r壗\r�O���C�@]���W��ɗ�f�
�=�������;��gb.�	Yu(;Z�V�Z��y��k���%ı��d��Q�8��)v�	\�B��c�ar��xǀ )NSƴW�Q�!��?�}��G��%���b.��V%�:k�Μ���l�pw����^+���"	�r����K )��R�oվ�/��ހbA����zaF�,�k�,u���_|;:ʤ�وd��@�ӎ��"�g���G��m�RW��R�M�B������x��}�Ks��5xGA�Y��0A�t�\9 +fP���/F`�������'���%��ft�Դf���|�Zt���GG&�	�z�����֎����O����#lW��W�닢e�𫽇���������ʛv�e:ʽ�R�J�����#Q^�;;�K�K��I��z��fu�4�P�)��Yf�n��e��ѝ�r�W*�q忾���7�O��m�Gm���/K�ytd�=%4�5�7�7F���5m�W=��ō�+#x�n��nm�ak�$�]8ų8���$nV	��W�N6ͬ�`=���J�ҩ�����
g�&w���s�fPU����Cx�m��=d��K q���I���I�OW6�YwMK�6<z��8N�5M_���,\?�W�;��� \���t���;Ep�ڵ��D��;��p�'���z ]Z�܄���p�-��~��/������bu�P��YYI~�r��ˮ�,1
�Xvm�y��z�=�^��թ)�<�1;���כ@�o�^������ft�®�c�Һu�N۳˄���'/���f`rz"�Ҟ�*H������˿��Ҍ�e�����\��C;&��<���Q��i�j�h�L-|���\MJ���:�V
�פ��G��`�b�ߣ��D���ݨgI�����wt���״c�J�=�����r� n�n�P�P������
�n�D�]f>��.;����M�����R�j��H�m�`ݱE�PS���(i���N��Ӿ2M�N��N���\cK�<��L)�(�;��"J-�v���G���Y{������\_G����7<�{W�-�M������o~��;�����prH���C�.�u�ajtX�_+Zx����OiH�-iش�)iFE4�Ynm����K���碖f�7�t�����ê+X�E��}+��J�����E��E�#r���ƿɁ��	�IK�$wi[KޱR?�&�����T�T�)����8l�N�J�Z�3O�~5�w���qf�F��l70��p�+���@q:G��K��h�9��Q:s䈓p�;��&_���܊[��O���qج��%��L_pV��	o�A0��-���D:�"4�a�4�g[����"�U^?x>p�;�4�<}��Ǵ���g���*/u^W���k]�z�%V���K@NVx�������|����U�ΔG�C놣�+W�����v���~�6�p�@��)rN�A!D�h$H��C�i&���0[���wRȞP����������/=���?����K�����j���~�O��ybԫ��غ��%����Bu������/���2g�
�*��bͦب#�HF��*#���Ƀx��7���r�0@��6��(-���WC�N����:Q[KǊ?8�D�Jh4�
F�դ�	��4����P��=�N_H�p�!��Ux[-�SR^P�tC�.��\�1*k�ެN��4����5i�ˇ5�:93E��Rp
A����ѨA3]M]�qC[>�w���;��mm��7?�=<��SQQ�\l^�&,�I�7/�/>z(��ޝ�a�h8z�X8��͡k���[4/��O�����;CW[�!?[,�\x-��D�(��\!��.۵/��R����y�LKn���8�<Wyׅ�ag現��G��k�׿�UWK�ꄧK�f�����is�y��'mʝĩ�/�� �*"�',��Z�a�M����$�-=h���ʶ묿���d�<��8=��$���x�>%}yx����8	����i5�Y�=@�\z,�o֝�'��U��)�Y�-�q�)�4M��0z�<$�Y����R�)Mĭ1Y���%�9W86�Ӷ��-���,d$������>�9���M���dX�b<�J��ˊ�߰a��[�>�;��W�UG;����J��\���C�% �@o�{�W6�{��ӟ�v�;��g�b�N�SD#]zgG����[�}���q�a�&�KP�QS'.e�>z���}�)b�|�k��Ӆ����A�ĘrR��4�s��nx�_���.��Ol��2�d���	���P�YN��ق!�C��_(xf[��C����2)0��bu��ͪS�����XB�d�����Ri-US��Y ��I;�n��(��02�ݒog u�₲D}���u�lg���.�L��e	����Z競`u�m� ��.+6\4���iSNSM2Т���ʥ�Z��H��f)����sh~Ы2�r���f��7=:�:��X�y���ηP��W���Q�������MI���G+o�Z�\~�����{�#3����²��G[�ķ�g~��{�G�9O>]rͶ0p����i��1���SZ�9^�{����*�,�A�N������u��jD��xqT�1�2�Ha��YS�6��ڪ��[5бUu����b:á:o|���mPe*��ݕ�w�q�u��v� ��<��%i�������>��5�OڰL�Gڞ�����e²�.�<5�Y芻6�����p;]���m���ګpɯJ������  �u+�*#���6��?�,��v�g������j�ƍ6����T׭� M@��Xr�ݖ~R6x/��#;�����%C��X=�7�I[^�n>|	ԕ�_�uo	$���뮻v�^�o����0U���m��	s6�t`�-�;�l�l�p9��)Ū,�o
#t�!�^+1]�3a��t��0:l�ۚ�D e���&\����(?��(Н#bh�0��[$������#�6���͔��uJt�ha�b�����LD�|�P#%�<t#�����ӊ2B�'73B:1���w&�+�t|/�>��?}+.�L�g�BLU�Οo��h{�pX:d-��U[NB�%8܌�����N�Z'�ڒ�JҰ�ɇ���ޭᘉZ5��di���֩7�྾��Y-�����5z8z]d���m��
Z��y�xh*j�]��h�ց��Ѩ����D��I����˫FFO���R(�t������M�����b!?�sgt��V�g���a����	w����R*��o��;Bے^�}�A���^�ڀ�KT��qԬ_z��|gs���,�i������UԢf'�Q�Vy�g��k�?�&�՞6K�����z��y������7f'�R­Q�uUiy�&�.<����
��6j���H�k<�$�N���0l��vO{��i5�a=���������~���k�x�ۊ�i�3nK��`<-�`�*E��$��Ml�0��5�)�h�(/��6<���;f��p�$��_q-�LYz�S����n�_��Ƙ�"��m˿vcݣi��d#��@<����yz��cp�p�9F}��!9旚�%��V2���\}�2�c��J@�Q�Ւ�{�o�<��j?{��0��j�Q�_�Nӱ%~�п��>]|z�f8��a&�jii6��=G��gw����`lc?V~�y�
S����t�L�h�j׎;��i�&�m��?�2ɢݻwo��e�}f��������`D��8e'�:WW��h>�O����ߡ�:��	�+�K#��
h{�##1���-�vI����p^��Q�0�?f������Vf���2}k��ؤM=@q��������x�Ąp�!X����4�.�Ռ���S1��3��/Ek��,O:��f�h_(W�:K:%ph(�u����Nh#Z8��Ff���7�i+Em�]ʵ6��q�ҕ��{%���h44-�8
�W�����������ñ_�2.*�WEk��[/�(<��ṻ�Wcm	�.�[�,�+�j�j+Z��R�I�'���̜.rnl�骮�H�䄅��9�bb|��\>���\�V�{U���L9E��`Y�:+~ZTת�ݠ%����d����#c�LS�RL;ʼ[��wo3��mp��x�e�xϘ
O��%���iX���I����v���=���$�����ȼc�S�O�R�<2���w�Iӗ_U��0��OI��Dg�~���m鹿�Oޒx�/K����ka�q˾g#f�IS&[�y�FM��[��a|�z>^�@:���i���ځ��p��7[�s��ws(��	&ۀ�����yģ�"��,�j'����+W>)�jLiy>����K��\}���G�xK@!�ƿR�Ս�ww�={������Da�R��\ߢ�X���")V��7���&�C�b��-��F���d3�8�Q�kK�J��+P&D�a[;C2�XiM�I�688x��-}]3G��h���%`���Yû�]h�4Kר2L�-��u��K@eI�qI�*�|~Q���R8�
 �G�%pr�����Pl�P�툥I|��S��Q�WՖ�dn����� �R�eLB$[��n+�� 68,�����<�Q�c��P�0z��P��G����MM�b�є<�
�⣠hيd�����+W�ͅ�Y'XOjVox2����Mh�H�j/�/�T/.7EM�|�����PikV)�6�Hy��ʍio��jP��߰!���)�S����D�=��0;1֮Z�W�W��{�}>��������7]�.�P�htz4��Ў�����5H���u�Z���9T�q�YˁU^q��������7��0��IZ��RyV�SPu󉕀���G�5��_S��UX̣.*��2�E���.<zs��6r:�i;zRx����9m�_:�BƏ��?9�=&p�Fw��� k���!�z�'�Sh��a;H�8��fiM��e��w-�K���*4`2v6^����-��a�θS<I��{<�4Ǐ³�����Ii�h��埅q��	�\��K�׷�o����e@Iݰ�d��+o8EP���͛Air��C���w�rE<����@��B��d�/�H��c``�U��y����r�d�GWj���z��������x�Ν��i���r)��u��]���q[K̾��2cA�������h$�if��#qlǬ�H:��tttBr['�0	CC��f��0�d�!fzP�����{XAO
���+��1Ixmp6��)#�%S�ь��	ER�S��F[�=}	4�����}Y'5�����u��$7��8�&�Q���* ��z�=l��>��NY�6cJ�cT�p��P�F��)�bʎ�M3��ɿ���Y8�}��(tQd���?Ő��/�юRok����htt$9�<b CK�in֌S���`,O��VG5%�C{Sgh#�Q���8�uQ����L��1�XM5j�K3LSZ�8��e��ák�9��lCӓ���3\|q�da_ؽ|yx^{�~��0��[��;?,׌�u��_�&~�G?�����*�'�� j���\^3V��w��֬ �-�ةL���Hǵ����xv��:9<�����E�XE�Oz�V����Ra>=�ӯz�E)U��v�,�I�푅��*P�U���e ���lОc�wk�^`��#������|S��w�1K�Hr�3�s����#m���4~-~�/����<1i��[z ;}O�I��]v?|���`<	�)���yHl����E������ ��L0�0�-c�~Ǘ	�8���n�|b\)��;n���1�q���<Q���C~��e�[������A�$>�}��X�����@�ű�:�S���CP���J��G����^A	��ٳ����p��?�%	�@sQ⬕��.;;;�Iq?�>�Z�Pa`(��\��8���D�ni�1e�bL�P)�B_l�-&a�Ƀ�Iz�[������wk��Z�<�xU���47����(�t��0cc����ډ�0]�/�>Ar?�I��(/�S.����[o]%e��2�l�	���iS��R�]Tʷ����v��Q�,��n�4��̓
���l�BDe�Β:ʠ�<,�c��i�J�|�H�n	��W���x�Z�������}ʒNlc#�ч"I�#4C6ʟ��+:���T������.����Tr�Нo�z�Z���"�u�Ɣ����T���O�Z�Nl�-�a&���4p���Zu�Eo{A�*[�c�����W^�ᒵ���K��>z�g��?�q|T�ڿ��_��Ɨ��o>̛uk �Y�#ˋ+��$��\8��:�p���!er��m�����i����������Q��X��U��UR�:�RCdY�:�����&�&�J�Wܬ�s��L�ȶ0���82�gv�O�N�x��흼��0I:f'��L�ga	��:o��\�Mi!^�����3�a50U���^�+$g�[���8�N�_�����b��fݵq=�Z޳a�����ڠ4�0b�ק��(�<����N�)`H?��;�G��z�}�h۵2۶m3�h�_Pݰ	W�����UjK���ztѢE��ʛ4��#�\���ճ�Y+1��f�n�b�?=��C�엒�-�Ӟ�[�ؒ(�������>�ϠQf�I3"�lX
����W��M��NWL*6����)!¬���P��Y[r(&VT�����;���v)V��}�{.ԙ6Сf�2����S�˲|ݼ�`9e�f���ٳ翕�Ы��1�9ֿ��r���,�����zd3���ӉtM����C�J�	�M�y��n��m�O���:m,`Pd�A?l�TREL��yq\ēBd��D�ĥ�`C#m���[M@'F�LU�vFBiKġ�ѡ���d�N�����'T��M��u{�ɢ��5N��BW�.����}��M�� %Ox�3no-��Y{'�u/Vs�����UF�f�.��F
�����{^z%W]|Y4�r0\�yM(?r(z��G�}��xJ1뮸$(,>x�H�,�W_���5����tI�w��4��DS��ʋ>q��,�"�����%忮`����m�7L�E|�"�ſ��9�bET�g&ٮ��])@]�=�:E� ���./����L����d���+^�~B��y�������
����0�{�Ǘ�̳��~����L6���9�A���튕�?t՘�Ӝ��;�$��yz�<Yx����V�=�I��;��$͔�3�+,Mw��L������xɏ��m8䶁R����wჃ��&q7
���_Ë�w��f0v``�;�~�Y�'�L��Y�������GV�uD����������|�m�̓��D(aD9�.1˖�uvv!�ڨ�K�m��pxB����wt�K�lQǊ�i�X#�ib�iTǖe9c#=	���_1#CO~�k_{\�߭�u��O]����Q�3:�#�H��O��4C��ؖȸ?�rݼ�P���y-�&��4:~�f�:�:++J��2�c�w�@��	C�ᡎ�݄%��<�F�e�.�������?J8�w�����Y�6�3d��h�e}�	.ff���"8S�	�ܭ�v�rXڑŭ�W�.���i�t�t�Zw��J� /*���/)6�Jq
�UC$�Z68_��j�c4\W]����Gt��2�Ü�'�8�ҼhVGķw���&fȤt�ි�R>���M��iѢ�v�ua��9<����x*��ɨq�X�7�5�q����hx����ɩ��9��i�Qo��� ��#GB�N�nS9i�[����F��fX�ʥbԮQ`�����Х29_��Z�ϔ���v����%�T7y	��i]����[ܪ}V��A��33V� �Z���r�"�g�_k�D�P��X�Kܕ�ʯ)-�ȸ] �ت�P 27m���;kj�-}`1N��э����9�)1$�?U���7�Cm��%�V�]��"���a����yM�Gm���Xja��ew��+�4���	���=c���]���|��nW��;���"xK?���o�A+���|x������+~mr��Z�W�pD�;u%��BZ����#����GX�uT���]"-����#��ݝw�YS)�A���G8�
��}���g���k�+1*q�xn�cG,˜l��������	T0�㒍hp���'���꫟��[~*���;k�����A��B7B64�c�ʋul��p�W7�T7Y�@#�WK���RL.����RJE��PT0���U:6��uД�-:Rʞ��E���������X�ϊ�
%|?����?��Ұ8(]��&�7��tA0#�2�
eKG��%z�t�jv� i���*��Yʓu��s�LA3IT.�f�H���S��4�p�E��U��s丝ب8����YgKNډf�tߗvʄB���u��L��L�0�w�t4�֬%��rO��]3Q�Nl�Bk�՘ă	�
6-X6_}m� �������:s"ڲzq�mY���4Ȳ�J�˺���^]�]���J�X�� A���!)��H+,+�B#)Bv8�_�8�K��˲eMLhF�5���pA� @�b#�ht7z�^j�W��}�ݼ}�����@w���ֽ/��9�'3O���Ƕ_��P����ݭt�h�o�؝���:A�U>̫wa�49֞�toH�R��4�7�&��j3X����}�2�c��|Qn�Xֺ_����L`��e0��h�wS盶�`�#�b/���6CyF��:'QY^`��dg��#Lv����λT�Mk���3��h��	���L5�&�n�e��5<�����QrZ�����;8�������8s��^���6���F:˴F�z���.��a"�w��|�;��^�2�J���]�.Ks6�k����(+ӫ�)]��2��#㯋��zc����3ġ��*�� r=��I\��8���6'��s��W��K��_V��_WWq�u90|����~��c�������RÅ@�p��-��G��+.K��nu�8�2��ǎ�Z���1��A�_�� �c�:
&�Z1E>;;�`
�0�ƛ	V���G��R(βY� �W<}��w����(g�6�4"(Ch�L��~Y8�=:�l���r�N��d'ס�}f�޽_F���b���A���η��a�q�év.'�.��:�- f�(Ǭ˲��1�	�:�3Y^�[�5z4��4�<s���:����e�����A��Y|v�:�c(�<�61>Q���#�i�4�XzK584�F�G#mg1� ���HO����*/���[oE��G�Ӵkt�=��އ�wb~2�)�R�o0�{�!�`oU���(�M�fi�����%�@c�=eSs�,�N��pK������d��#oRZ��(�#M��4����wN�N��6�����^������-�g~�~2=Y�9~4}��[Ӻ+֤x�8���,A\ρ,uD�����֚��h.�-���Ϝ�i�<ptW�f��5�E���Ä�iG{�E5iwONO��}��r��}MN��q��N����ZDۡ}���ضJW)��÷�%|�_�x	\5���.m4�pf�͞=����/�pOd?e�������K9���$�������Ӭ��8<n<\΋�9A�p�g�����a���*}�"O�<�y5,�V��l�eXv�(Ӛ�r������4�S6f� F�eD�+�뷂N��Y����*�ґ.0��,7ë��i��Z�9�%�*-9�w������]�m\�����#�R�>b��y�0���8%�k��c�dp��o�����+W��p �����G�}��������x��=}Y �o�}U�{Æ���)�ڡClB� M{5�a��6FhX΃�Q�,T(���zb�KK��i@�P*�
^R�UAܽ{��/~�?d��kк�|P�U.H[�N%��|��T��V��i<��r��w��\���M�P|	C������<����O�thvX5:O�;�#+�ǯ����D�E�G���`1�ڈ�1�q�o���R8P���u�޺.�8��u����/~�vS(<y��G�{�N:yFKC�aL���ĄiT'U�f�y�0�iP�h�|���H�����ЍNV�hz��b��w]�5ř䧗t䡳ol�e-��~f����f-��T}���b�ɼ�`��ŲBN������vcj�x~�+������k����Ŷ�;�uW�nw�����C'O�S���{�7}��+�\c.�<6��p��R�ͮp��r�����qf�z�e�����G'�8s��Z��Mr[k6�	x��� pi��5�`���G���#G�d@���Y�Q�Q�cP�r�?������a�>�S�N�.ǯ{W�VOqe|%�0~l�RX�-��p9�8�x��Q�s�
ؠ����)]ݐ���8��7�u�t	o\�Z�!|Y�k�}��٨�q_\A+��_���2C��9�������9�a��|���W�_�"~N�~�o~�����2�J|�ʴ���w�[������>@���)�
��xrY`���b��}V-�^���G��z��9���X5���x�����B�;���s�>������?7>��S]]	H�
�:Fзl�Yx2�ѣ��iF�<=�3"�	f�
�$
 Pb�F��*��q+�\��J�#��	�Pf���Էi���9U�ߢ������{�1��/6����9/
���.�~/y�Ѡ~Ȥ5ԵO��#���]��\n�>�>v�pg�4T�;�H�Yl6����l�;�Xߨ�Q��zq�]1  #~����}�����I'�8�0���rv�t=�h���V�q����G�;�=T��M����/�<��6��]��"q���ϣ�5��~S'�в�FM��#�߈��Oi��WK<�c'�n�9V�4�О��e�B�gh�`歸��;Ӧ�����p���J�o�"�N�^�}[�s�`�Mfÿ������<��g����SktM?z&7��6���q�9�&0�6�mb����U�l;=5�8�o����k>3�qlo���z�O&^"��놅��4>q�7:<�`��KK�F��ۑ�B����8�W���]�#ڋ��x�������](�xde>+Ε�-�_���H����L��& �����<�~�ĉ�o��qJ<�'F3N�6���D;ˇ6����>���'�qtuz�+�;�g�-˛p5W�����?���F��w�J�+`�_�����0ן���5N�S~�m\�<��.��_'*|퉼�[}��~A��V��~��W�Sa��V�X����#w�y���y��g�u��B=�߿V��_�}���c9���X�}|�����O>�̨�*�T`C �����l�첶S�*v^��2!�*F
�2��F�B 1-�(.��y��k�؟Ψ��I!(��
@\(��;�!'�y��P/ȵɤ��,���
�YA[)�}p���aW�Y�x�aT�¾�/b,��#~.��o��w-���������a�uʷ��o���|a�+�������G�h<�V��'N	��u���t�+\�GZBqr�B��6 �,�8$F�T��w�ƛ'����<o{�_{�5_�5�>��oi:C���
9���?/���UGi�� �F��9�����X,,<������p��e�=��&gg�Yօ-r8��`�~����X�W�o?����+/��O�޼5}�;�.��ǎI�}�������m<P\v퍩w����̐Ϸz&[��E�¾�F�q�'�����(�K}���9>}*�6�[3��H�g���X�����G+����?�e��u�4���Ÿc�FC]Ɇ��E���d#&+ù}F����,�l�!K�:��N�������;��p��rQ�������a5|A�o{�w'V�7ӫ�|­���-���,�ea����"H��-�r�+�-0�e<�1Q��߸���a�F�?簊��<��y�w�WҨ��(�����*���o�f��'�C�Zf>8�ˣx�'�/�-�a<_��D]��шr�����q�}�m��-���Wo���"��������5�U�����U��� B����ܶ���y������SOoҮA�C�jy<B��bt��u�e����FV���l�A(�y�J(ke����O�ɇ�&��ʤ��}$����`�>�ѵ�cJ9�o�t��� �� �UIRY���)��(|���\���KA%p�S(�V_��(f��Ct�տ��ڪC�hX��K�E֝Y)�>q£������:�S��W�[ϭ�	�hC��(�ƛF�0&v�Ґ��?��0�,�\��!����q���r�J�ď�!��D)���,i�QVg����=�ƼE���ܶ���Ҵ�Y/ͻi�߽��pE�5�Lo�c<�fZ��a�A���`���X��1(u*K�LE�^���b�`{C��-��D�pq��P|��t�G���ؿ�w�ï����f�G>tuڶiK�ev����7���b�x��J���4j2}�Hc���7\���۳\v���ĵ�#�x395�n�����}�MMO�Y����!J6=C�&,�U�+q�r������7:|�I���P_�Wf��:V��#{���p��w�;�>���C1/��[�7�6g��*5��u!�4m���/�����>Ye�x����̏��p�e��ez�F���ϰ���]���]�̀�y�CCؒ����x�-��oq�����c�|f��-�e�|i������6����!Z�X�&���k@�<��e?`��&^�_�e%����;�J�˃�{�9�%ua�V�T���ܕW^�]h�X��՟��W����|w((|�ͽ���_��_��_lA��SS�B��«ؾm[{##����x�	Q0�t�a��b�R�P�$����NN��Ha*�_���9t9�,�u9;��x��k��Vau�Su���IoG[~�l�_!]�Y�PX��;��Yne��{�E� \��|W�e��Y��!:���۷�K,�ài]Ұ�p�C���qiht�|�>�oa�{�g�"�L�w�Ky��]�	�SZQ��G��[#˴P���i౸cL#�8���oӠqc:4��`�zկ[��rFC/��z�����8Hb~~.fu���޶mG�n��g�x�Y�n.�]�!1�
ۦ���i�_�?0����̳���g���e�-������ab(j�a��wll]���4��..�KqJ��O��`�-@�ˈ�XJ�Z��g�J�n1H���l���^��;����N��O�O��6��}�z�6mM��ؚ�_9�����W<?4������^qe1�ncZ8C��ս��pS2iqz�8y�T����g�%�k���ho9q�ĝ���,ri�������j{���W���XG��:v��C7�:}Z�Ŷcq4�k,���Yֿ���N�6j<>+E�:��=���ҞÂ�r�@�h��w��qt��q�K,k-�+:��p�+�U�9��6�}�W�z�+i��/ҩ�7�'e��}+/�S5�o��*Z~�^2m�u�4�3p���w=NV���90�9'��/��-���L�wv���x�`Z�]���Kܑ�`_g��p����)�k�t�}�՟'�c��?(ˑ��@3<NTWz��[>������~�vc�q����!?EW8�U�	�\*V��K�$/�|41�.�?��7��P
��V���g'K<<�y��<�Y¤�����YD�h�H*�PV�i;�����
$]��"�:�
�����Å`���G�k��3�x���޽{����?���Q��/鳃����S���3��S�����)�K��!��s�>�ox"/z���������q���E,C�RO���0�����Ug�yo��|�|b����с��H��$���^_�I��i������/=��p5:��\�k]���L�@�X^�U�r�ǌC7���ٹ�G&�q\n�訆�{��_������m���c�#�p|{����^�Hs�?)f�L��y0�څ<1��v�/mt!�\`�y�yw�U��i�ܝ�%U���XK\z�i�����*��������i��]���ϟ��<�t:��w7-lnoY�W�36TL��Jz���L�̥���|!]q�u�i�#G�s���05�NL��$�Y�`�����o��3�5�]�E�D�@�a�q�gu����5��J]�3�[h�^��cEGL�B�/Վ:�K�G���/3�hO��l�u��;���j�~��1?zv�x���t0��I'��a{��8+�?"/�ȍ��?5�:ފ~eЀ�9��/��l�5��2��w	p~��ꆆ��H��xNK�&�O�e��K�);�8Jw���X�����ZZ���w�_���Y��k��7�L+��#_�q�������-�(��Ӆ�^�=�X��?�y��i��j�8x�Ƹj�u�]��J�]���:Y_������q����*�w� �e/���/������#G�6�uBX8�J�B�Qq�����޳g�£L�������.ڽ�3�V2�sW�BLe3:9b�s�W��܅�T���3}L����j���P����[�V'DՅR�М�Ύ!�F��$*���
g�� �o�&����q3�_Đ�J�C�ڡadi�2�>�����������*��� <���0��}�/:Q��V�S������@�#��Jt���3C�i��D�+q���m(�p�#�#�k8Z}c,e��F�ĒE��0��aIz��;r���p��TǏs0#�%J{�}���qͫx�a>�����2րAYN������2�4�]����4���ì����q�e�p8u���n/��y��t�'�K,�
gL1��]]��vc���O}:ͷ�ҏ����<���'��6��=�3����_��!g�����k��48�>:��y��_����]��A?sz2M�9��o'�/���Ԇ�g{���?���U����8� �w��%�WR�<z�Q�h�-��,u�c#;J{+�/w�F��V�L�1��K�e���$c2�#�7�"l�Qԅ7��,��.�E�x��߸���cޅ[���4-Ksռ���xW�7Oe�����̻�]�Y�
�����2�a���j+�5??+z��6�yp�+�d�w�!�*����s�3���d��Y���Oi~>�,4�z���'��F�����驧�r	�{cÐ��D��i�7����o2�6t�O�|�W�~%�W��V#�u9��K������˟���(�t0*�.�s���#GdX
���w;#��B�r:11���	� �NN�c�����t��\a��?:"��/����5�\��7Ϛ��x�a����7��u���s8ڂB6��)xU�q�!��'��|�5Tv�����T7��&����w�u��a��<�Ӣn�̈h��S�-.�l��4�4(�X���3���FP��u~y��q�k���S@�a�p�����3��$P�  @ IDAT�1\�XqJ�����O��,g��/�d�w$�֙�i�������;``M����i��3em�:�Pm�]������A1�
��[�ˑ���1���j��7�M�7R_��c���|�1[,Ol�D����ba�0f���H�u��er�@oOw�q��}W\�\\��\���6q�
X��R��#�o]{�w�,~���O���i~j"ݵ��c��4�5��83[<���,δo�����_��v��7����5ñ�k���4���u�0;�f��`Afq���۶M��c�UW����j%��Y��J��]/��s��H��*����WqϜ}A(���l>ڣ~|G{���3�0��<����oqă�CM1�.�;�˾�Kx\E��(��h��}W�����Jt�)��r�8�_��W�%���.���˳x��m����2�'�_ʒ��(�Mq��g|A��'���(���LG0�����+��׉çt���Y�3=�w �i�~gx�|�y5<�@��+��5��w��W�'���%/"���q��i2��>YW������/�	Ke�������>�6���+K��� $��Y��i2s�<�-���P.�t)�U��R,�0O�ѷ�z��������Gs�R�,J_�#�U
'�[0��O�>UpR[M*�
}/U�|���
%�i1�4FY#lxx$FΙ-�u����pr�LA��i~�ck!�_���'���7�t�[.�	�y��J<YTy&?v���|f^�;:�B�?;=Z������F:���܆A�������i�h���޹F,xl}�>���iiبP�@��?�|a,W�"�)�v���(?N�5���������$g��#-�-og��[�V1����
�"�@!����|7��i/��t�FR0�	���~t�^Q�wY�AX.�:�Q�R`�2=u��J��j�l�m�8YF��6چ�0���o�3r������3�Zq�xۛ���(��+�] r̅��8邋d�u� ���V7"ښ�%�KXLȄTw1�i4]~�ui��;�/?P���ÇO��ʹqxMq���4�^�?~���E�"�����MA�U�uq<��g�̊E����ܽ�4�5G&N�L�G}alÆF����)��0���WG���+��n܊̾���;�l�!�kX�pў�.��wV�3��;�G�J��S�&�k`�L�֧F7˃�oj��F��L�V�O��v_)߆g��s�}�T�3�������'�����gx�wͿ
���7O�5^NS�e��߾Ww���t�n��:l��O�V�����mx��2���|Wy"N��S��H�zx&Q�_i��7���lNG�De������ߐ��Me=َ��|����\�^y�G�Ǫ�h;md�FW�#�O�v�m�;'�~2�˒���ݟU�����£�#����7���}������Z({j���?D�@	F���S�l�=.���.b�&NC��B��0RP��	����ʡ�IE�0.z*�*����'?�g�����0k��	�����U ��Ҹ��Tؖy���O)�3��v9���_���{����o<���izvf�5�n�K�?k+3'y1N��W��Uu� X'}�\��~����a��� �=�,u?�#�{9��S]�Dz�h�Hs B�`��5��r�~���	��4��l+�U
�96Mg8����°���ٖ����jI�8l��O'\( ��p�L�84�l�9=��i��{Ba6�($/�?��2�v1�v7FSd��'l+�,�O5 h��o�s�UR�����,4Q�0XPv�����|��C��7��x��'R�ܩt+���v1u����o'=�p:��c�uW^��F�ۓ'&���)5d����ӑ��b���~�I�J�ĩ���;���@��<�	߇?���#���jڞ�y#u�bl�%���,�z톲�.�X�TH=�"�[�����(c���eq: YV͊x9\����
4�3�Ƃu9"P7�i��4 \c|��>q3�@'^�*������,,<kr�2�A���o�K��S��p�sZ uvQ�+ �J[��ٿu�g};F�3�ZP|��HW���LG����|�/a��2��^"_�0n�6�xU�UK��Uڤ[�I�e�5�N>���_���E�G�)���hdk{[&~�4��l�ǰ��6�N~�ӟ~�����"Zu�	V�����\"���~���~������Qo���㓣3P�bi^;
�#G3ku\��醦U��+TT��p��RISN��8��.f�S!ԑ�\-j������t�UW%��N�?�����~��~t����٫���d��P�����;)������;|�>XG]�n\�a�0��ǰ���c��I
]�ގ/�,���������8U����ֿl���x�e<�:
����+�uı\M�P;3d�"�}8q�&g��a��
�Q�g����O6hY>��aȘFG>�9�]1�u
zK�$�ҙ�u6*�m�^ڞ��-�\䑎?�o�ְ�w�A�62Jd+����Ņt��Q�g��:�� �%�ӫ�����8K�pi/K3�Y݇57=���*x�E��c�.2,0ўި����f�#�t�
rGM������b�h^�3�ѳ���,���kό�׮)�&����'����Lk*��j�Ϋ��������Tڢ5�RFO[\�ku7M.��4��,�ٳ��FvF~n������k��q�Ъ�sV
RW���}��vF��ڞ([ؐ]�YXw���Rʵ,�4���"�J��G	W�?~׍A��f2��+�)v^%�h�~���>�w���yk�P�B�}ۀ�Y]��h��$����io\�~�jv��*n	�ez*Ð���әaK|�!V���U�������7}��w�,�������X�ξ=�2Os8���0��/}*0^�60���]�_���EYV��<�y��{���,���4�*e�rV:�U� �p��Z�6
�غ�J؝;w��g��=���V����Rd���U��=f����%v��=�Gt�K?y�^�y�E�l����A��e���Ŏp��;'���������K�TLKA��|�#�F�J��F!F'����"��L��_}i�����иS��$��k�v,2�^�����%]�o^	�ND���c��y��:=o�~p���&ug<|��a(���0
�S�iG&/��c=�̃�B	���[ٜ;e�.�i\爣#��x���[��t�A��"<��8�#}�av�\��t��KG���0�X�74�&�Xrі�mK�Z��v�`G� �����*4����D�7���q����4u�;X�۶�a���I�|�&mY�z�h���F�x���A�������y��qI1�3�w�����<3�=藋 e@�����y�X���������G��k>���l�Y�4֥�������S?N]�)���+m]�����>p����NOM�IŽ��[�H�8xPŧ��83~<�L�n�߰�}a(��{�������Xkn��L��2�w~<F�=0ǲ�@;�`9o���K?�a��2����s�!嚊3
;u+ױ�Px��4����DXeX��������w����L����G�,�A��0�Z����p���(�`�?���:���۸<9�%���ĩ��	[>�[��3���o�+�˸������{D�Y�[�}�J����*������'�K<9o9��nF��Q�_�get�H����y��z�����)���_���K�틬��)����U�,L�>���Tc+�>�1�fƪ���{����=��̪'z���ʁU�����.�RЬٳg��������ER�/�����$���J�JR��aTm۶=C��q���R��0W9�$�l
�R0��W�@����[oI7�p�a�'�|2�$L��8��;����E$���G�H/�rCE]A,_p�3	N��B����a���:I�ێ��Ϩk�Ba��'+�A#�\~�l�F
�+�
���p�B�`�I�sot�*��v��VyΙ#��a���2XN��`�E���c9�N�oFR/'��p���/�����i�F���Ɇ�MEy�T:����G�QF�qM�#����֨3���̛u��
�a��5��S��xO*<Q'��SI���#R��։���3��F�i _�r�^J.
n-���E�j���(�母�X`Y ��B�^��ǐ%�%�l1Ȍ���Ժ���/�����������<:�>F�8}�Hz�G�ˍ�nlk�r�G���}�c'��3�S?'5������L�O�s�4��Ԛ81޷n�̺6o����/��6#��?�����0�?������;��	s�U��[
V1���J�P~�6R����2yiY���/�9����c�o�텇JY-�ڑᴑʈ���@TǙa��?���..�dӖ�2��(����y�h*W42.ށ��_�|�a�w��L?�!|��q3�*�9_���i�������#�č�L7����4�Te���e$�ǀ�O��oy(��_��:�F�T��/)cՃ��D[I~���#׭o�m۶��9�J�琷o��|����������K�$BC�Ӌ{ݷ����=��Cw!$��,?���G�h�3�gZ�H59�9�
�G!T:�Sg�a��r��[q�˓T�L*i
Q�qY_}�F
+�o^6��8NyǎqZ�S�{X��2�y���v���M��/�!.��C{t�0ʳ�!G~s�i�kN�- n���8���MV�ܷo���1 b���;4�uM#Ƿ|D����z
�~�?�F�<6~���,�3ܺ
l�#"fk3��uU�ᡓ~���#�a|c:�[7A�8t�qR�F����o��Φtsk�(%M����t�ۃ&h{a���Ԥ���6+���Pb��ݟe�	�ۧٙ�%��ߙ)�b<����f�\������ N��b�k*P�9 cn�%Ɯ�E�F7sY�d������)H�����a^_c�ii�GWO��,�<�Ǥ��u� 8oH;�3M-�N�4��^|�X<y"�B/Z��]�'�g{*=�7��_bY�7#[6�c�k�5��*�z{�%����4=9/��bff��>~�u�ٱc�	��y7�4G�ڐ�38t?
�'8��*�M��9s��%QP��>��Tn[�E{+��y�h��5�np5���4�wW�
��TxMO��I?��U��vi���7˒�D�o�gܕL1,���r�~�c��LC��K\��6,.a|�]�훼��/���7OE�*�u\|L��� .qd\�,K��h��#����kX�K*C'�(��iû����y7�;�g��[V��3ғa��U��M���(>��lX����!#��V��g�}6=���E?!����M�v���}�r}Y���3����^5��� Hv��n��׾�����#*p�fo�������X��`�K(j��8F�Q��[��h�#5޿��3�Q���9��煡�n�WIs�#��]��޽{�
n�Ql�0M��̗���Y��4J����lȻZx�w("(�a<���N�x(���2M��?Ȼ���cP�c���,+��З���Vvdv^	qP��ƅ�G�aᬕ�Wַ�)�g�|��G8x�H����@��^��Nv��eiY?�8�k]����ۓ�4VL+jM���̸�;���A	��6c<���6��=U.����_:�� ��y��4�vg�tR���~�#��~�}��v�g��w���q�.��vi�7�?�.�G
+/��7�N����s�S�Is�*}C���E�Y-�/��ԙ*԰�`�_c<=�tt�ՊS�S������ힾ�E�h-6g�gYJ8y��ك52��n���F��k�dO_z]�g>�����[,an�O��Mg��o>�Pz�+ >A9�x�M�M�.+N�[(N��^�c������8��M���ݜY�i�������&f.�W�%���̀yV��|�N���Ng�5���d��F\��̺�C#��m��N�e��j��x�K��o��w�}>�zx|g|�w��w(ڤ'�ix��TM������G]��w�׻�ϸ��t�S����_��_�A����#�m�4�|���8��~���X�D������"�%�ZZ��g:5U�3�v�����o@w���4V��3;�g�d��ӑyS�'��p�iU�r���G忲_��Q��(�����앸��Ce1K�ðR63K%�cU�;Y?&��2�z�J����U��}a��K�������G����Ƿ���k;Q�T<��#�d���؆�id� ���b���Y�t*�q�M�ilc�vŶ�0'o�9s*�ǰ��T.�b�����1�:J'w�V%!e�@�d^,o��ƛ�����O<Z���-�:t��菘F��8�c=��T:����FV���PΝAΏ�9<+�9�R}[Q�8H����������������bk@��ǥd�kF�(�s�c�(Al�a�3��暞%�:PᢎY�T�姼�E��u��n�X/��=����:l������ށ qi|̡X6{��T\:��'���Dp�ǻ���i�Hy؋��s����t|o޶= ��L��6���j����LA�Q��?&�2��P���|�V��\�������q���u��w��Ls�o�^cU����1�\��r<�B��BV�~YW�⻣a�O��cZH\Bhh��^V����0�8��ĔǾ{������%�ȃ��޴0������e9�����Ӝ��� k��N�:5S����+ַO�ucѷ0�����_K������w҆uk��nݐv#�����KO�!szN�@�a��Pc}j�N��NP}&��ig��b��n�bxtM���������ၾϬY���@J��Ջ�^=����l� �������#�>����O��p��1�HҞ\�@;��2W��߲�ON�uJ�r?~�X��-\I;`�����;�4<������:ہ�B?ۍ��LS��L���l�c�(Gt��4ec)���I�o��\��p�~I�#<�m�AX�9�Ǹ�����qeܾ�w�/�̃�sX~��oÄ���Z�w�+�����z��������_&�C3��4���gP��ߦ����#������#�ܷ
�o�a��L_��'��C������ԧط
o*���\a��`1s�I��)��;���4p�\���g��9n6S]}��X5��s�_�".�z��W���o|�ƈY�҈��A�`�b�ްa�Q��;�@ᛌ#�[6oJ�qr���#��Ȍ�ld�*:�P�Bys���BIeY���k��#ԦP���������X��Ϥ7�x#�8��ӽ�����3�x�4^�#��S���2M��پB���y�0ޖ	���d�K�M}�	�'���;�s�p�4�����|���r�ހ�H#÷�sJó����v�*9:;��m�O6^,;�bvf6F��Կ(�I8qp^Fd�G#�4D���{��g����1H:�bqM�KϢ������S�S��O�2G:9�7�+�9;l^4z�M�c�M���O����~��lQ��X����}W}1#�F�?��/���hm����<�:p�Bf~�m��oe�|6o���G?�dZ8�ܯ<�F~HK9 �F�"�^�ݠ������8`��L����@�RU���0F{X��.��C|3px:�;4��O���X�OH�h�׏�����|��m����u��rXG���� 'r�x��C�M��?~���_"�[}�y{��^��<Z9�g�9ql��<x��'N��������Ҳ�xy�)�&%+�X7�3�.����締�o��ů�iO����������a9M|���5�3��V�k�y�����V��i�w�#҆_�k%s_f<
�"nE?Ө����w��V�xyg��t3��~��f���;�d�j��|S�sE?�5Nv|��ɿ}�;?��Gٕi��;�'�a|V���x���/��r0�����x��/~�y��VN+�p-�&ɛ}\!���o~��V'Xu�/V��������(��3cu�c�=6J���c�]�AQDX�4�[�CT�E8�}r�U��k0��06٫��(�����eX*)�)��q�7�n�XJ�_vyڼyK�����Vz��gb�\Ez�\�:�[����ċQ��Bu�*F#���r�#e*θ�=ɻD����+]��m=2q��}��}���;]��A�m�vgf��U,q/�](�~��eߟ�J<��aoy/�ʽ���"�Tq�-0a�`|``u�n�O	벿��Æ�3ZFЮ,�����ƕ�F�o�a�;`�X8�9�Q����0�
N�<2���G":��!)-T�Wťʱ�pv6��)V���>#�����4���K 9���@�(�b/����������8�����zn��[��o�G�c������6J�!��f(J�����}ũ�r�FWZ��F�����CH{ar�XZ� �ZXIS۶�O�q]q�g���3���ڮV{l�pq������R��/q0�d�Ě�~ۚ4��,���~��GlM����aC=�����ﮅ�y9|��Ƒ���6m�+��M��C��]rd�"�Cޔ9���?��G���U���XX��yW^�p�L��緞Q�}�|�3;q�X/x�����8�ŝ_��)��M��2�����yWJ5�#.�<�Q��y����;�O�xPO�p��q�a}��2?*|�ٯ2@w����?�+���c	S7^�
Zu4��2�<�x"^�t�P��3o���</�W:�0��8�O&�*'e؊�A;˝2?�T�7L�(��[����M�N�ʁ0�1p W�e�Ŏ;B�B�+3�_�����OX��J'���������]����z���~���,���p����
!���
�j�Pfv��x�G�����ba}װ��RH*�����q�
��P�U"CH��)�4褽k�N��E�2�W�`����=X�j�ڵk�K_�Ҟ��� �.�{ ̎\��N"���.�{� B�_x	� ���GN�����g�R�̽/�55}&�V5��j��ү⯧|�����qd=��M�Z��$�w��_�}�Hi`h��>�0�%~�"N�<������8lC���_�ʹG}?뽏��:����'FF�7;��h���_�*��2"ݦߎ����p�����c���[Z~|1�$�L�c�h��I�s�1x"��*���ah��X(;�,"���6/�L�t�y1�y%���&MeE7����ۜAW�2[�[�.�� jqY��h��.p�X���wt����яߘ����z��{���uh��yamZ���o��&���{N��'�e6��f����<11�hF#��<�uX�ɩӍ.�.^e�|��U|���8�"�9ٺ$�+���Э�����ĉ��9u�a9Q1�G�QQ�:�<��Q���z�[W�u~.7(���h������q	Z��9�q���c���Q�B61��0��z��Z�EX6��\�#^�3Ӎ��8�w����oߺ��[���o��c��A��̓�4��|����I��H3������?ӈw�'��Z��֕p�-��F.s��w�f�U���[��Òg�i*����L��9yyV�9h�l�Q^
��cp-�xs���a5P¸��^ՓpWf��w��\}�:k%w. ������$\�@(b}������Ϛ*M*L(*�A"8B�mfo������:B��LW_}uڱcG�:��`�+�BYIS�6�T����O�<3饡m�g��^���֯������S~>���k�T�m��p��y��1N��}�o��Ύ����{�S��m��-��k�6���l�N$:v��R{������ǏO|��;~���Qxb�ic\�0�p�}�Fitd*yvnv�v�t��(���atr��&xi�}�o��z�c]��ebt;J��ѩZf`�kؘ&%4<L���ť�k
f���-��������'�Ƅx�����A�?0ļow��Xi�yP����x�/5L�?<	��aOc�?g�,. f�ɻ�<�O�i)Dt�����r	j��0� _���������0���z]�M���yn^q!���/�Q>/��JN`�Z�&}�a�3���s���4ŉ��s579�fo\�;��:ڙ��Mir]_{���������/vcl�8����h15q*}������t��7�m�����t�f�� vrj�yƙS���ݍ�	f��g��F���]=�{���<��/G���8W�NN��Ǐ��L,�eU��_�dWm|U��K��xk.�G�W���� �ū�T�Y��p��yY+q� �|g*�(�7��<�+�f������^6>"��<W�9r~�x��]��~�1NN���'M�G������3|���Ӭ�eE���k}��۴�tY�A�R.DT�	˴�۰�w�����:��+�"��P�"ig2%��e8�(���^����V�O��e^������J ���ݻw{����c��5�\s����}�����ɩ*�i[u�V������e�H��5���>'nz��cY~�Q�T	w�Bϓ5�F*z�Ġ@���
eOa�0R@� �0� "ϊ�َ`�XB@q�(��
�%P�w�H;w�T�K/��jz��WP�盠k5�˦���Y��>��?��d/V�^��C	�G3*����A�^��:�}���<�??~b��uNC��D��<+�YV�y[_�D;A��U~��a��	:a�'��r�0?(����z3R�
#};Z�h7,������s%�KCL+��ड�ဃo��7_.�wgE��3��[�1���3�>:�)�z(��7J8�9E�O�:�1Շ�4(|̒@���ߋ��-�T+OxsI^ut|1�u����Xˈ˂��ҩLPv�i�Io|'?M?�1s-��8���nyi9)3��/�iL+¯?�yf����&i�hw)�]aa��1$ќ��9ddOZ7��9�bӵW3i8a���/>�lJ'ӎ����+֧/��<�^�Ez��'���?v٦4�i+��7���Y8f����{���J���iϵ{�ٿ���O~���#����2i�T����������9y�osx���M��K����V^�3ک �W��ϲ����}J�������T�t�#�L��iT�4��,�L��W��£�Mo����s� ��O�L�w��� ���+��	�??�Ѿ��"��G+�o<ۣ.��i�s��W����7%>1Tq2:��hF<��M[��%L5��ӝq����ZxEK>��i�ַ�U9%mᲿi(����T.)�с#V1�C�b��Zp¨�	�\Ǝ�<�R=g�����	��O��s�_�#����(>W�����.�D"XzP^w����|p��4��y����ix44'�1z�P?q<�+�Q�F`�B�E��Ȼ�	!�VA�bˈ� }qt 
2�PU0u*g7�xCq�UW�2�ҋ/��_`�9��%��L�­�"��ϳG�к�Gz��R ��s�g��7���*+��{QzS�8��#���#W`P�����Nq�x{�]{�B�����N�'���[v�J��(O|/����*��=��p�A��kxQ���VC&,v��̌O=M��e�D��7O=(�1 a��h��#;`�Ls>�O�I�'���T�N�t�7m����vrf���V�l��\���Zh�2a�sw�q�m4N�d�V#��4�
K��Dwn&��Ʌ��6,�x2�#����
i
������x���ڼG�E�&S$���f�����m�������,z�H���n���F{-���yfŏ/f��������+v�3��������`�>~$]I��_^����R��=�E�y�0[�`/�L�R��oP@����H��U��	�ML�g�oط��o��6]qb���ԭ���V�ȃ#�;����|��|��%�5%(��%��f{,�W}[���Jo~�p��u ��pӒ���9�2,����Q�K�s�\�!� L.OgO���-�g�W��ߕ,¯���>�E^U�³�S�g2��0������io�*��q9^�N=m5���S�6 �$�\p��ϳ�����!<O���x��Y^���J��%��,�2�����8�_󋰜'�����6`���xB�W��܍=���9ɬՐKѕZ$��?M��I����o��k|��� ������qu��E����\h������
����P!hЩr�U��wƊ�P�u���a ��L�n7��ډ)��WQC��}�U\*Ww�ug�k�nN<�^~�����C�ٹP@IO���d�ظ��۟�����GX�!
ы��O�c]�q���sR�wy�E�'_=S;=����ΧΜ>cG��X�PxT�Gݳ�؉�ggg=�����^|�����184b,\����&$gΤ�T�;��ޥ�^��b:J�*޶��e<�DY�à3��f��Cal�Wфp
`b�H{�޽�����6�d���q��Ȳ����;�l7\�%}�h�.�i���Y!�G�3��:��ƫ��-�i1��RAf	��(r�/�c��K4����چ-�J�T�]N��H4���_��7�.�o|�i�F�-o�X������8�g�'��S\�̌ֈ�'z�YrV+�\x����ș)�8r�`7��s��i����.>�ģi������7�k
�zrQ�o]�+M����}������K�[�K�˚=��싞����`�`�O���T���ݘX<3��+/�>93;�=�<���#����(�i�p�Rv�``�_0�<Lۈk#��2��u�'�e��ݩd���k���j�z�<��ŷ����k�g��T8��R��%��i���Ǌ��hg���*���h�������Qw9m%�Aa���F>l;��O��0F:�:͊_���u�8A�?�ߙNI�4T���۸������I�q2.�CNf<�2v�CZ+Z�qj��pe<���U��w�8L[�G�3��>�+���>ʨ�I�)q}a���uЌ�=ְ�/�_��>������Ƨ?����zzg���b�iX}��X5��G�_̤&(�k_��{�����J�q�m	a�"�H�
&G����]�b)����7�t�%����?NV�U�H��"#ױ�A��+Tf�w���f{���3f�� '.F��kq��G,}�Ǩz���nzmǎ��p�;*��GE\A���m!d�� �O��25y{�8��þ�{�~���:t�.fb��~�j��ɟ�5�i`�/�!�!4 �I�z��S(�*����:��)�q聰įNT�����8�yo=7�cq���i�lj�D,�3����}i�����<��6&]��F�Q`���e���4�7�i�I�4�)|k�1���-}�H���t��b6hvv�勝�#���e�?n�ejv��p�A᪄�������3��#J?�\�2`I��a�+Ҝ�M�G��0y���I�0�i���.Ϝb��<G�;��^�������S��>8�}1�qi�,�"Xz��ޑ����ў�.��6�n�ߚ�nl�]_���|�o����i���vnܔ��ջ��={�s?�AZ�YJ����tH��ޫ�9E����E?�Ȩv�}nK����V��?�h�GҺ���+���E���4kl���}��ԫ����.-Lۇ��O�I(y�¬tĉ(�-â߰l}��S�m-{���J��W�Gt����W�G<��֟��E�:K�|�oݘHx«�)��o��-��e}^�=��\\�2]~V����̸�_�a1sb�2L�V��4m!���8a˼d�e�Tx���u8��+Nq��F��W���<����|�v߸���S_x�2�L_��\�S��E���7�I˧LO�_x忏�\���
y�G����vpͭb���+�g?��3V�Ȩ&�޲n��'�Z}���O��Kb��,�K�j\]R���d���c&���p�SO=�Q�G�/�8�*�)�2��g����Uz�����,DJ9�
���x
&�V3�G;��`)�Z��z���q|�G��\b��i��{�{�#��L���wX�����Oqd��l�$�YRq�<�H\���)���;f��a�7��~]u����9v���6��XC���0\�60ȥ��f���d����Ot��7���?ୣv��M�Y?� �ş������"��0^`{p��8���;��E��>�S�������������.%q�)g,��i�3@ܹ���L�5�qj&i�� X���'��`/��0�l��������J�°�K���&�=�����Xi�t�wR�o�Ɯ�#	�P�"����e��������ѡ��x�my��c��ȇǢ3��`?�	��c �����#��]��B^ͦc��,�"�-Nm���6FW�f��h��nO;�I����>�/5�W7�Uȧ�r���7Ӌ?F�n��o�5�^�#�p{	�{��`��bQ�w4��F��]�c����ƍ����}f���)�<n�,�xA���$p-����e�PP�m�U�D��\�/](��G���,�OU����eFE=~��o�x���3=�U���Cz����V'�h�}t��HYI��We0��U<�~��|���ǁ�`�2G�\�2l��F��tj����������imS��Ǵ�Aʰ�#�K�7�Ȟ�����;�7le�*Pq�𛮀�����-��ʴV������8���o��E��Y!�j锃X�"�,��6�ŀ�ƕ��'b�2l���|���1��w�:ՠK0��gո����p6����O~�������w.S@�pљ*cc>2&+��K�P���RGe��˕��BQ%O$�{OzC�SS �t����5k�,�������J�7mj���g/K�^}�5��4C�^���y3���g_A0��\	e�K���"�C�+�}��V��^
|�y՛�.�?��|��cG����=�L���0k��1�*�β`������DUJ8��g�"�s4���:�[�#�'�5* ��1�C=��.�+�m�!lA��_��t�6p�L�m<���oۃ�2�w'��4Hc�'N�M�6�����CN���S��-�w�?��5�r��q4�2���ȿK �6K��6K0���1��.,t.�]\�ЙE���a(��3�ݲ��t�*/,�D�-�	��?���a��b�cz$N|u_��`��r��\�������P�ᐓ�ł��8�yx�FC3���0��;���=�����)�9N���?T4︯����ii��̻�՗mN�b�ϯ_���gϧ7�ֶw�n*�^�+���3𒁢�Y��"X��y��
l�F�ў�����u��5�Wl���``�Dpu4[t�&��<m�?eE�G�h��7�J��f%6�ֽ�U
����]֏��ȿ	W����pS��h�����R�K�er�K���7��"�O��~�����@�2�ผ��ϰ'ڟ��ng���/ە���2������ě����c�N�0���Ʒĉ0ex�y���u@;��r+�+���3?*ٜ�g�uz�LW���)�y�_�>q+<�_�����s�+�����M{�=�~�V�[�b�]��@������O~�^d߸}�{9�
����{�c�^{�O�o���y��u�p�l+�@�����>F�w?��ӿ�'�'�!F����Tƙ�8�q7f��1�KK�ON�=�!?1�(���Q�<�># �*��������~q�U����R��u��豣+G�)�߬s`o�̍��{������?c���D/���V���غ�����':p�K�~�e�ы�����ß����P�֢e�Q�Tq�c�+���G=�W���_�+���?�>��Ÿ��0���i�a��#>㊫T���SN��q�<O4}�I_#�q�.i�Y!�Ù��  @ IDATҴ�hxx�� ��0یp�&���S�#-�������L�8L7�|M@��E¦M�J|�8�#g�4��^�n|M�
��q�G��^�'�|:n	�.�P�,��I��'m�4�h�X:|4o����<�BB�J11m��η���Q�<�ؘu\�"$R�A��&�M1�67;�^��+z1�\���K����5Ȓ�Sg�g8��ǲ��.���p-.�&_=c����w���wo>��1��12w��M7q_�o��k�����w��;���z�~����lf��G�7�׌�w�q�p�#�ٷ:q���������n�]����9e{A_xN�����3S��V�Zپ�)��Mi�D��:�U*ٶ���7�h^���#�u���z���a�����d:�#LzP���p�Tؘ���餭��J���TW1ԝ��M���4�o�@�FbT��x�J�w����,o+s䐑�1�[���d��w��o�r��L��n\�g������/ay��sye~G�.��驹ʰ���Ϝ���_�^F?G,�r��^'�\~�a�-����R�g��jc<i@�*����!��>�4;�R�����?EF��Uߪ��8�j\]xerA�Ȏ�N������=���/�4�P^*B*/*4�U]����m��G���ꭷ�*&0����Q�+�X��h��T>yWaą �[Euǎ���q��g�N���04��]]��>���L�o�=Ͷ������t�cL�\�i���y��]{�ˈJKgM�Wu6%O[���0�7(ϋ�|Y��S�� �'�w�;p🾽��O�19c�*��Zy!��I��;�u���.���͕�}�1��[s'�7~aP��S�@Zǭ�Ʊ35\�J_z�p�}T�.�T�4^����;:)�hp	"]�7چ��"-i�t�Zxi�^��q����m���=��mjo�rYi"c:�(�=��{쩔i�Ǵ	c�̣y#��N
��.�5o���%�%g̼ck!p���t+��bd^�P��J~W�ҵL�+OI{I�a�B�1��6��Q~�F�]�&��?aXj(�!;�e;s�t��4��L�,e�f�3�X:8�Z�#�GF�$~��3'9-�Y���tb��Ǐ���f4rD�@��%.���c𯹖;�&�(��,N��mtm��5cEb��7~��<v��̆n����Ĺ��q�X]0+�Ǖ�i��q�Rs������^��{]���uŦ�vM����K��`�{��t���>��?c���1��=`y.1z��N�g��\&3��O�VW��Q��[7t��wٖÿ�m�o�,S��Q�7x�>���_�W�m]�<�;h�.�������}��ǺN{�<FXI�$����4E����2�9\}�N�:~�-]��[9ﾍ'|���EX��x�i	Ե4�n�:h��L?�c��N���L?��'���9����9�a�wU6+�բw>�����&b�5���LSn�w0��i��
�P,���Gy$qH�򯅜l0�5}�]w��я~��Y��K⊆s�w�y�W�X������Q�6�d�z������{�CB��JN6�T��c
;!���8��T�ByC�t�8�l�K�J%Q\~� �T�֭]��o��q�k������:��z�:wYu�AS��q�
_��/�����G1����_��q�E��s��T�u��On�a<�N��ri$y�!�[�>��C�~l�ː0L��Oj6�X&G~#�eyG')�t��&�����X�uO>
[����~���r\�z&�&���X��]��W���m�A�0�&�tI�va����]��7~�6.�	E̽Zcc�#�M���6?2cu:�+z(����Q��T��}��c'hct�.l/�X�:�P^�Fq���̠�H׼�W�4��(]�m\�_**9�wF~��ҩ;��Oi������x{�vc��+�S���L9�?��I�Xy�H����93�>39����e�K�6�)8Tgxt��a�bv�;9��ł�շoJ�ӗ��J�>w,�?�>�Ѵih}�vj��⫏?������;oK�|1�bY� �2�1�.g�<�-��Y���bc�[o����{>�f�����<� |�l����Ò�Y8�_Җ��W���~��Zn������8�_�䯌�::����_ep��^����W߲tn�3��6�k��F�+q֕��vv�o���mzm��Y�rz�β����~2n�%_t�x�LW�%����6]����r4�ηi��0��H������'�.���xex�����U�����]�����^Vn�[��`뻏�K����hX)��ٿ���4���'������w�1k�@�e��O���7�a����z�W�/(d��J�jb.H�p�&.���W����t�1r���Q�(�T�|+d��n#
H��+�WARبd��@�_A��rt>R����-���]�w��̥�ɋsk'�ņO����m���������-�ܲ�4���\���+$��h"����ݻ�|���!��o�oy����,��<�������c�&����G�����(kyN��QAv��E,/�.��覃��E��3�_y�;��w(��g]5�8��`��.�'���=^���`��mE<������2ی���t�Y
C%J�1���p��;am�]f&ޅ�ᬗ3[�K��30̻�=z]>��T�:����{���X�5��*Ө�"�Z0�5'\��ԿEU����7y����?�ɿ��F�-c�ͫ|���e�5�6/�#��W��K��\�͵�c�cI���M0K7�R�%�
��bHqQ�,���|Nα�k��1vfOO%�|S��`��ay J��usl�:�ٷk��4�v�	�����v����XVx��������[�Si�s?O�7ne�l,�6�����w��4O��y����J*IU�*	��,�%��1c�=M;<v�D{�3�h��1a��?�c�c�c�1���������<$@�0`	B�G��T��wfe������u�>u2U��*�:y��{��^{���گ3����>}�8�s��X.����Z���N/��������ʫ�x�7���Յ���O���eF�ߠ�na n#�W����r�hC��X���޺�2�Ao�z��}�ш�Q��oܛ�3�*���Ό#ښi)>�]��q���p»|0(�_ ��΃��
<�ʹ�g���S�(�q�	�̳&d��}Mr���o~��+��Kת|kC�<'�N|��V��擶!��.�i拇5��A?˰�|��ȓ��\�*�����ț��aDy��7u��Y;��$-^��m�g�h������֭[[�O�l|�oY}��k�}�^S*M!�?�X��Ջe�s	h�� ��'?��{8Ŧ���'��4T�*�\��)��np�-2�-�Ə�O����[�`�(��IE�2U�9r���������_���#�gb���&��Ea�(��iT�Y�*�������PN�Y}d�m`���dk6�1prG�q!��8�]YQG A@��38��I��Q��O�>zρ��Ʊ�J;
'ub��8��U�4ːl��/o��ު�&�<ڟmM�_�l��Q�zIJj����#�y��'�4rv�2��%�t�0�����gnx����_��K��g�|�|7,��NO8d�wEg�ߞʩ1���Qn�]�7�c����Y6qa�̱ΨK3o�s��C8����G�[�8�B~p�b������4>f�p��!Q������!?K	�YҡK�YJ�v,O�Uz�!3��g�n=k�ܕO�KU�.;d�d�,x�p��,�S/��ボ�_}ܙe̻�Q�ANTdy���)N\���/�Y���lWɖұ>�M����)��3.߃v1�^a����Wm*F�{�;���_�F���_+6-�(�m�-�o�������āog_8Zlٽ��>�m��){lQ��L����<��Po�`f�g�����#cퟦM������(u�ʚ���a�z��z{7� ߈n��vm���e;��h5��@͵�j#�x����UF��f#�A����5H���6����`z�}��ک2�Γa���|�?9D���z�>��/��Z�2!��7�x̘d��7��;�WyD�ÏX��P�ɰQfqH�K�ґ��#�.������r���a��ӻ��Kxk�����I^j�3_9�|\9����.rϰ����'�h��4��_�n�i��❈��«����1�v`LǊ���ow8u�`UP]�� Z���9����z��	]M��ϯi	�;W���ym0ǋ߃�����9�bH倁f�	%��c�##,~s*�:�f�p%#�e8���L��T���qxT�˦��o("�nʿ~��b����߷�������?�x���J#Vx��c� Okž�,Ͼ��w=v�ͷ<�r@���,����z#�?���9�:P��۩TM���1D]q��o#�Kf��R�����ՁC�v��Ow��t;3s�-.f ����ј��cѥ�W"�9n���+���'��p�5�3˜�����(�;8_t�20@'h��,�Y�=��@8��2�w��È�PЈ�^t�.I��ԅN��j�Ʃ���nܴ��
����9���euy�Ec}n�Y*�f��̰h{��w��Lzž-`|E�mۮ�r�a�xVC��a�,q&O���k|�u��|���;���̤�C�08��7��A1 *ܛ�E?'#�����!j�)�g������O+g��#�N+�Y� ���A�#徯ʡԩC�!3�5�s;���S^���u�e�iM�<�Tj�8��b�p��e~���i;N���N-��Y����[Y��T8K�r.R�9f���4���k�@p����R��_��/{���ɣ�pg�����}�e��JNW�/O����n1z�P�w�[�}i��35]>��,No*F7�Y�n��X:�Sl�\�!ⅅ�bj��|Ը5���后�զ�Gx�߄��/)��;�U[����齼zai�O�:��CG_=�{���Y�]TF6�U��N��X)����;d}�K������u��=�6��������4`��ژ��kX|W�h���1����Q�_�&}��ep�P���.����}�W*C�ƫ�[�@B._�d�|ޑ]�l�df�V4����M�F��7;zƭ�o� �l�	K�,�8}��1P��ӠU� ���C��i��_U��sz��<�7�G�&��YZ�,��y�efi���D3]}�����
�d�L�{V]���q�����b���o���R�����o����C�T���^*Xw�.���	�dD���q���/��j�by�#2{��o�h`a�Ǿ(God]���u�+N#�c�HVL�Sk$��c�=�癧��8p�T��"U��ǈ�
�|ѡ���^ܵk׷9z��3���.���]��G�{Q�*w��e�=r	���3���AF"�Kb&�m#;iww:|��N�<����Y^f*c���M�0��+'�6�\4��B5�RJ����Vp�-p9����������Rt��5Ф���}j�KӶ�,Qrb��u8_1�j�t<����	'LXۼA<���g�� <��|������'�9;�;"��:�������+gK�\1��n���C�1���:�d�g��C\���?�=���h�a�;�TKP�_��@q��Ј���h䑗����u,�*#3�]e���+τG~��γ^�)�at���<�M����D]?%r�
ߢ�q�+�S��i�P������p�K|�߃;z<���غiF43v�
N�,fq�Ƕl+F�Su�����7������S���a�r{9Z^�a�N��>���9f�n��]ņ��S�)�����;T���k&�;1��Y��^u�K�F)�[z�zo޲i��<��^�Yh�Z���-,����o`�m��4N��t���+2�!�s6|�����v�*�U)c
���;B,|~��/S�yx���h�׿I�ϑ�vx���@������ ,�Jo�|����~~�~�}!�|�6d��.���X��>��;�d��4����{g�]jfϴj~r�/�y�M���5R�t���U�'.�t�8̿�w�,��?5����̓�s���ix����Y�s�X~�s��[�����Q���x̰˓��U[)�`�Ow��]�û��)?����=�����9�Y��d�����y]��֝�K��~�n����ԧ>�vN��0b�R_�EF_4dP&�(0�b�K��8WaȨ�T:*V�*�vh@bɎ��B�4J8�8�^�:1�dh��B@�5F5��w҇'�k�5��� ���$�-x�VU��/�?�#e�C�F,����ܻ�F.�&�T���w1������k]�NGhg����#8X�-,-��N���ǹ`��2ő��ێlv��6��m��|���d�)�,zt�����]y8C�\�C㐥m�� ��U΃q�Q���.�������+����6j�b�k���2n���ɏ�i��v�3����N?{��%�]�} o�qG9���qm�[K�欰3�����I`c6��ȣw�	����Sc��:��x�e0ą3I�������(�Ue��,�i\�~-sC&�K��!���p浾�cP~qW���/��.Ʉא��(7��l�!ڋ���J��y7XFh�s�+[��a�&��'��0/�/�!��`Vl#ǹ�C���������q2j_qlq�<w����+�F6wl+��~�k_-�_qE����(��V��9_�����8��
=����i���c�l�����mڲ�����oS�����`�U�C���L�ţG߷���ݬ&���l�����Em�&6C7��eZ�⅏t�A����L���m S���=�����V�����5>�7a�t|&��5/�x6��xx���v$.�_�0���}?�h[L�iЏ����E��4sM_y�N��~�_;9�+|~W����󞈲�-���	>�=��|��AO��U�_>R/����k������S�7a��4�����/���,�c����1tF�a�(b�]}�~Q�;��q�J�\�=����E��X��O��	f����5����EyY�������~���P�8J�������;P
-1��8T4Y�.=i���#�%N�RQ		����Ѧҏu�6�[6���~��}[Q6�q"{�·1hdRV��Tn��(��
%v����t������4�P�WD&�[;+|���ڎ���PǨ�����p�1~�����l�M��P�8n�|@�>9� ��	�����}j�fة�]Z��ц�\�E�-��/DG��xm��SNq��`�;���G6�cv&��;m59�q���;�bE����;bGk���	y��	�tz\�����L:	3�8@�B�_��w��Z��dv#�IS<�²��>��v�	�,��;��������}_)vvccv�^8tByA;�k@谑/�֔���(��0�M��|[&/ಁX˙b��2-�e���X^�[����Q�2��2�`h�k�!�g��u���
GW��#�h�\�Qg�<��Zx���O���$��w��܋y�����c��gW�)��3�&��\w��Bymw���v�its�t���/<X��7��3x#���Sg�b�v����b������^;������01{}���H�����:抾��w�<s�/|���c�z��0�cH׮]Ľ�W���&��f|#�;�I���W�O�gm�7p�y$<�`�y��E�D��D{d�����C�\�å�7�	��4�\�'>������\�v��pd��4S����	A�w�|�ǐh�X�'=ޑ�C�?�p��aWͯ����h|���m���%l�#��S��i9!�����:滉�	���:Ʋȷw/B���Fz�;p�C���W�$]��L�b J=��a �˲^�����|�EW��=��������Ol�xb�кЈ����KE��եRS�2���=z��1z��?��=�d3�R����T1��eP���.߼*U.��P�(Q��Ai k�"҈�o�hX�N����tx�{�{����U�����;��1r��8e�>��~����{�ٯK����kֺy衇��{��� �V�ة�����X;fڙ���vI�kVi[>�k����R�_d/ѭ����'�g;m3.��<v�6DQ-'�嵍��8DF3q�	��dU�*C\��g{��F| ��mMZ4�z��p,4�u0�m�5?�7��{�����,�1�<�do�֙�D)g���#=�7���XJ����ɇ�uDp.�1�ՄӖ��h/�ȏ�c��-���!���cvJ^}�;���2�K|�]���Q��|,q�U�/�m��]ݢ��W)�L���Ǭ�e&��j��x�
�̤�<�2'�=��2
'<�*;���6`~�O�Lsugf�E� �v����#^A~g���c�X8�r�Q��-��u�X.zÙ�>x^Μ)7�+6�0�ž�g��d�Ԇm�Pk��z��_���2[�㯝[>;03w����M��!�_{r��U��CF�G���B�3ȣZ���
ߡ�{�w�����_<}��M����2��'�/gSD�Sױ�ĺ΁�k��%�p�
�V�a��ͪ�x ��AcP��Ui�t�|���h����fS��v���ѐ�
u.�����|od��We����N|]��,I������=�!�tn�(>��2�82}�L�=�f��=蒞��hH��NGMc-d��5H".�6i��|_��E?_D_�F9�eMk妮�ʷ<>�ob�\��u�i�t��2u�K��1�t����+�is�z�+_�J��[���{�~�	��O@��f�h�^^/�_>�z��.�i�66Y���?�����ia��(���١r�Ν]f�4�ÀIJ'�����tH���v�z�PA�#�,bm���,�v984�btZ�rS��Û�h*��9���Z<��֗i-�N���Cu�l�(��COc/|�#��a�� �|{��|/����V���T�qJ��:�"�¶�m�N,;����ve�ݲǾ�����"Ѽ�Ly�0���0�C����*��p���Y��F��϶]�i�_��rzj��� t�}e��� �N��b����g8f}��N��kA�{�c��`��q`���g���RgS�IG��<��IWYH�w��O:y�`/��9p����h���c�.� p�P$�����p�B6�a�E[�ҰDv���wZZ�өQ���a��	o>�1��|ZO&�-�[yG����:��P��4K8�ֿ��ݪ%-��_ԫN�����і��)g썳���p���U�̕�*���0h9T�,�z[řeN_�0�>�h���v1>��Xj�|s�t��w�<z�`����U��o��{�m.��R���/��-�����<����.U��Z`�oie�lc��"C�xlrr�� �I==>2�u�߹h�?�?CsKK7�?7�~��v��lWփ�_&���U��fc?��x��K��hG��3҄M�k<��?�'m"�|���e�Pd��<ⴝ&�&�#A#d���h5�a�4��v������啟�G��o�����J��/q�t��3�tyn:;Q�O�/���o�3}������#x�n3��Z�i�����)˦Γ����o�q��e�k�W���:O�_ÐW��
5� *q�<��s�<)@��2H�����;�n�>B]k�:�;�(�y'�348R�9��%�����k��������9V ��?
�Yx{��X���ږ��s�ڮ��w(���	f�����p�e��ii԰�����-�H��7�Y�۷/�ˈ�Lgc�Q_c<�l�FA��4�N��#�K:�B��#��"��XUy	�S��<�b��Xӯ������T�9/�����a�(V�2PV����YN*xB�}h���n���b��Z���p����%^��87s�}S}1���6ӠK�~��n�2��(;B�Pϐ��$��3R� �������`�լ����ְ��i|��m���D'�A�y��y�����"���f�^�p���gfll<��T�c�3�����r�eo��i������ߤ��߷Q�7������Ӫ���G.�r���ӕ��5�2ʟm+�x��e�7��K�$g*�� ����	gVғ,8���t-�<�Oǒ|��<{Y>��%�c���8t u�|�a�B^1�i�q�h��y�a�*8ʩ����?���;��\rbE13�ǟ9�s�ؼe3�p8�g��H3AώӲ�5�gg1�s��V�g/{��Ly�z�_���mW���o+F�(�mst>ۭ�C���"�=)Ƞ�f/���}~����F�߇s�,2q��7ʔ=�1���8s��<�֩��]��[���z�N��K�����ڱ�^a�Z��NW�S�!]��j�)_��Hy04��7.����k�H�`���gpF���ot�7�&?�=�����˕x�����/��2ω��MD�w�^�'��L*F�N�=N������=��&�Ԏ�l�/_�g��.�L'����+���L��>iu|�{�M�kC~mZ�w�y�����F�)u!�p��3�Q����#�!�b/a�Q��#cG��v���i�1��
�Z��S�$�~���ҟx��+�7����H`ݹzu�|�QD)\�!oaY�v�Q(Gf���;w�2aF�����Jƀ�f�6ѳ	E%�񦁧��"�%<5*Z���~�A�QX�d���dG�3$Ew�Uz�\�̜��;��G���?�!
���C9����:�Ύ(;e��;�,�P��8,Z�W��W-K��*���ǹ��(��8�1j�ņM�d�U�ڙi02�=zٶ��r`qp}�(��t;@�6=�vu����mՠ������#�L��t�!`��t����h�z��!:v�	�2�%6<�[�(��D��#����yX�F�K8s=:W��0zx��+~y� g:���m�,�N�0�M��阹�Й�j�!F*G�+/qVE	�(^��M�?�[/��qŲB��-}e��jp�o�޹j�7㕆��
�6�|�ūS��̓u
��8��@y�pⲎ��Y-�Uw)��c��d�q�ٻ�a����T�<u�;�L��F>�܃��[�f���Sr�E��-�f������E��+���C�8σ���fŮ];�;�n+�N+����ɽ;��=7CǊ���C�����)��!���9?{�S7m�������	d��اᑐoD��БCơ�Bq0��+f�|F�Ѷ�}���؀��Y��x	�}�P��ty0_#.~ۆr;2-�c���4����'�{�ݤ{�X��%x�z�ۄ���9$\�d�qq�w�|9��ײ�w#O]�WϺ$ZU�����Ȍ;�x�~����ͼe��c*_-�L_ؚhz�<'���	��_���Rikq���@Q=�_�I��o[��兿��,g�c��M<A�>Y��1�*��NV�x��:���x��'�����;�s�Y�/�O���֫~�g����WP,�W�:�KW(g��ùzϧ?��(���N��0��r3�����	Q�����u�0�b/��(�:?:aѱ`�x'K���ӐR!���&F���JˎAx4ȸ����o��3����ߏøx-U�(�}���X��БS��a�����U��P��(��~-�^ൗ���Q��R�wS����DI��0"�'�c�X>(<������eGm;���̨2�aIN��]�\��H��0(G;Nq �hs�Z�&��'X��KGOXx�v(/���lh��p���qP���[tԱ�?������k~����!�/��J�,g��9���B��XW8�{{b)�NPr���ҙ2���9ީ%���[6���8��G�����oi�q����0�����N�J�[�	r�k�UF\����c���,lo\�
g{��B�2���ٺ3L��֭�	\1<G}�`JO������W�7�+�,g��-�Η�NX,g�~�o����Fu���s���3��qxFp��;˧%p��Y����Z����ku)a��G]ai�m��v�����[���q>V<����({���ǋ+{��6�/x���W'��Xw��˂;�8��&����Q̾0�������۷�����x1>���h�;z����>���;:|5�$�z��wL9Z�1;�8��:劗���N'�6L�K��x���x���J�e�*�\U .�.����&�ܨF�vHR��?�ٸ�]��,�"����HE��"�yl;A|�y!dؠϏ��_�y�W�9?�Od�$��~���V�$��ij��9�d�����ϻ�����\Q߾^b>�K|�9�]����nO��qE+���+`��1-�6ΐ�U�Ry�є�iW�K'�)2�zR��2W-�x �A'޻��~l���-��o�[q���|��{�5��a`蠖t=����+m��j�����M [�sYH����,��^�W@~0��<���Bg�#����
fb1�M(*SV0n�t�C+F�5��P0a�p4�PD*Vqw?���Ѽ.�洘&�b���*3a�Xc���)�1�2S�-2j�F�>q뭷^���Q����W|�)���;�U����r�ZDnm.7Ӟf�I�{��B�=o��.��a�^�1C�Y�\��� �qiۀe�|��ώ�6�E�m>�Q&9���8�u8�و��`�/�ԉGǝ��jy��4M��l[�2^�k}x�Sg�j�Y����]�_�r���T�%�"y�cv��wqo���Q|�N����ås��w�&�!�Gg`p�ʾa�}��py[_�/�!�F~x��K�~,�>ei9��A�}.�2�Ij{adJ#�"����EYɻ�/��@��(�Ύu��m9uti����L�:�g�!���c'}/��޴�����/�Tw�oL'�٬���3�1�X~�;��"��g�g�s|�ydh�����^|^�qrj|�w	���,1 ������o��R'8d�nF98��*���)M3�v�dw`�,�n��ޙ/��cŉ�W�C,�k�(ϱ��3W�x�^F<�>??��/'�s��+�ѿ/P�Wj����n���M�������>���ܣ�k�����6��Q��n�B�)>�0�צ�f���w�7�yO<������x/��6H�v�Ѷ��{�%�%��m\*�p�M�W�mઝ9���u���8����~7e��e���E�S�:^��c<���s]~ְ"6�asޚ�k��\�'��g���w��i��;�F�K��q���;��3���,�(�:A�������������Qoi�wJ�M�#�]�]w�I����������|.��|z3/Q���KT���%Zq?�Q�0o��[?�O8�4�h=������)]?LG���Aa�r3��F��E��q���#�F^��%Pg�:���/����?�a�T�bd鈴JL|�*:�
GK#�ߡ���ze;��|�O�m����e�0�7������7!�Q�0P�3 ��$T�<��#��2���0Z���k&�[e�H��n�������=f��v��F{X�t��Ŏe��j۩i �f�g�!�i$�/�r^y�KA𜍱��;`����Cg�u�haa6 W8z:�gx���ˠ����q���1^y�}�*C��}���x�O��t޳���怆��W�'����;9>���AS8y��1�Fе<�#ߐ�e�|1#�D����,Q>�c\�I��*�)k�˓���4��f^>�7��U|5���;�#PyNGJ9K�Y'󫃒����r@u�����NK���:c�#�E������^�sh�"��C�Ϋv#����ɳ|���=�_p��J�V|�dy��0�i|�j����cVێb�E߁�r��dq3�c����������X�y�[n+�7���8VsS,7�g_���2���Y\X���\l붛i�$���uő�����{)����l�13&Ѹs�ǝH�	�]��5C���m�8����n���I�Mn5��'��,/y�)	_�M3^�>C�i�0�#h��j ���/_�3d\�9��O�8s9�o���LӤ�E��f�i9��l����~��G�ڡ�p"�9�(+ޭx&n��3�t�(�&��k�J�ȳ���|�y9/���[�?�I�;`,o
ᜫO��X�O��_=��5�tY^�a_W��^rP�`+��D�,��f�?X��)�xz�z��$��\]f���Q�]� ��8Vw0u�f��{�]w�.���׾ǭ�\B��x�CD��13Q7)�*!�"JHcl�<��4E�2x�92��l���������@:�X�[�JPe&>�"�-�P=��Os��9~���?�,^�y����|�;�Y�Iч|��
_�C�k��'��p}y�������m��f~�2�C\���A�l�� Ù��b�b����[���߻F�r�2(�F8���R�)�̗�jL8������xw
�Y����t�ü�����4;W�-�/F�h��h��f���8O*�}�T�
��-'���܃�ȏ��΃tuV��2�.�)	���x��#��eNMd�P��8���	�G^䣑��Y�\2 ����XV�Eeb𝴍�p���LW��Y~@��7�!7�����?���+S��ı,9��e��x��:Q:�.O|�K�:V>�ot�p�4]��@Y&��ᘙOyR1��s�N���`��h^�^���Och��}�٩c�,���r��^,l�����s��rpt��7���6���w���x��q|���zz[1X�~��Ȗݞ-嶝{�e��4��S�J��/��;s���������]�&�����g/1"�V�2�9�ό�oSV��J��Y�%qQw �O�6�4ͼ<�/��"-���]UmȨ:O���x�|�H�k~7!�Z�Ӽ)M�*N$o�3p�}�C�2L���!��ݼ�&�V����<��6���3h�̉��Oܪ��qE��e"�:�w4Ӕ�Sy�̺2�(���i��8�H�*9|	�u���Ei�oo�/���)o��3��VF�8/��W�E=���/+���˕�`!���U�~���t���X�#!�#����2�@m�\f�Z/�!��Z�d�.���/}�K�7�|s�R����}�Q�E���ALq�`�0x�è%ut�q��F:�:���}������_���޹s������;t�D?�	���3e�s��>*���_��_��(*��W�d?D�/)P�D](��N���rF��E� �0����4�V����6�^IA�����yy�ۯR�]vB��sϋ#}���al�e�/pZ�崓�(����_�#��9u��l��%�6e���P�-�S�<�w|�HC<�������:g�쀽t��w���0��'O��y�/�C�S��S-e$>hZ�,f���Y���l����f���Y�K�y���o��_�cĵ�O�U3��2��,��Ŝ��N4=;oy��c6�x�j�e���z�}������ �������^�I��,KqqB#�����ёgۇu묺8\���u���Sg�4g��A=u� E��o��q�_���򔶿��.���(�JL_W��A����Ǐrؑ��a}��Gퟣ~��ef�8�ժre�&�L���'���篿�8��A)��'��N�����j�����-���l�vu�(��2(c-�Gs��7�oڸ�������}�Z'�O�C��=���n��Q���b%�J� �0p�e�o~d�9����n�(�0���m���~�#�|<��6R�ֽm�v�.'�bvʶc0��v���ChD�0)�%�bs���U�H��-�y�	�k��2�dЄ��F֪M��/�ȸ2�����K�Ο5,���_�R��=�cUB�#���&Ȫ��S����tz�y������4y4"��u�#��AY�9���/y4�K���`O�Ew�2{��?��˙���2��n��s�����w��8��������suy��[�^����^s�F�  @ IDAT�����l�lqꞣ�-���v��kP�X4^T*�Vi4j��X��2R
g�$��Q<�`�|������w�ڵ�ٱ���a�j�Q�0ؤag(����(}K%��0�H?�r��9���|t��[�KYb�đ��e�-:"��q$C�u������K�e�'����۷�,���o��>�j�:ce�a�3���#��6e��<љY>�iB�vZvat*4�5���#�Qh&8����z�@Tէf���/n��o�Ƹ����b��4u��Y�z�B8�u�3����Ge��:��x�2My�F�q8N��,��X����0K<�� n�
�/�a�A�
ǲ2�U���Hʯ�2�7~Ǟ-��FY�P;'��'�$�,�#�f��0f�.niX�LS�ɳK�����x�-r��4�&g+�ۮ�<*SC*[��h2,��f�O���F�K|v��Q���D7�8_<u��8S�bn��w'�7�m�|�!��ё��%������lq���,�p,�8���7����S'^(Ϗ��3�8s��;6R�|�v�v����ǻ���;6l/6�O�--��u�8d���a�����r��ƻ����C��$ŬY����l.�ۋ�~'��\h8[u�`���hFo�F��&=W	)�[�.�r�=������M��	��3�f\�o[J4y�+�ߙ���)+-ۚϤ7�v��2����$9��3`���JL��l����oZ��������{�4�?]!����%.�M�p�Ƹo�Pä<A;���K�euQ;~9~^���Eң�k:k5���<ֽA��CŠ���wθ�ws;A��xu��ɖ��ˌ]탾v&��R�[���7��Ļ����ك�9�ϓ�xMt沯�_Y	�;W��</Ul00~��y�aYMg���(�6p�0+8��I:�X��F�;��z��OI{c�?��{��ǎ�گ����ڀ��f����GiEq��T^�8I�NNG~G�=�ͥOg1�e��8h�8�?�q)V���p���?~��ij�(�z����3��1���Z�,��� �U���vu���G�V�s#E��V��1{k(c�����it~�"�sˬ3@�=L:�)amc|�7��lt��QN�Tx��l��7z[����z�+.�y�����8Gv�R��us��w��{��i�͛߻y\"������\�_9]ՠ���U���G��$8c�[��(��n�f5ډ��)��������$�G�˯��k�S~>[`�83^�#N�=kf0o��2չ���N%|����������ƌ��=�/�[��oq@��r��������4�W*���.O�]�T���@�Y������=zG�����5
�,�&t�P��Q���|���f��G���<��u�����ݻ�g=_��0{$�Ttq3�����N�+��bj����NF�G��YB���戂{��s�s#�x'z�)ڤ�aC?x�b��C����!��h�uD����!�
���#�{��*g`�a[�浾�k^�G>�<�p|�OM��5�&N�R+���:iA�6څk^�'>7q�N|e\_ �2�y�~3==�<����暐��=�a��HK�^/�Y��U>�2�[�;ш������nu�F{�8l�?��7馴���H�������-O��;�m��|6N��������LSO��l+�&�lɞ�8p����>��q�%�Ӟؾ�{>��N���+y�u��2��J�Tpt�;1~ggF����[JqƦơ�Ļ
��;/�k�cl��`�{,��ux�
�Q��C���ۿ=�Q�(��%fĦ?��O��:,�B�f����F�F�J;��=ǒ�Gv�������)㻌�}�o���?�FLd�V�vH�<{���s�޺;w�\d��kEF8U�������c�6��`[���=1�u.�����燓,b߃e����Ųp��)$ۍm�6���Rv*�Cf⑶t�Ѡ7ov"h_A���Iu�9�=�7�wg��3e�#&����qѐ���O�<͖��0��Y����/-!`�9���sy���"o����'́;x;t��l�{��U%/��D��>�QY�SNމ�6$�lħ�i��ˋ�����ډ&�ɓ��4�Uf�sy�u�㳲�~�rX?�(/�J��S'˲�l��cۑW��|�߲�Ol6������t��6h:�5�P*[G�}ߞy�b��qf>�X8{~��>7U�m�r���Nw���I����</�8��3��mӝ�����[*gN�,�٣����57�T����)�>p�hw��3���.�����ũg/lz���G�2�3ʲT�a*wG�-c_���_8|��ݻ�ʱf�	R�(��p�>���+�T�Ң� �������ڋ��P_5\~�s����AѦ�+��<�{�[�nj�!'�m�-�f .
��I�H'���Xf��F�.r>Ң��{�P������ኸ\�&�r|����Y�#�n--���)�S󶖗�;�g�^�~�I^����:j��\�L�e���Naԁ�dmy	�>|���?�ꨔu���ݐ?��O-����.6N�X=���������g��:�	h\�o)��{Xw�^�- e���(���A�С��Lb�0�oa�sUqdCU���Q�$���e9*h��E`�����F�`��_��_Q��m�͝|Do���S)y����p��#<>!m���������;w����!l���W��.�D䰨,��� u�b�Y?I�i���n�	I
~��z_x���>���9}��n��44s>+���������):*�--u)�,&�i4�_���d�����f��5�����D`;�/�4b� �q��A��.��~97S�;<2��{���WZ��!٥u@�Y�e� �����I�#^(6o���<j�ܹ9f;8�z9M�~�>��<�}�|��D�a����o������D8R��N�$�w���p ��䜭��@>v�w�,�0�f��X��~q��I[�QҷMGzK�Z�*K����-ۣ�tjL�N�� �p�Ο8�3�}��d��I�����iֳxL�8�cGyӱ�iȿytL��r�
���]�;e�%g�p�ĩ����A��W�>�q�������9 �=��A>\�$s�6������夜!+g4�}%{���>>A�3|<XyN���I-6��K���,��h�gv�h�2�.��bS�����f��c{�-W�P��>�������)��?�wl)�o��8�X����Qʳ27ρ��Y�=�s��쭩c��l��ౄ�^��؃�}���\m��;�ne��H��y)D�`]����"WA<�:My�Nx����3g����=г�j`�>�C��}�A�E�[Ue�6�k�)3>�L;���u�p����n���{ɳe5�2�A;b_�O.� ��������@Y�>K+�5��n >ޛ�]8��o@��T����T��˙i6�Ur��7䓓ވ�OyKx����B����g9o�m��|&=4��w�p�3���&<�b�C,�vG����f='n�F� ]@����:R%+s
O��W�K����w}�=���|_�,�V�6#]�_�Xw�.�j���Bɨ��Q����=���* >B�2�Xo��RɊ��P��raw�w1d��	:�{?F�߱��qFq�~�#Y� q�{�C=4�㴙���1�̊_�	���
R��������~��o��;��y�(*�h|K���v&��#�퀬��`�����H�ߎa��K̂<�OR���9�������ܽ�a�s�s��1c��s�t<y��Y�Q�^=��(a2�k�BB'��k;U&�E.��P�a����Wpx\^��f(6����ƺ����N��~�eaSS�2F����<���{��R.>���>:U?��a��!��A5��rH�h�r�lT|[IZ���ٺ�a�L�P�_��%���쌖�S^:r�c՞,�\�e���f�&H��@1b��g�R�
��0<r]d��4�K�s��/�e�Y�P&�u+�u���0<�����#]��3d}���|���ũ�'-d��n۶�>0ڡwtH�3�7���m~B��f�!�V�Os��aЙ�o?&;J���TmA�8U���ㄵ��eӃ8X�T�I������.S�x�:_�|D�C+v\ueqf��bKxKO������b�������/VhW���<Ns�[��ʅ�r	���ԙg�'���骵�
�%����@{r9�/�Џ(c��Ƌz��(G*"��%PEt�5 �͕�|����Q�2"*�<�8�Rw�ƣm��_ᬇ:�4��T5[�?dY"�mҊ����x�q7-��&oh�ED�'�5ߍ��G�|��h���`�Z��nN���&>~�r��I������S��4Lk�o�֏kaS�L7�!�W�*��|����ɧW3� ^��HK|\�?��/�����>�d��4y��ɇ���=V���N��A�����4{���w��O��C\��Y5�fA֟/K	d��,�z�^V�t�{XR�8:��߿߽��4�*��Xo���`�����Bz^>3O� �F��%z����5���O�D%Z7|r���%��u%�T|���G�C��4�0l;z�V��sj׃��IN3<�U�k"�كegyA�g>�a���4:�Y�v�At�֙�g�S Mc�y��O��zR�O$�k/��W:t�_�<������Xk��/�یl_������0�??=�a+�:��r�&��g��N�Z�:�	r�ͻ�t�lS��6k��cƖ��kz�1�o��<�.���5���,Q;�F*�+��~f�Cy*�|�����,�A�F��o�2��g�7��\�kyp��a�\:��脰JT����<�̮)a�k9tֈ�r�<����8�q��&��)4#|��t�Y�-�N��%.��T��,�vJ����̑��ѣ=D=�N��B�oy"���4N��jy��O'�M�赨wdG$��������XR�L�ϱgϥ��O���]F(^�m��3�[Nq�`��Ϥ+�P��fe�ռ~U��s|d������v�������7�S����r�����8j�ņM�oB�~�ݣC���-��Ե�s}��0��閬V,V�?u�L���aF���(���H�����w�ǽ�Z��m�s�ZV�e�q���D����1.e�|6�����B�9p�<5��=��I9Og}y�>�}�vm������~�ɝ��.�-R��e����|�G>���٤�	q�e�mW޲L|θ�4�cH��>��,�!Y|�o�'>���L�Q&\���̓��r�,|R;S9=ߛy�̃��9ݳ|�y�W����;�Z��`�u�#ѕ�o�m��?������?�$��C+��X�w�|��ԓ���8�mg�د��;=�B}�a���������?��saD*8\�s9K`ݹ��k�"eC���Ӊ�<���=��#��]���?�Tѹ.���o�0�TlQ*�ހq�.bl�{�?����{��E���ph�����mMC.҉�P�J���P�В��Ì���t������u��(w/r�c��ju�h�"_u�Z
�·sR���a���w��1���S���f��ǈ������=9y�g舶Q���h|��P�yI��S;Tˣ�,�
g�v��qXa�'��à��4�`���Ӌ�܎S���ƹ�c$/�_����y�]�؉������B��*�m�ٷ�_��Y�����t|J@'(;�t�n\*o'�GG�8ʯ�t�'�³+�)'-g���f�������8�F��eD,��*d)��QV��(3y��N�8�k�k�<��|���+.qЖkc���QBV�TG8�%塞�ӽ�lš�.�c�M�����KZ�b��y�t���<2����If�f�$���Q�b��t����Y�U�2�����󰌾�8EV���f�,�|K?����gya�U����ͼRo?�|�v�g��ށb�ئb��7��{Z�ɍ��N/6aC�����$������ε�E����3�_̟eY�m�����n�p����ZǦ��&3�Ț?�g?Ц��e��/�~^	�CQ���eHr��S��)��і�i\��L~n⨝aR������9��u�yLy3�ajC�A_�x��oۓ�	gM+�G�e��6��2M�2/�2gZ����ӣz��a�]�%�6�i�����������\&��2�i�f\�q�{��*	y�(�'=i%8y�e�r����%��.��^k�@~u@�<�
	��C���G�F.u�y���L���g�[���3�,��`����{�G��W�r���֝��_C��H�`i�����1t��*���wnmGiU1j�����e�(7�k��aG�UB�;��;���?��e�I�7E̞�7=��3����'��؅+�J%�4��z�o}�>���r�&�K�y���(u�_#�1��xg�]��)p�Q�0��{��1��,˜d���r�7�Q�����oR�-s�C��@��u���/��z�<�CPwz�3����,J2d����\C��<��mY:�{qh��x%yr���ˋ�Y�2~�l�t��=s�4F�{Gȿ3|����w��h�w�|ϔ����@EЯ�n�ر��Β��n��|�?Q�('���*ؠ�c9a�/�,S�ې�^G/��r�� l^��+�.m��{���������a��%�u`Z�G��cPF}a��5^��@y8cE���L�qɓu&?�_�TX�3f�t��-��pY�|�K;+Y�� E,<q"���YO���'�:��e�I��D8�Ҵ>�7�S݄��N��Z�'��Hd/{�:|��G��W�c����Cg����M𺣘|�pqn˶�'������8�ۘ���c��<�	�#�݁�[�žVw��������kdݳ�S}�'��\���m��Їl��|+��M薨o�)����y)gIiC٘Ά�Y�����+;����5��y���V�̸���=��h�l~U$I�ނ����e8���@\�_�%���s��l���^T�2lN�.S�%\��s
�p�.O�t��x���J+�����j��|N�5/�f�r9���4��gi6��g�u:D"��(O�e������fX3�2g^B�?�y�20ސ�4�*�A$�K��GY�7x�cr?:/��綒�.���H�\Q�ܹ���:'ɻ�X%���n���뤶Q"j$g�n©zן�ٟ݈�>�r�0n1F�p�s��q��{4�0Z�q��=P�%����:(�Y�ߐ�?������/�XA������>P|#�N��ۂ�
��qi� U�޳(�!f^��H���t�MS��*��,��۷��;oFvLN):[e��C�w�!�6ʽ�c��7�2ȫz�p�J��90y'u���5��K}vp(�{ ���E'&�vr�<^X�#�1~�l���^�H�i���H����y�k~ۡ�m/:K�O�0�������P̪�:�a�Ɏu9nod�>� ���)-��?϶7>1����511N��lr�i6��h�L�勃,t$�Q�J�VG�{cYT��w����,�� �7��	r�%�GYfc���q��y��F���8�7H� �p����z)�*q� �L������aŋ�gS�G�.���D2�,e�e�����l?u|�8x���	sR�"(�1@a���J�%�+��f�vk^�Q�ȗ���<��J�Y:��r�e:�{U�_Y����lw�5�q����b��k˓S'8��b���G�O��s�������V���o�z<���Bgqf������ӻ��@����̥;��E�[������nڢ�C�RC"�h9��w���S[�m�	pq3v�sM/������'/�4�W�5��p���m��~SǄ�.n� �t.����5��wa�U���/�W��8ie�'pA�r����`4�{�mW\Ұ</j��d��_�ƽD�����uz��̏�B��� \�sk\.g�#L��c��9�%.�Ov�}6�K��7����AQ�v��sP��&���yt��L|��l��/�<�	�
��zx}I`ݹz��� 3F;z������>��Xv���琌�8[���v�����Xłq���;��r#���~�8V�0u��`����ĉ�{A;�7�b��g��Ԏy���L���8X<�s���#�{�#|��?���D*v(���1a2u���GX:u�:�����!)����m�j�g4F�EpV4x�mQ�a SזǢƬ���%�]���}��vFz2ԣs�Q�=�?��ؙ*;Y㕗��!O�<!x��z�S�:��3��@,i��Ʋ<��e:��@�|��������9qGYq�p�0�=�=��Xg����S�Aߙ=�����{~*ܝ�e�;?1z-��`v���|�5�0���$��5�B.�
9����0��7�21B�I�����|�gY�yY�*d+���@n>~Ǿ+�Ia�йqv�z�1�g^Z~��o$�PKY��J|�*8L�!�V��ue�Cg9�/!O�%�!�/�>K�vE}�ϫ�'��rXf�)�/�"N��]�A�|+m��F���dJj�۳�*{m��X��������tW�塩�ž���[ON�;�g8آӽ����;^L>{���XLl܎|i1��%nގri�gqr�/2�(���8�aoap����o���'>�.��#ʬ����L��� T!����WF�w��zN�f\��<�f�K=��A�͘��:�h�G�S��ʚwܲo5n~������r��A�ē�E���tr�y2�p��ĴW�s�&��/yB��:I|�i>d���s]���Ch�5�� <��Lh�����G�3�S��}Y|����J�+�[<��'~�Ƚ��t/��"�S����+��T`!,pі|oy��0/�P���+1��O�k����u�]�Y��O�&�窜��:���su�W<��u�$q�>��������N>j��0�#���p�B����Qw�<[��C�q�F�<��g����������K:V�������(�o��n�P!�{���"�Y�D*E�F�u���g�!f���t�qU�x��[�x�č�1�訽
94;]㢳��"�;���z�:����Np`�-�,�Kۺ�Z*0��11�1f�(W�?�j}{�-K��<Z9:9�+���y��<�-b	�!/Ӎ�f�R���7�s�/�uGo�m����(�/6mڈ?Γ8�p����3��#ۭQ\��q&�a�kԻ�̲�\-p'�2fT���ԉ��u����a8�⻪M!���q^ʵ�?��N��%�\��l�te�A~�����H����^�_塜s�g�:$Ň�d�y��z�gg~�q�MX�Q�(�e6�r�N�G�m%�)�v�����b����L�s	��=ټ�<����z�4Gf�/t�P1G��V͞���N�,�6�f��Z���p��D���(k��0fu��T�~係
c�)q=��+�؎s��y�o�gv�]ה8W��ۊã�����������c�[8���sŹI�����aj�ױܰ����=��.OMμȰ�/=��������
��
��!D��8����֕�6�S;ƭ	�wƤ��Mpu;j�[�''�t����b� /��<�m�O�2�q�DA����7NW���ۺw�9��&�)N��)>��H���F�˟�3-�q��/ᤕ��Zn9>�6���8�3!�0֣i�n��<GR���F��¯��<����u�ʇ!�1=�#�g>e����e!�yr�x^����y3N��m]��+t�6�:Ȼ�|	�`�f�W�a3�K�8�	������+��:��/z����?�	�;W�qU�p�6ё���W?���'ل�ѡ����#�i�~,er�[��(0w�ݺ��@st|�4���]w��w�����-�Z_��?�×���w������ϯ�0�M��0x��S�3�?���<�-��~���{6�@���+�~�u��Ё����A��0]�t�����w��)�	�����G{��o����c������	��e�?���\����)WuB�m�`��|�J��v�\��R��'t����@q�@C�x{i'N�@m����x�'��G�)�����r�\z��O.�A�q��ٰa#�TG��w���8��'@~���[7���?�o�%��p�p��p���'bMX�}A�*[�2$LÁ���D����w��ƅq���S٘n��G^SE>�e��)ߨ#+K�[^r�8x�o�c��r�[��rȃ�`�a�2���������JZ�GɠB,�ܳgO�vv��A�c���z��u�CN�ˢCg=8��_��Jy(7�����ۦ����g�S�e�3�Ԋ�Fu��[�b������3���U��l�����`��`l��A__�#u��Hys��x�����EX?�Q[�+���=�+��'O�;��
kX���� ��v���)ۇ)�z����g��{��{L�m�\'\�)}���L�Ae՚����{[�<�z_y+cq�{�+_���]��w$E=*Xg�d�S\x�j/�83^�5���F\]~��7�Wu\}��(���"l��s��>LW���_��ND_i��M�g���H����Qo�fzw͗��3�E��y�p�(n+7~�N�/�$-�g�)�Ɨ�|��+X����=�	&��7��*�������y����&��������i���Gf���������ѱ�e%�Q�6����G/>�Wu0����נ֝��`���,� �ң,ɺ������/|aϗ��������p�QR��(�J�=���Q���a��I���^�f�����_��_��\����/k�3K6���}�}ؿ�2r����[W'M+;:
~_(&vt"�9{�-�<�~��2�|�G�˥��zl�G�
�p���r�t':4;��������K�9F��r�w9~��X�y'ˍ~�Ng7m�*���4��)��:��vf���;�o":l;7�Iy����e)�`���h;�i�k<�;fW�$����%�.!X�$���v���04��ƶ0�.q�D�L'=�D����Hw�^̴iLW|;֎�J]���\��0����'�9����a�Sa>��ey-���t���y�g��!K�� �5��2X~�"�V�Y������Lò���v%�K��^�Q��6━��e��X~�YV�-�p�a6+ڷ��#���3S��A(��3_�q&�}�Q&��2��Y~�N��qR#�8�#��*�ۃ��s�1,�luu:p~�8=��-�[�X�7G�#{�Y6��O�=ڟeQ���f,��{�fU��$��A�Qt��*XE�2?ݝ?I�.���Ն7�PϷO�.�(ۖNO�q�U\�}gq ��b������,g�u�
�P۷��n�)�3��N.����]ԛ�G��,������aPr��H-O
������6�=�3#d)>ꊄJ8�M7�{����Q��r�h��)����$\���O���x�&��Y�z$=�%L�⽎��pQ�����Bęn��������/ӳ�)-���y>[~�&9�o��U�4Ǚ'_�hį�OR�\Q��3$��̟�mg����	�:Nz�|�9�]�π5O�Ix���l����n�����GW��~N��.3�/�Utb��o�5ڟ���^R��z��_݄ni�����1h��>��.L���?�W	�;W�YͣԊ���ފa�;����,�q�K(?Ll��(��-]F�c���K�X�L4�P�y_�
�C���{��/����p�^V��˟��n�C�o1�n�x�G9f�����n�iPхa���(��rB��Ї�$�{���KG�a@^��r'{�<�=+x���u���2�N��y�ް�Sz�Q�W�C��!��nx�op�`4�Z\ڔ�h��i��X� ���+���eW�:K����0����vx��F�@;U�٦t���z�M���}��8b�:e
̪�g�l���%.�h������rC�:���0F��)r15u.hˣK�ԡ�A�l�0�O�ʆ�����Kc>;:�E��4��NH+ډy����̯�H��˶���G������^���*{,�Tf/m�s��-��By��8�����7���M=��"�!�D����({�HXq�T�Ǩ��rx=���z��YVi�ρ#ˤd�Ig���И�zA��,��on�%��8�v�mӦ�q����8t�9�Xv�GyXdee�Q�qZ.eE`� ���L2H���l���
����ep���\q����ޑ>6:V����9����Do[X.n��w,��+{�����<u���g�׆M��y������o�k�;��#ǏΟ{ÑÓD�|���LL����vE|�x\���Q���X�@i�N��1$��32����u|�'�:�q�w����1m�ŕ�Q��{�Q
t^���{_�ub~�qE����,�9��L����#��yR]G�K�ig�'D}0^��W��M��[��rH鵾�.�ő0�~װ�7�Oz�I�bAx��7!�*_Ο��qE>�\H��g8�m+�{�N�,���f�7��;�y
�p}��,��QG��y�/.u���댋���I��X�X��w��ݱc�#�X=���s�/���l�^OXw�.��FA�0J;r����>��O���q���l(�����`i9���BЩ�7�?���*"Wt�D����g�Q�VV��	��W�W�,G��dj <m;�v�c;�!����a�F0O���?������t�sGi0�q��@n�Yg�P�3f����uGG`�V#�:����γOm������6�M��^���ۨ�8�.�pV�eU.�Cװ,Lީ��Ѐ͝r]�Zm�:Xβ���N8�D�G\a(�l>;B��0Wɸ��e��Ʋm̶��4kԉNV�,�D�������#[?";[���'�b6˲m޼��o/0cQ�a����r;p��`�����)��K��8>Jk94ʽ���w�2�c�)m!ff,��a�ӹ���a��N<-P�%Φ�CBc���)Ҫ��%q��F]��ț�S��CP�W&��7pF���'Ņ�P��R��2ζ,��8>�.e�,,�u�e���?3%FY1zL�3_Q�.�s&���F��G.���-f�t�t�u�(k���������/��!��UГ7��'r��P^�/��y�x�.�h���h�3"�c�y�C�yrf-��N�<?S�Ȇ�>x��ٲ�8q�u�����g�ϔ���Z���,��+�ٚ.Z�����;���g����:�2^�Ӳ������G� ��-�eD��)�~��Q���{�ˮ�P�ԩ[�Ʈ����d�Mq�EJ��A٢$�E��dE��,ۈ�� ������Hg���=�F<ȖI-�Hj�8���3{y��u+߷�٧oU7I�#���O�s�^{��מ��#l6����R/��o�p!/�U�h�L�ηrH��;����@��F
��k���z)�Mm���xX�7BT�ȧ�Gz�ǔ�O�Zy�[���MmW
��z�_�?��;�0�� i�H�h��-O��I�%l�5<��d��I����K���Hp�;�q	dY��'�W�+N)L@�S?�l�K8�S����T�?�� X�J��n���h�l׬���y?���z|����:�������e���/���K��_�����Ր��F�W��U.�)ڵO=�ԕ\
|�>�a����DU`T=���b���ذ���F�S��4~�ޝG~��~o3V�hX��U�����mh����rb�Ɇ�CŎo�WMh������o����s&��Q��	�����7)�"F��/�n��߮g��%(��ߟ0#y?3WŹԿ@Y�1�������c���(̛���,a�5]�E�Tt��mi�ą���e�G�g�,>*�vxvt�_�3�O�b(*��XF�G�2�"�����R#��̆x�2F�^���*��ј)�L�7
�=�X��?�f��A�/ԻX��I���%�aDP��#h@��{����]���1c�ү�/������߿���)��3:qjȁ.�q?G��3N��ƴa=��������eG</Δ?�E�	���~�R���|R|�8�Rl�y���
ˇ��k�(ӢA)�*��]a +ڐ8���)�ߴ�C?��oa-#|��$=�Qovv�P�8�u��L���^��G�����Y�b��˄1�܃�>$�X�$~�i�Oi�.hKC��G&���X����n�&����\6���9�i���'f��v�yvr�������/�&8�dhq�9�A}�^�j�֐��;�Me=�O������F��W��K��Ü�����x��ޛ�8x�� �J�WN>����6��K'�X��ڟH��7�+ߑ��=��qW�[ir(���
k�Qр|���29g�	�*xd
'e>ʬ�e}��g�2M�Njk��)�'��r��G���0�)�A'��w���?�H�-c�<S�G���~''\ȼ�_ƻ�������_��h�[��g�I��;�������o\����F�D��ٙ����|V8��K�����<�i�9�,�턏}���6^x�����W5hw���&�Gq���ݗ]vٗ��1���wF�[uoz	��!}��WU T�������_��e�L�ܹ3w)����@�	e1��b��FqmhhH�!�a�Q�8���Y�G���oQ�_��Sg���O�X] >��6�%}6h�q�ot��K��n��4^���U͏��o�ߎq5�~�m�a�Hu��P
���C�IiU��[t���o��_c��/Ը�VJ�ff�E�{
���=�����(�/��25[l��o�T*�a�\�I�עH�:ʣ�X�1SC�eU<�����Ђa��J�yA���?]i�Ō�����d��g��pep�T��?�N��a($�-�{!N��1��R�踇���#�Mzҧ�4��X�{�L�4M�����o��*�H);Tڕ[�w"1�|{H��5�0&�}P�ؑU����?ߡX�['_:�H��H8�;`	ë�V+
e%���|�F�a4�𘙲ͱ��\�2�����>|U�\^j|e��Wn�'�2��%�����#���ήndQ��j�<*G��<�_u���7DZġѦG����0^cI'���)#���#O��*��5����<�z���e���c�����f��wu�O�dM�gS͉li�/��퇧�� �e��v��mq�9�R�v�|��H���}$��ɮ���uy=�q�������7t���#G��g��F�"�)�ǒ�U��N��Sy6��(�����*e=�iU��ۀ�w(��6�u+�	o'�5�q*������*��U6���m�#<�l��)���2R��L��oq'�Iǲ@Xԅ^�#��$<�K�c����w��$xq�p�����?�Ma�V���.��/����D���N��������I�O��׊3}+C���d^l���A�8��d�}�~
+}�D2����&\�[��4��:�»�����GO���BO̯�W%�V��7@1��@�ފ"~�/�x�P6D� �D&e7s&�QoG�9��#:�UV1Q�A1ň�g%��Q��5?�8����W�������5�P�JC����0x<��F/���O,,�5;�if��q׮]�d=��z6~e�P׳�ꖧ�~�
u[~;eg'�B��yo'o�&�楗^��W^����⠩�޾�0����P�5�,;���<�C#����H9Ƈ���X�%�Y���Czu��k���g�2>���!���ԫ /��i�h@Y��L�#�xv�6.kD����a��cԥ?���^��A��vFBg1��n���3��i�WZWβ�?:s�ƞJ�Ɯa*�<1ۦ�
��ڷ|KG�qE8U��x���/9A�˔�c���h�E�w�P���[\�M���o�W1�a��^Cn��t�5�9�  @ IDATn�#)n�,N��'e�+��)n�y�3[�ѨQ��!�Sz~Sb6Ox�*a��a~۾�oMf�0D�A�P��Q�⑮y����ڲQֹ8�P~Tڍ#����N
kڤo:R>�{����v�O
�/k�诹�j%o�Y�������ToC��)�evmb�<�ϻ�5�X��Lf��������Lv�m2۹eGvۍ7g���Z���>מmn,̯9~�wϋ/�Wy_o>����^6�^u!�ô��E[��y,����ʷ�q)n�o�@<��Wȯ��ڇ(C���e��p�w�:n�O�G�������O��?����S
�wȭ�q��,G%|�%N�B��q��H�q|���A�-����'l���n��[hV�+��W�qZ�����$�py_����+��fۑ$?�[�/��;�o<]+NaJ�h�����Ǻ_�-�e�e�U��Yܴ��5�Zr��}�ѣ����=�����?oj	�Wo���D�����oGI�5�.�b47����G��%76.�Q	V��+��Q�sX��p��}w�q���B{|eG�����������wĻ�G�H%7�gC��lDi��W���2ʱ��f��S�i~Si���9��e���3����	e��!̽,��i�4��a<���/t�
�w߾}W1c���n�S�3*�<a�ۑ�3��S��3-�},��s4���fX�qF���1��tx¨ؚv�	��/r>��TF�+_e��X�b6Bz��J;xs�ת|{����&˹3IaKũ��ԥأS��g�IЌ��ʴ�y�Ұ�0��]\����|Z/�:�˔N3>C��T@��$��S�5M�'(��̟�%9)+q��2Eͺ�<5D�X�Y(:��F�/i���}�:��b����dk>$CD��.Õ3e*��?yS�L~��;�GCԷ�ũ�lsL�y��o~�q���*�8坶�Wa?��͉��<���s����o��2%�<���M�&�:�Tľ�)��l��R�owgw6�I�3�ͥv�f61�Ef��ڻ�.�n�|����'&G�v�Xǌ������d��ޙ�&f�u]��w�޼�W�]܉5��է8�bzr����#�˘�;;�6�a�-��y�_�h^�G$�����p����3�/|�e�+�#\���
CH��;`K���p�~Qv�#��'
W,�.=	�0�!�X���w�W�$����G	���wJC�/�T�ŗ�~(��R�$_���
�h���g�Ore�y�S�-3VZ����&NԿ�Fa}>l��W���mܳ�$�%\��q�V<�Ņ��o}l�,��^� �����$'>��a�?�G����^[G�o<���?��:��"�nP���8��@t��`���p2�׀ݟ设W%p.	�W�ʯ�Dm8˶�E�������_�s��۟��z'l�4��7ڛ��&�Ge/N1?^��&fb������UA�D�R)Ѡ�����``�ث�~:�#���_���(H;��&P�㺍����J�a(A��{�VOs��n��Ǆ5�o�p�?����O>�T������ 2�uG~92۞s�6�+�P�fgb�VgW�޷��׆�e��E�E�8�������3"~�����'�'z&&'����M��ϻQH�%�82�i�!��{(�$&��:3�W���`[��W(����a�i.ac3@����F�C�
͹��|��jl�g�9-����gIX��Fy���
|(�*�O�}t��!��t5�,����j�h\��z��
���7ׯ�2x�w��%y9J�Fp�Aq���d�?Cx3�,e���ݩb�DV��T��W��{�f.ĭ``>)6��1��2ϡU<Ŭ����xq�|�o�����QfYj��.�8�.�:4�{a��`(5��1��]��H��M��z�ou5��MmBq�L>���2�u[����gf*�PY�mTh�auhҕ�ƺ2�<ɷ��Y��0��9]q�et�uy+�	}0��#�v�������)�HEݥM���ɬ�(N��'�
�K���H�ca�����0��jЋ��1X ���BZ�Q~�����2v K�,ǰ��4�f9��xf�����l�tq����8��&6P�D����Y��!���Q�h�X�z�)Ӎ������U�_�\�"O���:~2߻~zhx��{���.-�8Z�:�.�a��V�4��R9g�0U��OYL�ΰ(+�҇Kʲ �m��,W�_��m��;�9夼p��_�6=� ��8"��˥�|�ϛ�9\���ҧ���.�_�<�j�K�.���I���P�ki|�ś��S&�2=1�,l邾ߩ��p�V�5<�!<d��i	𐌪�vɗh"����C��I��������7n���x����_���^����.������A?�'��_?�EC�wپD��'p	k�o� �����'���ǀ�߲�ڸ��_u�x%	�W�$�_��,��\h~������~�
H��Lc{wOmM�tv'M�Q�5=��{����g1K#��6&*7�l�Oe��rc�A�t�w�w�}�m��~5qxd�<�����F��tV 6�*#�eu:Q7��	�!����Ν;�����_|���P_���z82�!�~���߿�� �S�#���zF��TpT$8����? ��މ+����/~�k��S�L�x�v��񏍌�����X����L3��w���9���Y5�5�2�(K|jhә�i��b�J�Ϣ#&�0Je-s&��U����.�^"��t�$�8����,����:����Y�u�yt�I�O�p��jx��i*��㎈+�.�܁��
w��Y,�u�<uq�+Js�F?xY���	ø�Yo�t���Nf2T�dn� �[0�M��)�3<Vᯌ524�H[�H_A%�LC��k|˗�7La��Ð�8�q}��R&<��:e�a��:�<�8��R�\C��d�o��k4�~�(��[c.��ӄ�Ӝ���`Bg�	�<q���7�!Kz��HS��0tf�f#/���}i����55��� /�����_RjST'�W�[YG^,3�weE��=����Ai�/���)?��Y;�X�^���ɦ9]p��.Y��~E�YĨγq���]ؐ�t�͍��qU^���s�q��:��K���gE9Ѥ��rk2�*���R�%�Çe
��VӢ6�E9��),���_�~E�)�B�|'�7ȕ$��2��������a��r�Cb��������#�3��'X�?_�"���cyK�)̷��_�~!��Ok<i�Z���l��p�J��~+.���e�_ҋ������y�}ȿ5����*\-�����>[��T�B-�Vr��<W�a�7,=�U�h��q��bV�l��e��3�m��ٷm�Ǻ*^{���_;�j������Xu�x5	�W�&�_�p[�.��+��G����;vt��C���/��f��maDs+wW�"4g�&�(��0�~��l��\I,���h8�L矖��aE�T�4L��y��V�v0"��|�����
��XFu��.��c)�
����J8��M��o��_��V� ��B�v����o=���9ҍ��	�n�4?�D�k��Dqt�r�p��7n<��z{�^���rW��s?��ĉS��qbb<.& G@���}�"�.�W~�/N�_��݇0��c����8M�ʍ�~;[dǨrMY��t�S�ո�jXhx�n�ŝQ(�a��y.��E8��"����c��T�(���ʔ��2g٣?cy���34�U���8q�Ď���S����.���q���S'��q��z�y���.jo��-�>�{�qZ]ѩ{W�iD���Rȁ�k�y�Ba<(K8�.�%�%��0�O�WvI�S^�/dF��>�1�<�C!)e��տ��
�bV\>�/XbI�y\e�*cٖN�;�e���>��x��)�E(���R�����ǥжcċ�N� -'h�!fڕ�a2�4|�m3�z�[^���8�O��<�g9�_��j ʟ�$M��2��`���'��q�@Dq���" �ram#3X��e`.�b��|y�<'$��nq]v��H��ߝ���j�77�ˑ��Ƒ#��'N��T�6&q�e�+HS��k��S�-�b~�^u�ռiyB^x�����Mp�V	��K�^?k������K4�wx³<�_��x��"�dL����E}+���-I����ʐW�%�z�-��F���ҵ�U�-+-0U:����L�|���FU_�~b��V\+���W�[�~���)^�W�&�<�K���Ð���	O�)+��[�l?�S���N�6�t�����#�P�'Ю�S�G�G����oڈ�����^M��իI�$�F��C��c~r������kN��;{b�������l���=���H���ksӍ�ӣ���٬��6���l��8��E*4"*-v�6L6<*�*Z6>4bc�c�ދ������[Ǯo|衇n9t��}6�*)�ǥ�6`4R^,�h���w�g(.��9΁�}�;��a���s�O�m�������?x���a���ٹ ��T�c(w���vr\�7\�gǎ��X�Yl\z}%X��̓�o�=G�U,�ťa����L�'�j?��P�M����m0�}���>\(�~�\[.�WQe9{P�UB�W��>f ��X�K��oG>)�*�v�,<?�U�]&�L��]��}a(HC��CYq��rxB�y�� y� Bo�X��4�)���$P�A,��a����n�&���dDҔ������,��9+�q/��E7G��H_ލ�CU<�Y�lKy�?��c�I��|1~!�Pbw��Q���C^⑞�~ˇ<���m�ݙW�g�)W��Јv��%���֨�x���G��9F�����̀O��ۙR��0T�K"\����(�.��P1a����4Z���%\̨�Ne"�I�4KG���>e*o�(S�!7q�^�-��uFX�=a�y
�1ԋ=!.o�aFk�U�Z3�0��T,e��dƎ�<=;�]y���{��`��뮵����s͓C�k/>D)q	)3oUMpָ�������]�,������u�<1M�~�	��ʪ��;��?�ek[���-O�6}J\�o��lE?�n}C&�o��?h�?������gɯ���;9�M�?��	$���N���y*~ %�s�6��[�U�/':I�/K��a�=�_��;���
�w�I�i	~K^L�^��R�_�R��.�(?��B������� ���������!�s�97�ۓ�X���:��h�;���?�xe	�W�,���Cm(`�{z!�bi~�����Ʊ����s���|��%�r�Ԯ��7�7�ךӣ�cG�/>��6˪�����~Z�ǎ�Mv���	�;��m|h�Xu2W�1��Br��8ҟ��}���l�^�<xp�w������G���Za��԰��o�cc����+4��^��<x�w�3W/���ޠ�������Wx`�y�A,#[�yOt$eǎ��T�#�BY��?o���]���?����k6?���ƒ��Y���ѻ�8$ âǼRYuɖ#�*�>:�i£��,�Bb:y%�oˁ��
z�P��CX��l�AZ�Ph)+���G�^E^�(f6 �^��,O�ko/�ygt��Uw����;�b�	W��隧P�9:}T��;??�!U�%{33ΐ�$ϓ��Pĝq��$[�xm����~���_8�ue`�o�K�e��;ϒ0�be)�3XIA���N��S�I���$W~��b��/��I��x�3�2D�I4�9ʟ|�g,���(R��ʊi4m�WAƱOK�F'�җ�_Y褭_�K�{f4���+}�3����1��M����?3;F+hbO���{��ka�KR���N8�a#�J�E�I[u(�y`y���H����*KF�X�{�B��x�O"��rf���fIi�.���&�00p�[��?��Og7�~{��oM>2=���`~��Q��Me=k�ڥ��5�*ߴ#-g'%��-s�Z�[e�d��~��������J|�[�yr~KBÔ��N?�[W¼*tÀ�|�\ŷa�.�_�86�H��9��_�FZ�O��	�	�+�����\�� ���VYǷ|����[�k�K�ӻ,}�+���,�Dl�Kx��N�|�3��#��[��/dnZ#bI�()��U�����1��9�ښ�']뫏�v*.
�o��69���;v�O�$��qխJ�5K`ոz͢��������Ng׺dәg_P����C��>��/6O�47O/�oݸ-�����7��={���7��đ�=�c��ʮ��[�磣ۏ�טGc�C��ï�y
NC%�HeOi������ �|%�<ᖷإ8��gu��?�;'OnF{@QRy�5hkvf�f�����[l����ћn��!�z�C,�e��KG����m_�җ�߳{z^�f��,�;�.T��p��S���P�jp��Ȏ/����ֿH���	@���-,�|����o�:u��	櫆������ک�X~J��4�˲�qy��.�b�.�Cs�}:�4n�\M8��z�E.�5�a�kH�س/*h�S|>R�7�lq0�kD��B1�RsGymfk��I�&�m����uf�j�͑af��V��Y��l.ˋY1f��P�'��Ȣ�����N���qߔ��:�m��f��j1g����M��T�I�3o����:a�R�,��h�8S�2�( m1��SZŕ��R����Hxeǧy�7��3��_ɜ�F������S�O#���q�ӉS��KO�ɘ$n�y3\�4B�G�̑J�qh�s�Йn"C�<���F���Q�N��@�*W��	��QN8�3��[^M�p��	�� �c-f�L�pQ�K�E�	��gi�7y�4m�By�C)� 	f���l�|>=��(,�\��5T5��'F�Ν-e��i<ۼe}��]���n�)�a�ߩ������}dS�Y��-�Z�;i9s
/ML�(')m�#�����$�<�!�W�1��M�1�>�2~��G���O�����v_����(0�<#exT���/��J�����1ܴ�D�Ip���J�0z�+߭��[�����?A��oY��ߊ/���w��i�wV>�+���^}`[�j�Nl��
���%���e�L���2M���
0�!��1��6�m�U���.[�l?VV�T���Y����.���6�� b��/�6[!� �O��)0�nU?�V���N^�Ph*�=C���k�6ߝ���?x���O�^����/�8�������-m�%��6�]�w..d{{�~r~�953���Xs�U���ƾ��y��Ŭ���{������M�=��l���RAw�j��n�U*7�g���?Ĩ������z��ǁ����O\��o|�������P�Oqo�J���Y4|�ţ����Br%�IN|v׮]�ķa}3�ޣG�����|�]MM��N��
��@M����*��F���ﻗ\x����s��tr.2����Pncrj�"fpf��˨�(�*_�G�-)��uvdɉK�}L���-{�1�J˄p��T�2̎а�Ngy�{PT��e)|�否qt.�sϓ��0#�	o�}�a�t�x*�<͙�g��ߙ+⡼ƽK1[�m�o*x����Br�i��wf�8�3&�ɸ09��ڜBѵ���f� ��̚1�׉�2�?ǻS_��3�P2<	��-ZӋ�B�)Kӟ堟r�?�o��~�C�Xz����'�8B�1��&�f=���;��{Ǌe�� /K�3S
��ʼ�4Z��/NqK����D̘���.��
�o˔{���oi����,9y�[��F�D�ϸ��3
0���	g��1\g��R!���od�/6PvCw�H���u�wc�Y)eY��>�L2[5�\~�e��?������l���~��������)����%iR��fB�&-˚�3�3��Z��s�$�PxM��+\�Y�݂c�T7	�x��D٦��U���R����?�������
|���f�^�9��NJz�a)m�~a[��SW��G���
�p%���J<����;�Z�ē���8+�V�Nil�O�),���N0�~��^g:�-��w*c�p�;pR��>�y\��~ɰ��,��b��v���3����V��q���������`F�����#��U	�v	�W�]V�H5M7��XıPͼt��'^x��={�f�h.<\�89��ea���~���l�6�f���'��N=wr]��>��������ٵe�HϚ���F��x�v�����F��s�U�8:��H-
�<��x.홥�ٍ�p������V�E�#���t�����?�𻆆�c��� Ϋ$���q�n4t��^,GFef��w����_�^�ظ����޽���}�kw���m(^hG��~)�y#��lj��@T��9��g���mߵ7^���o~�F���j#��ap|��ʋ'@Ɓ����eV���_�t۩���\ѡ�&~5�a�~�:�(3v�!�˪�юѱ��TXяC!�#��dZ*~���x�f5Ō���t5�{�X+_�4M���..˓vi$Ĳ���'nD;[
c%>f�ٶm�Kc/�{��^_��e���qV�{�(��Ό�Ǥ�qg��0
��� �a�oK�/։04D�AL��!�P�5@t�%�kL�.�l�r6-	Fy�g:����L�����Ra@%?em�<o��gBA��DW^4��y��֘�-#�#&C(5�� �>҄�S��o�X6(��,P^J�.ʟ��[�FX�!~�L~�3}�_([�@�OgZ��E���j\��(��Q�#N�`���/-�RĀh036�R�If9�3C^�)�+'"ƒJ$��	9�;.ؑ}�c��>��{��7d���1ku��|jt�k0�8f~�1O�s��6���d顬-P��{9E���m�����|�Z�J\ˌ���<�)�m�Iag��P�E���>YO|�bf�M��
�r��/��R��8���M��R����ģKohD{��R-AU���	����^�7��0�RV�o�K��&�+��Q���x�a+q���M�\)�S�O�KyD�E�4�|R8u0�	����G��?�,+>�ap'�'�G�l��)��}V���������~	�W?��^gX*��}3���sã�=����N>�b���/�\:t�+?v<�����T������j�(�������lF��ё�nZ�[?��_�е��Ϯ���:��<q�x�#O>����� W�l������u�>"�!��q��x��N���)饑��~�+w��]\���g]��I�uV�O:n�Ν�bp����H;G�:���8xNopOd��LХ�<�ܝ_��W6p(�'Iu�*'���g�dބ��R�L�pf�n�|��[�}��js�~YC��%�ڞ{C�݁A�oP�/��.�Y߸yc0F������+� ��=(�By��I�b#,����
���QqF�N؎�5��gŴ���j1�""�)�D'��0�AfaЇ�om���B�_j�&fFX�����	��Et3�R*G ��� �G!�cHr� �#���0Ĳ�I���Xv�L�ʟ'��O�`Vy�~�k�Y�\��|zj�937
�F����}K�Vy|��QQ'�0x�Ew��R�B��+�^ˈ�@���!}��Ra���8E�8ʔ8���2� ҉�8���� ����Aa�}�O��;�U�Bh��L�.�F�W��4�����o.�-�Xf���2i�kP�!%��IO�M��Y]�O~M��O+V(�*_(�Q&5���L���H��
E�߱�~����	kz��6N�Ic0f��_�b�<@�X=��?��kM���f�s���JIۙ'���GFa��zq���7�3�������훷�"�SC���{�S�Y}	rcs	�p�'�B��N�A �/��d�۟��N�M3��LW���g��3��7q�%�W\|We��Q�J:~�[�Bf�mƔ�D�/�Q���,�Qލg|˃"���jg����W�Y�8K�'�O�cz��2���N� V�>��q�8��~��!n�dx7p����"�L�����FI3��p������_��w!�"?���~�0���Oe$ߑ�O��'���0���r���E���x�-}��1s->�-������Oe��I���h`�}�������6�6�8�>�l�]���E]�Em����<��[���"�7�qE���Ƴ5t63�dk��6GP��ᬏ�X�A'Y���/��`���f��k{�͘_6�ˁd|�,R�V�����F��)n��7����̩���{w_6x��3GN|p����ԋ{���ᬟƢe�$�,)ɖjmg3\�:�S�GX������Ϟ|��ګ���|�����Cm;wkB
�����3s��X�ǎ�5��X8�b]J���E��J�6�J���Ǐ�Ӹ"=�j����t�#?z�m���p~�ot)�eܔ�P���k6�@:���a�9�"��'>�o�{�CȲ�-{��,������?x� ��u�үtY^�T�x{��LtJt0�詈�8n޲�?��mW=|�%�����ŷ�%�,�z+���o�>�7��n��T%bG�:Cx�:=���x�NW;�2^�Q�T��Ht�v�*��ٙzq���}L�%NZ��� q	�X��#�TI��y��sc��#�9�n��<Up:n������0�8��Hs�}_���Y'�2����k����O�P�9f=��q����i�1�j�S�%�� "i���u���r�ξ0&0V��G����2�t(��U|`G22���TXV�Ny�|����#<p�����C�\(O��3ӭ2c{�|���?��aN.�����U�Y,���HQ�8�B+�#͹wȈ�|���y�쑆o*[���|E�����o��O9��ĕ�.A��k��i��RM��7x�\��I}ф}I��� �Wi3ݦQ�*~>�|C�����?3��C���ϧg�p��E��.�m���l�<ϳ$P5�}�{_���ޑ]x�'�8�~0?p��䉓��>9f����D���V�D]AU���{����Kuҟ�	!�%L��x�Lo����7�K8"���W�,�H�2�N���o����e<'������P���?��q��0>�������wq�]�:�7`�3�˾��m�G忂�(S`H|�,`�S��sV�Sxz��KL%��/%���_��%�'p�q�n��� 埄۟��7O*�����*��)��8)Nq_^Ж��.x�m��e1�{�$�ڰ�ər��iP��^xᅏ�ܹ�{�%'���$����g��θ������m�9}��or �%y�cw��Ѷ���M۶��et���h��ز������n�c�py�.tc���ю���-v���Ş`hٙ��T��N����jix�C���&��.<�9���s�dS�����u�M�o�[���d��E���E�����6n�jlp?�8?�o~�~d�T~�b�����;���w�����C�*\���<r�{�������,sUn�p�ռ�K8��K�e�ޱ?��?\���>w.�/<���z��EQ��8*�*�6V��1�6�6�6�8f��)��c�C,��3���-e;���~Ȥ��������C߹�+�QA�Q(.�h�8㈚F6�
S!����m���>�/�d��CȯGzY�y1��̬�N�(�9���7ڐu���[������t	��k>� ^a�����C�=�O�^�ؘ	��҇�����j"��/q���a ������1�C���T�U���.��I��[�~}� �6���,QA&bY��j�`i�F�vs��3_����S�}�C16�^�����,��w�s��%��h`����5���1���eD^&��"��Q�!W���-e���r�Bo|�+<��C�i��0��3�FkRT4,��_�G��y���1�F�yQL1  o�
��1d^��I��o���ɓ����IG�Z{G
Q���믢d:�#�g�Ǭ���/_�K�+�-n�&?җ�o���<�;���B�/�<�g:|��#�V�5�<͉��s��"l|b4�����)�|���p⴬q�Mv��~=����K�r	��\ ̥��$��#�bf�����V]ʗ|�����:̥�BzfC�E�L�
��G��t��|�w�J��	.���H1oZ����q���!"�U���Y�\�/YG��x��2�ޔ}�WD=�o^��l��I��K�A���l�)K�X�Z��d"�<:�Ҭ�ߕ�f�\*��U�)��ao���
��3�)�h
7V�^F#�k����n�6����8���gx��e~�|���H��(c�w��7= G�d]���t�k�~�^�����e��`\�K���u�LrY}��$��2��@���Ц�?~��O�[w�������sD�#�Mf��G�;�:Ɠ�ôC�n4g�g6q�X���?�[��h����j��3���a�|��u[ۺk�6:�N���}k�X�D���6�0�!MY�����z��aÑ�C#���i�}[N?v�̩�9j�C#�t��W�ZK�%������������`aM�~bn���������O����/}�w��]w�zq���/���ĉ=�'�On�m��H�R�rI�m��o�0�Tzxfh�N}�_�ſ��+*2n�X����]��/�`�_���rL\���x�ҫrHO����ɢ�c����4��f������R`~s��C��һ]_�җ��C�'��p��3�l`V��m���{�ct���4�ӣ׾��_���Ob��&C��$|���.���Y
�qF�w��NG�����{y����0��[;�҅!-��ٙ�2ģ���y���S��7e#:M����U�o������ �_�P������H� g�J���ז���0BP���a��}��Ș��ޫP�9F$Ҡr�e�ٖ�[0P�]�T���[=��o�N>Ǹ�&�')��(;+5�v�r�b��3(��]��K
5��Tl�JbY)�pᔷ0��$� ����pT1��;�*/ַ�5\�+�R�1A��e� �d@�R�!��|34dp1Ȃ���"���1_)��(ƒMO��HQ�d�)<5�?�8P'f�T����O2.�`~�7i��G�|+�Em�F�*e"��a�:������7�c��K���@���3��jCi��5�TI[5'&g�����4�Kr8�`֍��ܜ��b���Ҵ��]������\�r�Z���,��¥��a_�ڪ6��vZjtp&��Nk�l��<�,�A����s�7���HJ�Ou���+a�?��>8Zh.`+�),p�)�7�G�]�֛���y��I��p��~�Y�M�觐_������<_de�$�J�� )�v0�A!��ӫo���+�|�o��i3��_��x�y�� %#���^I�ep��[N_]�V�����:��J�Oe��-Dl{l��C����m�N��+�$F���q���ǭ�p���3��S�1��V%��K�Ҋ~~T��֟?������j�񧮿`a�g-qO;�\�D<9:�u����:�c m���)�Z-,�5F�X���۳9�䌋f'Xt���ޞ5���f�^�Ȉ��u��͛��B��O�ă��l���(k8Ǘ�E�������pcit�V��'g�Mt�},/�A}bR��r��>;���5�����Mrp�	�秦�ONO�Zjb�@��o�������{���_e��ه�����نr`!��Ǥ��i�8�=N��[��)�Q~���%��#G��|��\��o
͂�SE��w(=��V��������={%z���a������@'���������|�����?��}=���k0rC������O�eV�#�׎�|�䒋�~��o}�V�x�d�Ap!�͟�g=��7n��;�<_&fXֆ�b�B���V��R��5����9��Z>PB���B�^�V�~�Cx��hQ���;S;Ug��=�8��,;�����e	\�5u޶�XdF.�a\����0�>�g9`��17O����f�����ܯӅ��h����֒���xu�p�4� +�BөR�:e��"\��o&�U�#��9��)��GY(o��)����_Y
���tE��%�(�iF�#C��8�8���G\杆N�mX?!i*O�S�c|*�u�&�ew�P�E�Sq�^)~܁E���Cg�u�w�);�3�|�F��8�2�B�!����
#ֳ��0�yJ�Bѓ�(;iʇ�08��0�g���rj��𚣟������
˅x��9�\������#�g>����w\����z{���G�?�8����0�y��6�ZT�T5Hxl��:aV�HT�x'��-�V�Z�㻄[f����o�eL��Ov���/y�+���u�J���\�iX�]�SCY�`��β��KO]�q"�-�~�M�%����~��R�V�ɏw+|���t���w�P�*��K���
�8�I��Ɲ�]
�]�&\��q&�š<S���Fl��U�+����]�e�<�'���u�o���� �n��w�>YS6c��x�����yX'�߆YR�0�G@����IiխJ�g��Ƹ���^9?9q���腋��=���c�Y�KL�4�ڤN��ǝ6��gIFc��S�x;{X^A�Ԥ���"nV�04O\F|�[�8�u�۪�4#�5����iF��(�%>�'3��ю���FP�8�)똜��L-f[ѣܥ;R�f_��..E�eRm��f4�z��&���#�3�>��OG:�I�	����n�������]�����z�WX��<�Q�7���f֮oA�b�C���h|4�"Ұ��)�a��Bc9G�b)�Χ�|��G�����4Y6d��Tg���aC�#nFۣa�$��c���=�������o�"��_��W��@ݤA�Jj>��!υ�U�^��Ѱ\�$PYF�D��m����o������e���wN�g�}��b{˩>̳�,;/F�r�[�G���S�&D�t����'e�[��2`|JaJ+F2�
���`�&�����#��x�|����1��4O�Z�*��**��	�)�ai��2NJ�<X��}8t%f/�`6���XV��щ��qB�	ih8#����5<2��2�´9m�l�۵������o��b���1������挘���a�(��;�ȷ�ąrb:M�3=*�+'eLF�>�2i�T�&cHy�tǌ�a�%?"��P>�����Q~�a���'O��iO_�,��4x�?/i��ae'���A��'~�,�=Q�[>�O��{C3]��{Y�"��/�N�M������n��+����T
��Vn��p��X����R\�S^�͖�vE�dB?#��bvn6G���ַ����{v�'�,���ɜ���!�F��)s�q{��0�y�>���T껿�xP@��c�bP���&E����OY�L_�������7�>:��V<!c�B�rLp�qJ����v >-��	��y�G��{�*�DGX����*��ү�
��_
w�&�,��ET�K'�3��߸0J㣔YD*�,㻄o	�t,�qY���s��K�笴�AY}U���Oxx��4�J����y�"��~l�=�N�	�U\%�׺���V?mR\.mM��e��	���&l/�Eፘ�V%��I�a\���^���\��w~��]?X��=�h�1;�wtf[.�ξ���ҝ�x/�C�j?6x�Ә�g�<�bj:�����8H�P��ռ�#��;jLC�e�-������umu�����X����A+笈��|si���~R�;9!��~�����*㊪|�ޞ���h̡YͣL1r|�������͑Ņ��ɩ�D-���S��sGn}��_��'�Y?N#`c�j��ƯGYx�R{g{����.`q���1�.��Q�Gu�efȹ�O������?��,��bZ�&o��F�QLb��NNW�`M ��_�v
����.����s҈Ho�?G��衇��t�w`�lsՈ]b  @ IDAT��4�E9���['C�\�=R[�H@	��Z	��yqm���͛_�e��K?ti���y�e�>��[��o�p�B�ݨB�Q�aՀ?��[(�ߐW�
��R��̢����CD�ȖP�1�Ji��F9Q�����؊;u���x�Ҝ!��+~��-.z g���[oo�xG,19ⴍpO����
��ťA`z��[���l�o�"��̛|���4�;+�`M��L(��/��6o� �	��q�v(�lX��s_tД-����BIS���O�[��0��Sʮ������p��e?�?e�odp~�<V'N�M�H�tE>Ȼ����̰��j���'#�)`4���B�1%=e�c��LCģ-C��R�j.ma�[�֨�>iD��n��~���w��L��4��|+nˎ��)-�X�n�����h��k�cظ���#�%��n�Z`��8�,�U��thK�������W_���o�v��;�y��a��=���u�{�(b��Y�0x)/���j:��e|��7UF��!�3���~�G�:�qQ�}�f]�zV����[?�u�c����	�
oK��x��u��:���<3Ly�we�T8"��Y%��t�K��^�>~��
�%�+��ğڱ�>�o��ʞ��'>x'�E�[�_��gE�������x�΂K����x�qA��N��x4U�(�y�[V~���0i���J7ɹ����7�fj#��b����o=-y��&�ټ@����n��j7�2�A;�~��D��U	$	�!�+Sg�b[�wt��8pٮ�e;�y���B��5,㫯�:�{��v�K���4�+6�z*�������O7������h���j�߬#F����f?
v�4�KIO?��Y?$=����)�}�f�q8
�y��kV��������v�u�8T|��5���Or�b�e�=Kc(h͘Vڿ0=�غuk����?�Ч?4t��w��DK�2��m(�G��Ο��kֹ��O�v�Q�sy���l4��A:�2�7�/0��5U����偯�}��V��qS'�2��u�LE�Ľ���/}�}V����ꗽ�x�7����=Q�$�����H�U4��\L�wi��7�m;/ǀr)Zv��q퓚�#�.}Cs��7��÷^�N����<����?���Nx�����Y���T�U4�c;�y�5�kr���vj�v�Wttvvvdvr>�L�3�/RCg��0��]%.�d���Ō��.�c�9V{i�/~�&�BQ��9�����Qa���3tM���$��P�]�fx�B���L�d�p�[�X%Y�Tf������(�V��Pl�>}z�=�(���2��)p�iӆl�����Ʋ3�rb�RY59#��u�ւ��a��T�u���^):�N�,C��#ũ,�Ƣ��Ż�����x�x�Y�F�E�R�T
��,�my�;)9�KG��t @cL��s˖[�V�T��bO'�j W��si�E��=Y�(�&�[M{TK����Sa2���H�<�ɳ�X��=�Og+C�3-�4��$�D�4�WYf��ߦE��}���8��*��,3��Ӱj��ץ��r>Mv���ٽ���ܵ���8�3�}V/|)�V�����c����X��P�bqxdՒ2�e�P�?yg���W��iӑ���I��N�ʠՕr���;�
���w��-A_y��X*��~x�?-d�o���g���TJ|�����?����w
_�}&�g��2]U�����#�Q��䉲fL�嘲p�VY��յ���m�����?��,���[pW8^�#��(�)nI3���;�\�Hq�|4�	�����>�e�c��Pn�+W�u:��$�0��>v��_Ck��+�ܿs����6�ah�VIЫ��Mo㪓a��KK۹����ַđ�VH�f{��X�Q�x����9ۼ�'ܩ���7��������T���̺��9���s����f����Ά}2�ؐa@�����N9�l�D�ͨ���&6�_r�َkޑ��tg>�0��x�T�ű�/�<�=91Ҝ���X[�����̩Ņ���'���_>������<�G���?ş�S�Nl������ɻ�#b�Nt@�."/�`Vd�mf�P���5��r���������Y�ZҘ1����8N� #^FG�G�p����陉٫����?���W\��gZ͟"A�ʠ̖�:t蚿�˿���g��r�ۙ�NB�<����矿�l�y��/NXCID�ot������֭�����x%�������~���N������͓�S=1�{{�^�Z&N�+O�В�iʷ�۹��1[dG�o�:Å�љF�U((o1+�鷼P�~ҁV�ͪ@��|h�1{�4,\`�Qf}�k�_3�Sٚ�uQ��'H�u||��(��|5���2��ۉ�0	-�)�yn���C����I�����]�<�Ņ�uN��9��m
��tO۶l�Y�	�nM�������hSv��#fO�W;ڻK�zA��w�,	2s�٢.q�9�9qd����i��x�Hz���U���Ґ	��0�~��Ǽ2?�w���\JT��䙧�^��d�i~��_N�*.��|Ky��*�a~k�0���᧋˚g����5�ͯY~rgS⩻�{�6F�R�r�����AG�C8��(��0��ϴK��$�/����R掮|�<����-0S�.)�υ9� �;�1e���m����A�h��&�����l�Y�i�<��8��Ð<Ѳ�ɑ}�1��R��ά�����棇N���>�1à�{��m�%��oݖ��g'�����7l�䩡�cǎ��&�9ݒ;(��� Mu*l�vf7y����C�ˋ\+� ��|�ȟV�7���(��$��a��g���/�x�%8a�IO��e�<�2+�.�����|W��aC<�������7y)υ1�}t�I�6��2^�{�g�_+}a=���?�-�@�N�W~��Ο	�8�6���7Nr����w�_�J|��"��$�����Sf��+�qy��>�a�i����F?�^q��Gׂ7���8)��߸�W�q�)�4�b;��D˺�3ӦS8��si-�� �1�_u�UO���!�(��A��e�U�*��Io�*5��Ne�B@VX.�UTQ����u��B?©�tLD c��N����G��Zt���XZ��c�v���+ߚ��NtϦOfc�P2�l���.<e�r����K܍s򻇛?9y4�PɎ;�={�p^���=ɀ�139�0��/�袧�����I�7��~�cA9cv��=/n����Vdƀ�.+�.^;0��۴�ap�����<�����?��N�J�LX���R�QǢ�T�ӹ|Ǎ��Ҹ&'�8��z�7/���5=��W�e��%�;?����k���A��:OXTV�9:[b>���0k��V5px�����뮻����Ӎ~.����_769v����O��b}���R�P�)Q,�vf��Ogj����uòc�H�N�:N�F�+�Tq��C����2�f�T�U����|T���46�ޤP�B�t�}e�e�+P����	��o��w1SC5Cap�Wg� x$��,3rh�D;�!-3[Hn�l�F3�V��L.��?�RrA�y���ț�z�eC�"��N��R��7t�ʡ�Lfx��odX�M����)L��)�P��AÓC�Q�>�b~���h'�s	���� @@���|�\P�IYI��A�<�t��
c��bT���f���.]����Ka����o5t��Ι摦���V��`�e�e�'�(7+���$9(k��_��"'6���(���8�W�jE�@vЎ�1���'ő����x����
=��� ��2H�i�r�d551�V�Y�8�k�pR�-r���)�m,�ο쮻�r%O����ټ$�pY.�+�@�)�O�`k=����6�`)��N��Y�e�/�)~崠��-#:�>ʳ��JC�n�0�T��?�R~&%��JC�J#<�#��<-�F���~Рoxr�Kq�;���ޭ���4�n�o��	kMs�I;�ߧt��'ϕ�ď�~�į@�Ot+��~G��Gq}�Lcr�3�K���m�����Ne-f������*;��~�i�j�.�ƢIq�s��#��N�q ����I�;�������<̙D�Ī[���$�7�qe~e=�1e�c�*]TT*a���1ttD�I���i8�U�/������DhX���ߴ9�_����z;z۬��?4*ӣ�ّ�fG86�i�ƾ=�kjf9����q2�l���Ћ�:
'���=�gX67���~v�ϴPeB~�4�i���@)h�2>��x\���tj����,a��������Zf�>��DeI�?��*�3�BiB�<�����o���K/���%~~��C9v�\j;{���}�N���n g��y?g�"X2��ر����\�[y*G;�}>�d�ڏ�w7Fܟ�l��ê�艣7��N|rh��M(p�{�:
k�\t�dm��^ag4"�-<�g�0?��g�o�C�Q�Տ�FݴNYfw�YT�_�W|<a� ��1E�4�~<`���:���"�%��(��=�:���oe��\>xj(x��^��P¨jN�O��m:Cُt���T�33;��ɻsOu�B`�����4`t�ů|��m;��4��2��8	���Kq@�:"�3K�GZ!߆+�b"����E�0|H+�;�㣟��K�0X�͸�_\�y$��d�\��a�4`G�cI���$�&�o�T|4�e:�����q@F^��8sI��y�ު0D5�\V�a�F��LU�?���ɇa�9���&~y��h$�e%Ҫ��9�İ�^�ŋ"�L���`r҂�0�X�ϐV��$K�Y��0#����V�F�8F���h?-6��+�bzS~q�z�C~r��*�X^���8m���2�AK��3^�o�$=��p����2�5�	�A�,��D�4��WfV�p��)q���̚q�~�Fq.d(��]�ՐD�gh�x#�|"mޯt�ӟ���g�~������@#�D�7O�?�d�w��wԙ���O�~�zK�~�ǵ�l�NX�_�&�)y�0���ʃ~Eq.h��7nB���D�
�O�a�~D��m0U<?�]��+c������h���}�l�l��11 �?��,�}��c���&Pwk��M�z�倏�~��#<�Zu���H���B��t=���*�֘�ei�B��<�epVD+�n1�iE�U���68��A����Hl���$N�QgƁ}�cVj���ǟ���?�ia�5�\e���\,9Ϩi���t�Q,���+�\w�u�0@�w��-t��R���(�����(��$�� ���j4�����56��e\=��c�Xo'�/�j((:����(m	�Q�QT�z�[n��7�k� ��U�������M'ѥr����2T�/�X�*����U\UU
d�h׃��1����3��(�0:1q���ȇO�<u����&��q��\ű�vf�	���0�����h�;y��I0<ykz��<�V��m�g��;d� ��T�!Z�܌�ƌ�qHs��O%�٤�zOt��Y�Ufb�ZQ��1p
�$�k����qb4'�����5��ʇ�_�q�&�%�$`�q
@g��V��TP�c����r���5e^�
z���*6�y������N��E�gf�(�_K�n�5Qg��B�	�#RΕ��X���&�Ө敏NY�(��V�.�+eL���.�S�E�̓P���:��D��������J���:g�L����5��+��<;��3��G�E�1d�yyR�����4���b$�g�G�+�6���1/Z�!N�F���;p���<Wn6����Ɲx�e�4��a����@F�O�^��+˺�½��\�L�"KIO��2�w�}w�]V,����D��=Z�ej��x�<�d�'��oe�]�Y��~��oyNx�pa�OTN?yް��ӕ0��w�#�U��.qWx�u�K���F�XG�ҿ�'�4��jMt�>Cy�gx�o�Ze���1����Ua�;�5����e�����@���M<yOrO�H�u�py��Zd���)/��_xq���|��0��L�M�~��Z�-ߑ� (���Q�h���T�i��J�B��͌�~Ұ�؎�;�m�O�3͉�=��֟R�N_�dd��*��[����/���F���{S�N��@�ꬌ�/Ub�hH	��d�P<��f�c�0�hg���T�F����fb1cS�,'����?߿o_�Gɟ{����C��`<�R6�1�\&�l���yn��[s�6���O0q�������y�7�|�9/��yd���n���t�����m������ހ�}�Ν;��_#5���?��'�'Q�o��R�8�Y��O�E�ν4�(X�({��;�2�7զQ�׎�tG�������n{��/����%������`��Qk�ʽW�X�a�l�1�2�c�{��w2c���~ڎ9ҵgϞ+���>>8x��ё��.԰r��uB%^"�W������	��D'm8�1� Oª.���E��� =QNT\Uڥ��ϥ�e*��]�'�lɓ(�Y˜{�<~��,�}k<���gP���&)��p�(����c\Л]z�e̐x���K�0��u!���Y�u���?�]t�Ët`����=aq�\� �g���V�ά-ğ��Sӭb�1�\RG����t�U���|�g�Tf.E�\D�e��z��/2U���O�ٺ�l�m��[%��3��%|ٌ��"~ayBY1oS^y��|��:~[�qV�#�]H���Y1ۢg^�tB��L@'���K쭊����Ұ
8ˡ����w�/�5g�L�DP�ĕ�g�L��WV~+����#.ý�����<j��L�G�<!kq�~�pi5W�E�G�+fq9"�c��8���ly�@C�y���gX8G8����Wƌ~���},�\���C��4KyV>�Oچs=#�x�Lǅ���s��`-3-�ߕ̔#O�/a�]�Ť�̬S��9�W��V^}��HX���'��?�|Ż�Cx�pH�W�L����]���ޚ��T>�o�o�}��*fp�m�[����e1 �����rH�x/玲,H����N��g��L_�٠�;��|�)_yM�ϖr�2�)]%\E��_�M�I��wU�'a���p��Q��'��c|��,�xB�����P������y����<���?���ǳ��'�W߫x�$�+m\!�v:����]����
���he����)h�Ur64�O ?p�@t��L9
��'�����TYޗ���K�&>߳wOs���|��e_M��|hd�c���G�=-�މ�������v_|�E�
�Q��������hK����^��<O�X�l��mGilvÈ��(J;_x�����_���/b9���\��1S���;���������{�`�����ի3k=�ؒ,�G����m�1�!�!7�?$MB߮�1uoU��?u�����+������nBB�c�0f2`F�A�$K�l��s��9zտ�����c� ���%���ֳ�i�����5�-�:U��iӦ�,�u��׻;��oE@'�#���l`���|F��B�+_�՛��S�/j=؞��$�ȹ�N�<L]��[�򖟠�c֗�D��a�K�9x�v�z+�ΐ��iY�u�({�HTj�&�!�^�S��ɮ(�\�{�ߎ���9ƴ�\��/>��3���0?d<���H���eK��v�lL�fc���͓/���8��v|�dd�Q�l��:����Nؑ-iR=�a��:�|)�����]��������%��ԹR]�[xG/ԓq�D'E}(��ݼCCI���!Oq�s��1<=hV�4uŌ�n�+~e�q2�8�ul���r����(�p^�6�v�r�Y}N�3��RGC�#�)e! ֌��^J��H(����a�T���������&��G,�O����i��Uެ��'ғ7a�5�z�,��bbdg]��o�DȜ5Kl�BF�>�NC�c0��E�uUql����~�zH���q��T�J���1�Ś��G��GѵW�1Ŧ:Z'p�����~w�;����$|�X����e�;��Y��z�r(������2�K���<c�>�j���2�Y]�{ꇼ_�[�\��h�NT�	@�#vJ���a�Q�s�cu�ϕwQ���g�cz�%.��;Y��+���Y)���`�x2�����%��O�'\��m��L}8[<sh͢/ފۼ������7�TҒ��������o��L��Ǥ�i��_PM;'���S�z��W�3(^`ܠ������Hj�8�G�{���)ڊ��[��Q���[g�s���A}ӧ?��:(��h����Kc�KW^�|���__3���|#�ip�v�NSI`�h�ѱe�
/��Ӭ�:5sk�Â�z�>�3Ƿd:Z�Gvs`��I���s����LM�β�Ew����?�۞~�-�<��s�~����M�>h���)_�j��Nl���8����X��Z�=8�;0�F���o����|�4�tЉ����FЯ���k�l�b����馛�-t����� ����{��}�s��Q]��I�@e	v�����:�SLYј|�G�a��S�O��~��/�?�~A�r���_��J����7�6�X�=Y���+늼ʜ��^���`�&������L�!�U�]�I�a��::a�B���xVDX�s	��g���:*&c��1u����5ϑ�G�l^�)!��l?	�qx<E���������;��c��������)G:s7U`V��a�C�;mC����6B��t��a&#�Ve�·��#�2}%�b�h�+oե��:o�` �Ѷ<�ѵ���j�;�������Ƴ�Ҫq�\q����L��L#Oh�L���`)?A�%�U��g�5�8-��(G�ԗ�[�L'Ց#e���1һ�s���?W�_e�M��j=�&���`�6񜩒��e����S���9%��4�ܼ�9��z��]�qSFn*#���O�~��LNs�M�5�����|t����U8��"��2����t�Wƹb���3R���HtE�&޺"^���̵k� ~幄�ݬs�I�g���E��<��>�,/�fWŦ�	T���^8����'��6����*�T������mc�O[#@��>JS���,�Z��7]��#�>z�l���*��>u$�8��:�ʳ8��-e�4x�N
`ޖ/�f=��Yy
}����^���L�J��6N��I��x��W�[8����R��M��k:�'B��|w;j�{7k���B�/��7p9�f���r���q���Y�aÆ/��>L���A��0��3��Y�\�q���X]L�4���G�����9#��1�4r5�l�y�y!c(�"ǈ���_g�g�t��Y0�P�u�/��3t�P�:®P4�ē���^��+��r�ۿ|�����5�Y/�|�?�bza��T5�h�������R��sh���(�+�rm�::���/Goټ��IgQt�st9�����י��ō7:��9/L�.:�>�0B���/�8�>R��O�dg�]C##u��8Ú6�Y9=ӺkY�0��Iv����ߧ�d��JO�l�2L9^̔ՏQ�/��]�n]�k�6��<yi�g��]�����`y+qI�Ȼ�u����.p���o��y�/n/�(^���|i��$�TMNx��$t��ӽ&3�O\��K/���(#IG���������1
5���#�||`?����kNGM|��/_�#�}1#��Eс�ئm�,:QЌs�n��{��z0�%yW�>�庴�S~e�A�����)F��}w�)����"���]��p	N��<�U����<�'-��e��O���"˨�y��(�A��L'��o{�\N���R�n����NF?�lP��4��,Z�!���X��ir��XO�a�u�g�š��!�<�WvԌ��z�<R����t�疃|�;0�d�鴟���q�� N��Ap	#oG������eK���)s������wn��&y�~<�z۶m����-4��g��|1\�%`)����iㄩ���q�,*aj��yԧ������wk�?_z�W��Z`^B��g#OYT��I��#}��]B���n�[7�ݲ-�"q�f�m�~��#����*N�����o��g��|'���~�sH��mu&����B/mw�Q��q��|�x�$�8I��>�P��_����E��o�g~�*��<��;Y�Q��v��
�)�] :b;L�1#��G֯_�(�ۧ�r��h2���������ڹ�#��L�Z�ѲX㔆�~��f�T�����Q���q6���̈L}э���ӳ���ד�p20giu���mxi��x�o~�����g�]w��,yzѩ�S��_} ڭ�N�H/R�"�@�V�w0*�E�e���T�E��h�-vDX�D�Ky� �6Ε��H�G�t���Ǿr�7�x~�r�ڟG]��S��ԭ8�����F�5/����v$ԉ�`[_;?��O�j��C����w���|��ލ_�Ty��b ���vv �p��w
C9��c6��K��j�0��|��(vx��#��WK��pm��å�8�j}�ِ>q���j�i>'��|C:%9=��!� /[k�l�� &��-Lᛀ� k�.�f-����H`���;=�i�ǜ o�ȏ�[��V�X���v��)߶�2�>��T6��S��t�+�q��[]� .c#�2)WY�A�B&�Gb�/��`��s,MG�s �p����7��Q�,�U��{��7�̫S$϶��9*����^}4N���ѕ��(���"��B�L�dJ�S�3^�>��dL��q�"O��}��x�9�`������ {S|�B���Or��L��b�
�q��_˔�@��~]���d.��sO�NQ)������F
<N3<�9�fE�1F'���]��g�����d�M+<+g!�ӉIF�&�h�y֡����E�߹��;;���t\�1fN8ݼ}��U�{�U{WmM|5ʓ/ V��'�l�_a��}im9�.m��Ua�sI��8�9}m�/���<���ek��ӻ���wOO�3�<^�x�m�i~���>W��I�ߡ/o^�2ޫ�+ƙ��ҌĔ��='H�DF~h�\Ձ����FN�ȟ��Kz�_�o��|�Tx��Z�}�["���'uD<�>�~/^�^<^�ի�qTȸY�ϴ�ݚ��ё��Se�x+|����m���i>j�qi����6�>8���w���e�C�,���/����7S%"���y�88��+^��7n�_'�}�5.�w�i4�v�3|��������G?�1�0�aÆ��c`,e��$_�}�yѳ��������8��{xѲ�c���߆�,[:}��UW_����W���x�?\�b�ϯ`Cp��&�������w��Hã������Rd^�cIC}�w�Α+�C%�#3iP��!ćh�}��������_���bt�^F�
x�_��_�����6S�Ї�Q�|v.���W\1�T��a�`vnD�,��v���
�Ϛ�o|�#�N|�T!�xZ��7���J��O��fߙW\��m�2�zoq������b��|��"���c�����}��U�+��8����{F��(Ӑe�7���������UCS�_�Y�q�#��8�4;_�pF��.{l��~S'��.Jg�,t��S�U+9���QpNw�Q%vpc$=3e�x�䌆D�eJ����bxx0���*�Ў��y+����w6\��&4����f�x�'�@��i�b��\����\cT4z2��Ȑ�8	�1�e��-W^i�2���I��
+��kO���V�WZ���Rn�GL���u�%��5έ�=��z����̈���dӔ�x����&|��$�^�T.q#�����R��B�j�o7Ǵ��nF�?�<��b"J
�淾ZG�7�!�����/sVw��R6��;~,���t�*��#���������w�ó��Y��y;�
�#��hy,���9an|�4.�K�ߏ�V�
[�э8ԅ��d���J������
��T�񮎭?\���[�&�O��[���$N��7��=���7��K���.H�4����n�/տ�H��VV~��+OH����(L��x�[~kޒ/�U����3)��o�*����ߤ�<�O=�+�r\������%�4[���je��+�����墼�o�i�}����E�|�jl>��w
�!ڄqګq�ܼ�[d?"� ��3��Qg�sE������b�n:ŋ����[����Ҩ��^���ܣ�üxÀ,�K�9�����:fg��p���=M^���x;�3�FFGO�]�9g�F֭��b�gf��������E�����|�0�ΕQ1Bm�|�3󋔎T�tC�0ٰqXp�fs�	�I��Cl��]�@�m ��A��b��G�Z~�m/D�od@g=]�.�a}ڇ?���a4��RO����G���Ї#��Z�1��}�R��f�3����]�>ǡ˻ȓ;�o�-[V��\ǚ���2�:��7�^C�)j�V��ܳ��/�w;f��r���!_k}&��O~SW�W��v�.��tF��c��w.�ҙǵ���*t�|�6]^��ɑ��td��f�eF~�I�����v?��i�c��AfT�(ga�&h1��g0��g�V.e�ڿ�@�= ;gg-^�z���'�B��l�+��v��D[ΡvU�6lt���^�9�̇�э��W}�u��s�SW�01�x��ԕ��4��O��>: ��_z�SxJ<��N�3��p������z,qK��QF9d��:���&�~�&�6eAv�TF�q_ik2O���r[?�|�,W�k���c����|��`>����-�MT��	�8��z�#�*;�Ĺ�Y���)ʉ	�fI�iB��zN���'����'�)�����j���3gY��ݸq�2uw�ڕ�ut�G�1tRx�3�{~4R_��wS�}	s�O��a[|�V�(P���9�*x�Y�
N��4��e>�
���;^����[W�*���1O.+^&��5�!��N����#>|J��*p�K>K\�n7�O�[��$��w�sՓyZ��������Щ�[�K���K\�[��_�Y� <5��_�^b�o3��k(�$�x	���&u"�m�r��]��=(��r��c�w~��c�6�G?wv�?�A���y�J%·�Dg�sŋ��y�L4����m��5���A�#��~�tw���=���C�{����o����^B:47���y'dC
:�8U4f�Eq�!��aa�(����h�\�f�;�u?�`}�]�@�±�A_�k���=��y�4�N���cP?��l0:�px��ʔ,�uXg0b���]��ޅs���_�{F����o~s%F۫�r���ܹ�6��n���p�4#�ek���,��t�vhě\��ĥQ�1��G:~��H>��p�'=F�馩����;F���@��Ұ7?;��5���GG��)\��F����Z�������)v��t��`��!������ibKqd�Hߎ[�bll5�/ϲi�.F�f�֯w���x&Y��p#�f��F�<�џ�)`4�d1�:�m3���5R�F�
�P�Vi���5w"�;��K��W��Wn�{i��kG��?iق\��&�ƌ���Y��)�u�-K���`�[����JGi�!��g]����#B�U+Ww�-	��tQ����&����2��o�~���n7��M�J;�z�>��8��R/�&��n�b�(�f4��2wD�!�LM���RG-�����A˚�_�f�ؑ�)�y�z`]���0�p��(��8V�����.}���fO����������<G�e��Rӟ�w_R�����_`�W�����ĵ��:��S'�c�:�L���毺��L5ɇ
���愼��VN�����y�g���8�?�D5j����;q-���Vd	|_z�^Z���޹Z��w����Qqz�L�?K^�f�6�A�
��<U� �sy�8���_˻��j�eoz�s�_a*_��*mG�Q��]�X����y��-}�$q���33��C�Iv��:��7h3��n�>��Ug�s�B4�g�}�Ƅ�1:�q;e��RZ&;s��s$�9-=�gC�A��AҊU�!��Q�O��|i�l�4��ȓ�N:24n��e7������=�a��㼮�ׯ_����Ί�gF�RF�nc�ʏ|��__�RƬK��1�Е�~��l���{J� �P�Xg���%]'֩S���F�ak��q��=���rޚk�ވ��	�+�߽��K<��N�,k�U=�1���iy�ó�n'�1`�(���o�g��s4�q�6O�W�^���tҦi�[��a>�c��]�\�-.p�|�8�)n��ѳe�k}��x��V����c�M.��-v���v���u�I1n�6�����Wb�f4E�W�+W���w�1f{m���G�f��3m�}OL���΋8��ԩ8����5�(G�r��N㔩+�+�[��V��s��A*=�G�o��7�����x >�^�Ԉ�+��쳸LW���#L�Ϭ�ԹU��|:��(�uX,3+�[�ć_y��#`�,D��ݍ8�i�_������yO�V^t��QeQ^EO��R��x�0⌉��'we���M��U}�7�t��$�l���2�Q_���Iؙ`}�#V���e�<޹�w�>��ۻ���U��0���r=������G�E�=�NDӖ��.ѿ����)�TCm�����^��\�2�#��t@	�]F�ٳ|KZ;z!�9W�3Zi˳ҭ�*}uZ� �*S? �N�y�{}o��:�o�}�����0���q�ߢ��"\?�i���s���L\myV�.��P��=���[�����etc���;��2ݶ�?�/�! �ou'��/mN;5Y@u`�S뇰�x�o�.��3nP�T���J�>}�����sD��a^/�~뜫�W^��򝕣RU��n�=���\�6�]SFZ�L�X�F�=.^4nik#,.:�)�#P;7n���7��=n��7~:���
�W�X}��?ތ�܎@�Р^нSF:tn�Z�E�;8�U��+z$�U���q�����os��u��l���)��� �}���7�s���ف��_z���Ίΐbl�oӌ���������V�ҁ����Ax돴�e o;�J:��NS�Q��if�G�॓S�g��
��0��.Z�;���hF�<ch׮'�W~��rtev�z��Q���z}E`y?�p!4<�f�A��D7��^f0��u�2����A"��A5�1�P�zt�k�θ5�k�:�o�o�*>/B��[�U�� �.��֙ >�D�0�AJ���]ɏ�q'.?�P�1T�mU�D-O�78�刕eL�u�`�m��u�甉˶Ez�H���K�U�i�aM�!��$�Y�%�yI��0N<��#j��G�o�����*y�����:W1zS'�43-s�(#U��'��'I����X�V�_�o�:�����^sMg�g�>���G݄)4,che�P~�[�����Sy���Fs{�{�7�"����\��6�{~���|���'����^T޹7�#����{���z�N����%4�O�������Y��Y�L�^�<�qs���?���>����Qh���E_�w/�[<5N��S���?/��*�
/�su!Nす�Gጯ��w��<��Lﯿ��2T�m]����s���8j�S�xk�W�,�ār�� ���!��o3����?Vt*K�a^/�~k���L�/�S�O�5g����{���V�lPM��<��l�� �|�ȩ�p�};��kҶ\s�5��5B;ynz���7�NC��Ӳ����җ���>��c�Ѹ/%>��ѱ۩�����Wv��8=�m۶��?[Pcf�8y��x����}�O��O�z!:ܲe�BB�S�  @ IDAT:�Wa��'�]O�9����r�Q����R��1���b�ۑj����(djax4δ|i� �V��j !O�h�qSor7]X�J����i�4�4K=�3|'�#!�8$�A�0_�ONw����1��>|$���WZ�Q�X�c|9#�خZ�����G�ng���;�@T�b4L#Z>t�<��"�]���xxQ������ �`w�,;�1b�q/���ȓj�!:d�C+�r�;�D�ʯ��]�c|(��i��⳴�W|�W��GGu�C�����q*�N,<&^����~�����,9������OXyP����Ȍ4\�e$���ՙ�w`�R��˨���G��GC����7�p$QƩoe��Z�楲�A�Q6�˺��a�]���Տi��L���D�] �Aa
�i�Qͦ��ǩ8۝I�vj�8N7�$δ��7t���w����
����>�L�Y�2�}����1��W�z��<��0N��p�a�w����я���xjZ���s����|p�M��Ժ�W��m�ԼPme�i%]|ѿ8�k9*�'o���Y���-A���C��+�݌��g�05�����+\�m�f���'T��a�+l�Sq���{�=��-�f�_�[����Wxi�Ph���c�;�U��nP �|�y}���{x���4Ἤ󶣾o�w����^N���f[��YQl��Gr�����}���w�e�ЙH�ü^�;W/��_$�34�`z�O�߬AhH�����N��8�ޤ����U��4�����������|�馛�b��������b��=���E۶m;�����_���|�6��b�e:w٬QC/3�t
���)V�3��c�G�d���O|�ӷ�~�_ݞ���e���?��O�0f71j�ַ\�:�.k�b�Sf��˔'���ɟ�ӎ�vj��ۀ��/�u�04�����ڨ3b�)�#6�ө��M&�A���r�q%}?�WG���[��j��'��7�;{��A��zG��Z��,�����G�]�y��XC5.MFfu�����&w���hV�@1��p���t��.�k�qS�]�E|�&�}��Sȿ�CN�k<�G��h�_8�	?1<��;'�jh��~��-�E�H���P��t���I^��Z���:�8!O�T�:��s#N��r�����2~y�x��+^�����(e�]1u���2(���:���T���+᝚yj,f�G���7��i��鍳���/�у�H�Wu+��J8uoPa��u:��S�\���:~6�`D�M+��g>7��a�妛{�����o��X��}�w�Q6�Y�@t�z&P�sE��A��y7�/������X�E������
�O3�~��|�0q��{l9��)��;�`Fu�Oߡ|��m��p&]��&�B���o~�ƙ���Y�%����^��2O�C���K��O�S���Zޕߋ���oqy��6���]�5��W��%��YU~�o���<\-_��	I����T>+.�6(jz��:���V��[g�G�U�%_����i�|��Bﳸ,/q����߼��3|�rjq���~�iӦ?���>y~�#Dy��
�;WgE1� &]o� �������Z��ֲb� �^8����yvZ�h�ɉi��3�j�r�F�6�&�ʠ�,0�l,=$�a��g1�����^�gO��۷o�_��_o���~涽{�e}�{�F^c	gchf��(t��UWhH�'��{����!Ӯa�:%.ip}�uj��|���1_����1p��U�~������'����\p�+ο`�v�g�����s�� �f�9?��5��3�K~�gaɢ����'Y�"�:Ó��G���̣8<]:Y;A;>�k�E�t����:83��~al�\2Վ��v��uF����9�>Cyp`���g��q��V�� ^x�7�p,��[�����:�V����'�:��1���>�۾}wzx7X(S7����aa��Ý_qAg媕e]Sq��(93j�ʯA��qp�56��;��g�8טp�j0C!VCuΪAa�Ό��1q{�c�w��1̫Ӡ���u`Խ��JC���cN�IG������YV�7��q6�����)���q0릐�)��	4C���-FV�1��v�k�>�c�Q��ţ���C�ϳ�#���x �G���2=qh��"�{�b^y9-R�̝�|���k���oGϜ5�������غ�����U���LR6nh2�q��<���n�x�c:s�2��;��f���q��vOu�d��*zH���`]{͵�������nz{�����G�]O?�Y<&5�Y�M׋��� ����G%�X �`f���g�R��YΖ�!|0���K�ǁ���w���&���% ��^B �|�=���m��"K=��ͭ��w|�����{�#<�l�u���.�%���߭��ʧq���5�t�,Ǆ�FaЕ�y|��E�o~+֩������V&��c fV�Iߴ�.��J\_��g���a+-q
W��gӹ�������ޏ#������G�+��l���$�ߕgq��c�����퍰�y^sڲ��l�i�A�?��ng���q�� ��t�#���s�h`޹:{��L9=�W����`��IZ�t��
*9;֦c�Sd=��kj��1�Mcp��4��Mϰx�<�1��4h�qvˏ9�ȟ�韞)/{x|;�Q�9md����w��/���ܿ������Qv1�<g
#vLC�iP��ƍN�������`pNM{��� �!6�����ƨ�X7�WS��1b5�s��W�����O=�ԕ�+.�����Xc5	#1~�1�p�����N�/�T ~fJ�v���읢�h�L��|�f@.N@v�ql�o'j�َ�K����"�iF��5����;��6�m��8��X1Ț+�0;�-2��o߁tīV��_��<�:
:QL	��To1#��D��c �L�ф�����8I�u;�8���N?���f.q�4
6F���Q:5�K>�>�3�uF��`C����P�9�G��!��GʊT<�Q�Y%���W�ҩ��
o��X��o3��(B�wc��I��+u�hh������Q�p�V!_�m��a����/��h�a�;�Nq�X�������ㇺ�)��˖�/����;6��oj�z�� 3�`S����5�<��F���QH��;�W.BI��T���81
՛bc�F=b�#iR��g��Bʔ��c��O%��b�(��{��Qcʄ��s����)z�K�묶s��m��Zf�O_���&z16�U�'pS&B+��K\�/��6W[�|���4<w�B��9b�`5)�S���'Ey�Y,a���:Ll�7����Z~��|�o�?��E C��'.��_�^�Z���x��Wx�ȇw���7�)�����-y�I}����/O�_^���W��_��Wg���|m~�>p-}��m~��|�M}md����s���<���3mR�p��յ���^�C��>f��g���]�v���)F���_ �Y������^b�~#^bf����4@cD�v�(_���\e��ti\I��l>;~8E8���ś�0�1���e��wfh���׼�L9��׽Ά�71mݺ���_��׮���9v42�c��a��8Eg�&��3�/Z�^{=������~g
�_ӻ睿�)S��a�����|c��*�M4�Uܸ�ɧ��4]eX��Q@$TD`�ʫ��9F��P�FwH��t�n��tw���9FH�����_�/χ�����眖�(?g�.�oj6ԥ�t�Ix�C�K�d�h�q����#uU_95�ʺ��3��ب�n��2��b�d@����U���یFyZQ}A���������M��ϗ��%)c{���gx����59�2�ꋓ��"I�	
�t�;�)���#E�>��<cP)dl��(�7��a�z��w��i�^G����j���=��L��\��_C�>����W."^3�S�n(Y�UQ�Hn�E�x�I]f4��9�
!�V���cYϨ�m�TC^s(f	8p�q�-�ȉ���Flҕ�����&6)N�)��B_;.u�%\���A�<ޣ��Qs�w��:���J�>+0X+SkM�7��1��#�)���>M�ۚE��J
���ʽZ�P:)��1�~L|���X<O��+�+Ծ�`to��2�V9[��볽��s�ý���H�s�H��Ϻ/rp��~1�� ƦI.#�.v������ �`�ĺ�:��'I�n�n�N�$I�c'��ҫ��Jz��>������&F��ܞOb��%�%������:��MX�����b�.��n�M����G�V�P�1a�`�L�Ӛ�\T�������Uh�J[˴�d�-`�S��Qwm�U�T�͕�8vCf��F���I�Q������M�}��\�=���s�WX��7�|2�n�Ep�/m���wI.$�
>�=�Z�Ӵ�6�\�~�`��R�qU�{I����$�d���H�����+���.e��ߧ9�_�z�Q��Z�-�-+CtF`I�����7]0R��;�?䔔L����L��a�^��������=��\�������?����,��_�<DB�ٱ��A�0ΖC�Km�Ҫc���zƕK˭�Q|�T�����Q��/��|�Cv3��7YV����!�2����i�.Y$��+�7�*�����Xr}�Z���)�w��=����g�d�ХG�#1<�r��g̅�]�-����ra��?v1�;����P�]��>x����r}�e��!��e���gf����g��.m��cty��Ի�*rF����*�F���s}?�T[� ���b��M���_r9������(�cc����#ۈ!� 7#z���a�u|��o���73�a�T�\?қT�'�dB��R�OZ���hnҾ0����
r��%1�]�{�[�/Ъ�Į�`�i�k���'�����*?n�h^��&���h�eUX�����J�#�K��Tae/{�ոÏ�%����
2�}�f�=K}**��<�l��L�З��N8�����[}�h�d��K��S��v��G���t}{��*�-�>Z�F�z�Ә��x���x�:�Y�8]����3��y����u��~�$<b����}"	��:���n�OH=�W���_�}=fsɫx�;^B��s�������j�����)l���u�)n��u�?~�e��r�Y��A;�Z��/�ߴL��t�0M6�kV���I����u*��~J�)�:�C�8��f��A�nK�}#��B�NZ�w��@���V�j�i,5�ט�kBc�S��}/[�^�#��P^k�xZV��DW�=kI�ξ��Tiyٴ���N!}M'_T�~�n�ܨ�Ʋ��}�����pHR�VFQ�^,������L��#:A�U�� y�?�`[�[E�J�&\�G�_��x���.�,�&�A*�1|�|{�7AC��O�L��t~2�S�<�^����o��d�Z۬�����'λ	}�8å�+0#�CL[�۰v���R�l��R��ʳ�G�i,'x��;"��͡N���M;��u���K����ҍ�f�+��A�]��E�-j9Q���H�_�@�N�����'�q�:�}�	��������p�0S��U�L@N#���_��3r+ۥɌ����I����)x����
h� `�G�l���T����֮A��i$s��,=-�eƤE����S{��1�{X�D��~�!��_�J3n���3'�S�ݗ��Г��,��|r���'J�5�Sx��A�P������ˇ�@�a���W?5x���n�vWVv��iA='��pl(��-�6�ˏ;9�䧑�ni���!~��^�7�@pD۷�����)�g�o�����-" d`,��46����.r�i����ƫϿ�Z�h�r�3O*ar*(��0�t+�.<�e���C�����=~�� �t�~|���Ϋ�R5�ݶ����,���8`�<6�N޶�փ�P!M��1{�*z�BU�b5�`�F�w�;�i/drM�N�T�*�k��2�v�Q[u$>�gD7ۨ� ��I��R�{���e={�<g����H��r��יJl\oW����1~�������,�=WJUڤk�s��\�U�5Si_u��ea��r����ӫ�U�ޥ޴�D'�x}~�Է,j-Л�ѵ�>%X��<nfj�<��+�C���l����Z͏�VÒi�M!�'�KJ�P6�|��,-�y�*$\�]��E�s������h��P��ts�(��Ui��b+�}o�ʻR>QX�l۠����`��[rC;�c��[��(J����师 �x�Ǣ�|8���J�D�ZgC���v4.�jC��Z��J���&q�6Q>�=�	�>6�]YH��r{�=N�#��Ȳx�"�׿��dD*"��PSo�$0/�b��i4.C��7�����'�U��L�0�����x{���y���X�5�Eu�P�]������S�Ii���
H�B��{�5Ü��{�ʐ�D;�99_�=�_u��6ǋL��s���^�x����PNMz��b*g[�Ġ ��1�G��Pt�d;Ub,�1D��x����9��.�~0�kg1���у��_��;�$J��;�py.�^"u �9�wCO,��b�9�T��S��_��Yb���0�l��%�*��7��?�Dl	�RU&�G�^k�7����O��3AS<�slp���m��8�gZF0��KP�h��wϗ|"�N�D�i	���>��d�1�
�����_���ɸ�[n�<U��y)�)p\�%��1,��Dx�z:�|j2��0yg�C�щ��Q�r�w��&��
F�����83U�)����������f����u��8#����n{Ȁ�O}����p5�s��6gF۶����bD�"?��56ڼ�1���P�W?�"�M�OxYo&��͸g���+�Irzb�L'C�8��ɔ�>{eǁ��_��K3�R%"�ϧ �	�g�h���l{Fn����c�����?3��������:�*�"�q��\競�	�el��!د,��H�S��b�D�V�G�{�7ܺ��8nҔ�K��p/�6���}ܦe�:�#F����9����^���J5�ͽ ��V6���QG����n>�\�iH4C�(���d�m�m�Uc�?�*�Eb�m��a;?`r:�V���4�0�Uw�n���y���=�L�<��?�k����굲(�('��I��GmV�8�nM/���Jh�s�]����Q�p�!gr����ܸ�r'�$�￾ջI7��2�JI,V�(Qd�)��N�"�F�F�]%�DP�CF�̿�t|D�����(g�3g����<ΓK��o��2��\��M��xl���ҏ����@EyML�.79�v7�G�?��Í�< �1A�?GGYm!׋>аSk��bd	d$�;#܆�%q۹�$j#Ŕ����n���*J	�Sp��{O��
Hߡ0W #J��N�ж�ލn��)�eo�
�!�c�=[nr�hLd���I�͂;x�h�o��-c�y��	G�q1y�U�?�O�O�V�M�$����*F�l��[�S-p_z�j$M��s7�#�<\,�����))a����EG�o%IHr�,�c�s4nk��Y|:��4�rϲ<��e���n����?o��2 �-�׏,�<�K�$*w\����~#֒�1F��p/���Hn~M3�h	�W��������L'�#����D��������?�8�)\L�o�Y�d������_d�.�����]U��f`���	��b�KN-��%�=�ǽU��&ߺ�M	W�0�F袕X6w�������Ma�&�I��-�?��]~�dfÿ.���f=t��)��a�S���X��G��xp"R�9�V��8�dl,��}z��2T	��xcYy���.�'SC���Z���gY�=�Ə�YĎa�����
*{+*��b睔��tw�ڵ
��Zܖ�?�|) ѧ��U�FmB��i�e����{9^��g�j���+�h�:x����{�`Qg�рh��N���@���-�5�>fӫ��@�P�d�ޞ�ֲ�w�;�_xT�<V����ZE�G٧�"v1��f��=�QF�Olǭs,;-	��#	�����z���l^��xt�|����������H�����z�y����l0�{��Ȍv2��o�Ub�`��	jM]T�n�&f�%Zl�c;;���X�����4=�^�ո!x�0�3��f�'��P�d���٧^ܺ������4{�v h��]���]a,�D�1��l��C\���{�P׿�3����*�1SeM�T��	hT��xyҸ�a϶��Χ�ar�(���G=ۚ�0�@��oZB�����H��ۭ&�%	�[g��fiwpl�Y����V�"��<�b��k�Se�ł��A����r/�v���3�CE��?�yI���A��z!8�ļ�A��Ʉ�P	�zo�*B��x-8e��i#yM�P�g��Y>Շ[Z�[�>ٖb����{S�(GVvD����dE�R�g�x,|ٙSI�X34���X�T�$K��IiN�0
dd��l 4Ob���,֚Ǥ;�k.%�w��6A2�|�p�g|jƑ#U�l)^n��o��V��2�?朑������	�����OR� :��x합��c���$�,1��3K.�\�ڝ5�3�s���Mgt�;��������#�)���\��$���`��(?�j������z7j3���c�&���M��R�9�7�tu�a��4C~d�l8�N��'��Ge�D����3h�C��S��M���w�Ӕ��v�Y�ã�>��#���b��/����2IMb�'ڂ��=�+�p� ����ک���i9}��Q��h�c�}J�<n]rj� N��k������7��U`����褝1�!�p?͕`4�o�<ɋj?����C&a-�m���v�Nԑ|\xuM��`��[ڸ[�=>#J}�_�&8���'���������I����4���Ҿ^+7#��6v9�!+B#BP!߼������]�C�oQW���f]�'�$Ӹ)� G�S#��n�z�ã�5��HƞՐ�笏܄�D�yg�/_�x]�ыb=g�D�`7.��s2働�#�>�l��c�2�⭍�G� �L�-z�6
(:?4/���0y���u����ف�sB��w$7bhj63ohw�	OvB�E���B�g�&�����ϗ��(k����R�!�;i���X�7�l�V�S�?]y6��(�wi���a>p���>�'ka�:S ��Y��G�2>}���,\��x�&
��L�$��[�6'��LY�����'m3��|[R/�2���X'��� �_�d��޹g�iU>&KPI�-�(���h�V�W���GA���"n�7j��l�Cr.������f|���D���=h����]BGV&�Y��x\DYD(�pT����g�� �Ȗ&v����3bEMK�Lo���*�;��&-����O)�χ�||���Ԭy�l0e�0���,WYV�WEvA.d�O�x<�e��6h��Rq;ƹ��#�J9��]Vd����`�����h�[�Ҍp"��hj��)��Pv(>
�r1v��l�KZ$*�����J.yB��+����DO��|���ɛ@��7�EHJ^�S���+��g��>�c��Z�Vڗi���ٺ���s��#sՏ�*���ڈw��+b=p~���N�w����N��0nJo/��Ʈ�=�y���3����TF��J��e)ZS�t�O?�'r:�2�*����Kǃ����o+Y~�{Fol���߅Ϯ��^�)��K�Q��f�ppa�؋+��ݹ׵/�JG�%��#e�Gj'����*��y��EE�eL����Uf�G��6jx�Nqd��k	��ցp���e	.F�����6s�i��(�@�H�:IY���<0�hm>��V�9�%���l���h�F�}��3f�B���|�� J�/&��~k搎��妬fB���O�����/�0A@~4��DR+�|��Δt4J���$w0���}Cp�D���L���`���
�}q~x��Y�\���D���A$O+����:#79tj��쪢��nY�M�݀��D���?V*�v�lfx���)o|̕l���j0�`��H���(1K)�»?�����KI>p-�V�5wQ/)���d��-/��N8m�J�
:�k�$�+���Od�
�D�W�oSz�G=�o�@�'�缒`V��#֨���N��c\�h����F�����hf���~����� �����9b%�$cK.3Q�z���OIĀ =�t����yP���!���f������$��I�׃�H���-�Ҵ��m�w�D97^F�t�)Z�/�2��I�`�p�zBa&O�Ͷ�d��S_�ߟ65
s�|�Fz_�9)
�4���{����I���V�w�z5
r�3q�$������{\̬���.����Q>4h2��p�l�(�d��v"ɢ\��]�mgY�k­�8I��"u��������C�{}/�3���{!ߖ��[痥�`�&�{X����W�����D��V�z/�}�Ws�P�������4������Gz?�7�+�?d��F��$�Ho��j�V�"����q�8]�����V㾈�{�W鉒���^|�ޡ� xtX�dv榕���͋=���uR�{��J�Ѡ1���i2�g�Fb$.�3Vj��2�=�8��sI�D��w$�Hn��L���D���;j�'��]�^��p|�L��v�f��k0[�y��ն���$��O|�����<g������l�K��ɝα�u{?��̼����Ǫ�h�t��9�vwCB��5a�k����4h��'b&��\���B���Xy�r�	�v]�'�{���V���0Uܗ����^���isl9v���r�!M���b ��ܞ���en5�������=ԁjܾk��}OP#u�g��K�\=d�Qz��d��ޭ��éM��&H7�
�Ƙ&�7�n����Do�逴5tEb�_\*��G�8�#��-��+�vpI�Q�a�S��^$5����2-�_9D�i�k��)���{��l�)<+�9���R�����% \'$7;�W@1�Gz��b���{���u�`Y�jﻞ-��/ �O�c!��;�ֳ���R�������L��5����4�˘��~ `-$[A=x��ZB��m]
I��r@B�`r5V��>�.:�Ɯ�m��IA���c`��W��uM"���>)ѷr��}�A!ގ�hM���?�{ي�V AЯ-t˨����0�D?sc�rN+�<�
���c]7��W�9�p*�N����X�
���C��L�Z,�s���FD�/Z��1���Sl�C��sX|7HԲ��T(�~܏<�W��v�~V�L=���)��{��]�L�B�T��>��(�>��+����W�v^��b��{�U���D���7M"]�R�-���X��
������ ���
��O�&��Tb΀X�\�x'������8s��5����3����7��`����/� )�Xlb����
�1]$e�@�ي�����4̺
r-,��z�S^��"���>�W��������o(�b\����`��C� [��o�T��'#��#����JP/�jW�����g���%�A����9'�9�^��U��M�F��G	O3�������{��<I��}��?ݩ�?���C��K��cޟ#f�cY����hߩ�S�$7![O�s� w�]����o&X d'�ƛ��*�o2j��J���񫰶U�O�#���>�ń�S�a�^46�#�+�o�}���V2i˚(dF�="V����B����u�:�I������s���a���9:���%��o�C$����Qz��ts&C_�pM�u����Ӄ/t5��]��X���5��0��Ig_�4�Eڐ?rg�b�Zڟj^T���l:o<@��B���0�����ޥ��v�ͷ�C�(M6%����ZvR���U4A� ́�M{f�]|d�n�@gC�]��#w�gekQU�|�폟fpZ�tn�����pۼ�*�Qx������.������m��u�MU�W	)Қ�5տ
���S�/�*�p�N����8����5�XݧC��R�HZ$�����ȯ���eJ�D�7*�����̳P^.,5���{������ Є�7�4�	eD�E�C�l�7�* Dl~�2�)oi�2�a�;A�m:�6o$,�'�LKf�s��}L��w�Ųr�t16\F(��%�{�d���߾�,��j��v)50�W�!����}�˧�p2o�-��7C�͍2���R)�U��0iS,w~�6E�W�W?��.,A���̌=Mp�쬱rx���{���{�y�豕��Ւh���`���K���v=5PgG�TdL}�k�JH��[���f�VD�5�iT�T���ƴ��p����{P#�N/�A<��q�o�a<e�[�� �R�_�|�7\A�T���(_�\�:+��͏=K�?N� ��Ь-%r�9�Wzf���F1%�����%��lܸRb�	g��Cz�.��(�o�[�Kq`Md�n��O�9q�o�Hg��!�{io(1��f����4,�Y����ݚ���n��?ܑ���t�aMi�D�m�V����q	e ��Z�0�����x[:��q���n�WE�Pp4���/�.B`/��^h�8�"v��\���P�3�Ƞ�����_n��ݪ3z5.{3�J]�4'�UF�uR����Ɩ�ɔ���{@Ut*i������&!%��;9jHbQmI�������2�\"��>�>l#y�}�R�ݳ�d����L���5����@@i���A$��H�r��(6
��jH[�.mvr�`��B ����eILL�⚺��ozX�oQ�œ��t����ϼ:N�M��1C;;乴��tWyc��/Hf$A����DG�l(o�k�ʩ4c��+����'1��/LP����х�ay�G����c¢�׉	�Z&���	�k,!�|�D����ή�[b�RUr��`�揗�1P����mZ�Iji�ɬ'9�3�f�1�\D&6=l`���{���(�b��f����B��"I��Z�����3���W��_�N�9?̬�\�e���wH���;ペ�^ZO7�~� _W���+� �N����\���]���}�a����/���O
}m�︐kĴ���d#Kw��o�I�rmL�N��m)T�&�6�&�^6ٔ���z]���TӀpx&��=UQ �Q�I���~��V��d '��B$���Yx���|Rk���m{Y*���{W��*I|����;OX3UU��-5yt�hH�d�\��>l?���8������1��م�	Ӟ$g��3�16�XO����	�n>�z�c��S��g��b	n����
�Wk֪-��b�G��A�=�/�|�W�{��%�Q�	�\_��'x�K�a�]���찞Y�%#y�Q��I���AR�n���;����O����%j�b���-���E�I@֕G��YQ�yT�U���a+�_�=g�����[nIM�rT\���7�l>��T�gC��$�2���w�?_r��JF���#��ӕؘ��	��x���ٞR�D�jj6c��gľ����Yy�ah'���u�
~�.��эP�FU p`�/~/N؅5��}�E+)d'�
���e��KV~뾐�'��"�U�b�aM�/�[�g���J�ۮ"�a��lB4���\���ޖ�=g!�h��r{�I���?)jy�G98�[���ƺ�s�o�`]� ��t��.2���7�gtF��Ң����A�\��=�􆛤�"���͏���X�YG2j��'ľ-�c�ho���n�As�$�(>{�ݶ#����Y~=nR��Q�!21��Of����	���˴ʍ��p �1Ⱥ�Э1K�^�� �n�n'��Ӡ8~I3���(T��@�苜l�|+!N��5U�9$lƢ%�L{�[�^'w��1G}BB�e�_�/
ۍ���zbXI�Pr�{x����_��!��e�E� �QC�۾������H�Ī.1-x��ݥ�xϱ/��R��!��:s����.q�S��e	���7ra فy���1�4�-�_7�����V��[d�Df�7|V�C�0��Y7.ֺr'�
b�J��e7��6�i���)�̦���i|~-l��K&�>�t�8 ��c���9¦�ɾ�"���ݞ��I�t-Ej�+T{�U���߮����e��D�;D�>�|�g����S#����u�%R_��F���AYR����{���w�i��|�%�Y�36wi9�v��٪��o��e:��u]�̰�O�­�i�:YjcI�xB�8^�h3������ �*�t��G�μ|Q�����If����VB�1�Ǫȕpi��08y�uBԾ/�9~�pך�3k���2�F��a��D�ɼ�m�Y�����M�8�j�۪�_�R^8N�����Fjd�=;X،��7w�J�?��4���p�s���(�����?ܭp����.@�3��4i|DS�`��E/�HZ�a�4T���
��	���.km%\���ORg��4[qS�
i���C�F�d��`�]ē�����n���A;�ew���^\��v]|9Y$���<(���R}��<�-���Ҋ���.�}�z������8%W�ΌL>����W�Y.��/;�cx�1?F���@����[e�^�͐�K�0	������K�Xz��מLr!���سJ�"�zy��V�Y� p��U���j���LDU�@^/�&��o�s�_�W�NBZ�ٝ�7#���Z��s�LY�Cۣ~ZN����Ckx�BZldy�i�8���O"]s.ϧ-Ђ��lu|Z� �a**��u��N�7=�?�f����	��S�x��_�T��=s`E�x�O8(�SOK " ��V��Hf�����є.��ɵ�<z��vD��Vg�Il-Z��9���=-�#Y�䣓gїa'ه1o���a|ܕ�\�ۯ��ȿQ���:�'jx�Rż�kn9�[�8i	L���d��2��p�M>��M�OdGq�?�ޟRMR9��OS���[�Փ��r���%���cUL��|�H4��p��~fws,���\�����w�?,����Dn�P���2d��^I����������T����+�=�W�,�;����iH�O0+){ɺ�ImqO��ja���dƔ��N��(�`��8�_�9(������� �ѡ���Epq�����6ء�\�K-��ݔXSU>'"���)�}�Y��Q��?�./\26h��j�C#�Wt�+彝�/�7��V:�X|<����u�Q���w5�Zb��b�ZD�fY�;�af����w�]���΋dϲٖX��6{?۝�>t �<^Y�A��C���{��sq�it�֝bӭ[�-+���n֑��-S��+��Q�\���z�m�b���UǈKO����VE/3h�R!�f!�ي�Y�gY���ě}2�w\�����VR7��X��h|����;���bo����y��S��;���(J\��J ���]R~;Z3:��G�q����;j�FP�N
K.f0t��0�9��7��}��J�� �����K��Ik5a>�O�Gh���Ţ�&uD���_�C�W`;��"��-�;�FQ�{^����ndq�6�1c���.�e��ɱ����4]�$�dp�����5�sF�۰1jER��}�&Y'vSiW�a"k�w���X��Oi�$�I	��a���5���q߁B��j��vUݣf�%�,�+ڡ�G?a���Ǧ�u�p��F��e���r�u�i���� 2�:c��<X��	{������D��Zrr���¯w7+K9r������*�lN`�k-{��S�R���?��&1<��W�kII�ߟ1�ޠ{%EG�c��1�]Jz����C�T͘<��A���C*����A	}�!?fB'-��\��rt���G;B�<w�����:�K�L��1N��~G���2(f�!P0���v�L-����8j�) ���mϩ���E�_�������\�g
�I��9��gʸ�W�x�沧'a����e ���$X�H�^�������@���{�G�*o=
`���'�g��Zn;t~�����ر!���g⧊�9X�]=Zp�T:��@>B�6w����Ur���o�Y��a�w��HI���e��oؽ��MO���ۻ��L�5Y';+eP}�l.�kW��ir��܂bZ�<���i)�cVy'-��x����o�Y9�8}��u]��c�0����Y�quh��� �գ:�.��8��'eD�O>z#�	9mg���5in&%֓��ݖ6ӎ�Ɲ�׮$ �OQ�nD��dn!Kb��&'��X���g�ϊH��' ��n���G+�k�zMDK1�e�=_�ώ�~S�j�y�-�>�m=����QZ�q�h���ֽ����z�׃Y�\�[*�IX�k��/�9���6R��3�)����z<�U�|l�W����և�l���$ "��.UM<S,����uB��dgy3df6�WjfzXx9���F3�w�������-7��}��8�?
�t�d��ȡ��q~&/���=��2���'X�%�3	���#11��x���`(M��<��M?�\��{>�loֺ��q��l�%��͟��NA�����h�)���ZY����j��汰�=���d~�0�V��J�"����H�p��6Ci�SE��u�!�'r@xד\�ET|A��zk֞�Eq` D�q�(�(�(�A"Ʈ�Y^��z6�� �'-���gn=ΦF��?�o���o�S�� ��̏�Ιr�6
���>�E�R�	)t�3]"[t��>�d{5t�@�.~�O�ś��#��_+{�O��=�D M2Q�P�W��nɝzt~�V�F$�z��5���>�[<s1nR���ʪ�c~,�P�����_T�b�k���'Z��qG�!�RO(ɿ�;y��j�C1�>���5��g��x���gU�'�ߐWO�Kv�q���׌GE����,H5� 5���َe�b���k��bJElվBT��R=h�����"h俘2���\��D¦O��*R��k�/�j�r�'�����p3��]�j�D���
3�������iǽ^^ѠWb����i#S�_ҧi��)P�/ma6����W�QFSqW?6�yyK����{c�p�E>�3�ee��������O�3��>5�^e:���ƪ[ʖ�?��8�!3:��e{�_��[��ޠz����B�wŜ-a�vb��|�]J|	���:T�����ؓ$�.1�~�;!}��VI��"���\����@3_��j��tJ�A��1��B���7�2�$��+�+��?߬��g�<�%�jp���p���;V'�����<�<��) s�2�?ُx�O�	�A�}s(��Ucj���fx�	��ID �ĄO#�t]���	�� w8�I�W)(�րL��ֳ԰`1n_^��t8+<U�pQ�γeڹ���6�8�)6zr\Q鞽`ȿ����U�$Em7(%2\�n�_hX5�j�b�,Vi���2��Ϥ���eP� .j�QW5�<�O9����~{a�Gz��A�+尕��{���6� �I�?���6{C�o�"���1�/]�bz��#��A�#�Ƨ�	侌'��n�U����ڍ4$���G\Y�F�wU���n�>��σ)�ϴ���zጠ�`@�9�k��?��I�ȱ�-=~b��'�%�3 5��j��XhY����<�C��/\mC"�2�` (���o�N�-��Y��ѩ��,�*�4���NҎ@�D�㬂X\ ��|�W�ƩҸ�˳!�ޝ�����ֳ�k4��)��C�οMB���7H)Jow�����?{�-Xf�`xAm�=�:�:MԝT���鵶$)
2�]C���f�q6�1�ەp*	�ѷ�Ԙ9
�\QDWy�@�!�yy;U=ͣD����L�7�4ޟ*O�|>c;��&d�V������c�ϡ��#ǋQ����3�f��܋!U�b���Ձ'ۦ?*���pz1�O�U~��@�]�Va��j0�!R�n��R��\�=_�2�=ŝ။a���x0��c�D�p��%@��LC�=S����iܽ��_n#s$��/цʽ�߱,��^'�a'�q�ӓ30�x ƌ��B����J>QV��A�g�K��>CS[����ݬ��d�B*�p���*3ʕp:�����'EJ%f��$���G��*+�u�k$���#^A�[�~r5�c���4�'��3N�c��h�ݨ����v���o�ʯW*J�o�O1�;�s�:c'��e|�\X�ઇr�=�9�"�>��58��W�����=� G�?�Q?��Z��g6���f 8G�L��#���x��ߖ����Ee���C~��6���1۩&�&�_�|m�u'8$��ٯ�U�2^~�2��.�k���xFc��_���ꪌ/��^|�囂�����Cl�!&�p'�%����Z��Z���6@jq)Z��F��L�݉ڦ�����<�^v��'�l�rYwك f`��&��?�7�n(�x�����I�ө6;�)��\l8Ǳ���f\ք<ǳ���W?������r��8%�f;M�v0�倘5�:��]᷽'t��<�{�,��5���Gf����1�Y�L�h�h���َRM�l��T��k�$�uJnf����7�H����;Hͦ�p�V���o ��-�\��G��{���Kq���FTN7��J���)*3!�PBqd�$�\~�GH0�F8�gn�=�a�k��+6u�i�,�w$H!� P���Y���];\_�X�ǫC�L��̫~��y�d�/߰o�� �s�b�U���ӟ)yG��RMR�U�ע�N�{�_�d�B��l��j�`�=ւ0�60"���Jy�"��U\f�S�����??_�alE�U��\-�.!TމbW�9��
��Qǫ3�աy�,����j!������O��ok��֖��%=nVgO(�vV?���d���:TaV�F��쵥$k
��I��j���2�m֮.���ψ�<yC�����9�FZ:�8���9�ם��Oq��}�݉���F�����{H��о:����|;����߷�9s���ܜ�9ͩ>NB+�V$�pǮ��\2���GB}�o�V2��T����b]���<�|�f-s�k&�#|�{���ģV�=tIkR l���<��z��3�Sn�=�ސ�2�_;����T��©,�0����3M�[e��?�p��'��0����7�	Õ�C��K��s�"�Tf�B>ڄBj%�V�&a��Ixe��%��Tֳ��k�EǶu�=N����eujmRr#"���>@Nj3������M�/���Ǟ�{}����!պ,JW#>MU�KR��OW��E�Zh����&z8X����)1�_2��1�nd�u�N�g������^3:�X�Qf��2��Xh�]z�or��6v4l�9_�U��0�8)�ӕ���F��2�{���CDg�-R�3�	Q^��S�N\����J�MK���v�]]��'���[Y��G�Rn'�+�Ѭ3�ђ�NXZf�,�,�ѿ�WG������/�DD��9}�cmJ�dj�jX�9�V����F�<WDU[Q5��\1�܆����M����8�~���x��AU7�6.�'��ڵ�6m�EtQT���X�\g�)��_t����>0�P���Ȣ����򈹧�W�>F���cL�^'��O''�R��7��=bFb�վ���n��,·Sb����c�N�N�̪�x�9�OX�-�R63��̇S՘ u�xN�b�;A���Y�ՙ�������8���ak!ۅ#��E+�g��%��V��H�擑� ԣ@�HӞ���d�,8�q�&���h8�p6���۪V[����%6���j�5j�X��-m�.Ak��;vm�XAĎĎ������~w��9�뾎;WA��+��̱s�3;�2�&7�
[z ��W��#�!]N)'����ݡ�V�@��鮓R ]��I�59�(#���c��P·{���S(f�8ɢA�ϚL����gt�I���2G���{�Ɛ�S�Թ��M�S��)U�TJ:o�t"�]O ;����e�ȝb/��0T�9z�C�ZF�W�P��N���7��d[b���Qzhg*�� �aFz1�Uڌc�
�P��y�b�	X��إ���"3�j�}��TI2C�sOU۩S�S:��6zus�R%���񷖚��B��y7�U?���O���e��ڼj['���R��l���Pm�5v�-O�$�ї{�h_��6��X�d��Kk8��|^��`�B	у�l��x���$`}�ǘU�r����?�~e�?��O��BsFn'�k{�=�Z�W?�V��v�5��]s��L��k`��%UE��ɍ��s�v%=�T��(�g�U�w��a�/���hzc�[���g�R��t0���Æ)��y@�����8�vWAZƽ�K!L2<\d!�U4��f<)�{�ƩhO${ȸ�A�B�"�/�n� �ئ	Vy[����:��
�S�ޖ����	m9�#�}��9��M+��}�iO��>l�xT�+*��{C�6����)�v����}�Br��u�;F��������}�S^0Q���օ��N��������l`e;���.�J{���k���u�/�K������l#�)6F;w]#�F�������Ӽ\�����.t���_%T��Trdb�_*����v��3*d^�̚׷���#��.�,�̴8��`�y���h��ß^�I]��f/=��"��?��F��Z>1fP�Cɹp_4b��&T1"�!��������&��F6w`��t@r��"9η�����?���=:G����5NLI`IJ{O���y�ʬ�f�eHy���^��-I^���k�r_��?]=Co:;&�6pB�|��a_!��t�R&d;�8S�抖�����V�O�A#��!�YYj�e]�'�0�$+9��M�=�X�4s�*�뒛}	bϛ��~��u��+���1�<���=_{�G[d������kA��#I�������)�Q#6�cR�ް�Յq��$9��$Ĩ���%�sC�Ӻt��s��x��F�"��w��7\	F��J未� ;�kIC��`�DV:��,P�"r����F�Z{Y�m�7��;>��i�w����'g���F������C���	��o<���'�[��u���>mg_|�ԛ^]�	��Uk�<4�!�&f�n�2'���4������o���})Gа'0)ݮK(��3��{��`y�F�,32��#F�{C,��3��2dr�Y�13�V�����P��Kf���G�z ��a��Q���ebW8'2b��_��5>�O>��A�W����ޱ:��z�>�9(����8Ռke��g��H��_��Gl���y���?H�[������l&oe�A!X����2۰$d��%��N��U֙F���<�f�z�]�m��B��+\�ON����M�~�Q5X`݂vTC�{`�K������q�=�)�����eQG�ws���i�#�*)I�v����t����
���3��6�LfB���<]�\"��w�k��;_���[BZ���9���{�;��m����C\�R�0T�GjKuɠ:�-�ܡNk}�<ܓ��u����^]d,yH;7a#�*Z	s
I���������o��έ��>�5�t閵&����$\��GƲO����?��p� �fF���}1����OG�����Um��'C^�6�
~�;�j1�#�r�)~�2c����:A[)��U /(n�Z$���]��l�J�ϷE6��t����B*yq�Q��p�q���ߴ��S}���`Hfn>�z�K���3Gy��q������d�# <���	2P����F��!�m�y���\�����t���(�8��4���K�WCt�#��#�J���@v:�̥*���Y����u�	�TmKr�%��o����k�\&�Kꭈл-�ڤv=���p���/l���ѹ���~l\�sدe��Q>_��;)�w�"s�{5���lD���J:�����D��[����y+�rv͊�r�?$^�7���̱-b��:a��1�ĸ��J�M�����`�)�hp[XS���� �/���Q`��V��*�y1�T��ΒyZ6��1�/:�u]u�Y}���:S֦Z�*s�Κe3(�u��w�ulWZܚ�Z�U&�"� .1n��dZ�(���D�� �l�O����`�h�ځ�m[���F
�O�2^����-���U�
������>Q�_ϊ��oWlx$ky���:����6&��rw����q�h���IJ�������{��I�Y�,��˛�8ޭKkQff%����.����2�����w�67�6qd��:�Z��!����%���@*��݇D�7w	5����:7�d��=��<�C�)G�OЍ��_QE�uk+�&����
���Xg�y���ݍ�z�J��a/��֦��;�p\�ۃ{$����|k0e�4�/$uJ�,�٭vΗ�
�1�%7�r�w۴��ˮ�X�\:�rn�ԇxt���h�pW�j΢�+���>�Y���j����k/�b5�3�J� G@�^�a>��&)k��k:�aF�Mo��	 ���}^�Q�z{���ֿ�=q�KB4���t]��z���ӫ��'�Z�T�����Y��5�@�cI�B�7�\Z�6��X*p,'HD�^��e׬���9
�0�*wO�*�f��C$�ε:��/@J+�Oތ�15�5l�lv��r��v��7ޒֲ� l�w�\�9�����u��W5��pu�h8�TUyL��������t�"��=�譿|G��վ�yЈ/s�ݳ�T���\'���( ��0~�Ur|^�����_$�rוǄN�'1:1ބ��
;x7�
���Ƞk+�_�=.�8�*ɖDA,u��bͩ��7m-�,y��Կ5�d�}��
�[:�b˚��W�5�U���yLoQ��{�g�^�7ˌĞ�\��ٳ�`�Oֵ��	&�X���PH�<���1�j`�ƚ�������	�'�bi�m��~�]z���u�Sm�Ͷc�r��I#%�{q9 �O�7��*�E�H��0ؼ֘��3Ʉ;=����x�=-�W�U}��0]��1���ꑘ?�J��òZǣv�W��r��; f�9�&FR7M�z�Gě
��FpjV(����cD;����C�uF'"�]���M)��Q�t���4d^������'�+Y��!�,���L���'�2�W���0��0S��ʎg���z�U�w�:}�r[]B�âS�c��<.�tX̬��:�J���Pu&H6IIm�a�߇GnY�����Iۀ�D����Fy���2e7r�o���*��)�3f�هsO�؀�RXkPq"��,��mE�>���i0�q��LR��AL�Ǣo�To�h��i�N�u����s:����b�Q@�����oY�|,?�og4��8~���HƼ���%LW��(6.��O��q*��\�lpr�i>�.�҆�p�Ң�8�o����,u��Ś���u�e�p�8j��R��c�A��{��!���-=_����VX{	��Z���x0��'�����/��hF��k$�,�!�}g�� zD�� `.��!w�����A1�D�1!ҋ_)B�F��~~ZmZ����l��4fl�t�ҳ�W�1wk�/X2W�b�����Ͱ-��_w_=uw������6*�A�RYG�\8�����L�[q)���t󉌘�il��;���՘�[� ����m|��¦��#�ֳ�G���='�m*	ס��*��v��F0ڸO���"M?��g��%^&��T����9j���ny:��8��x;#o׫2�7��T�N3��מ���뽔��h�A�r�J�iv��FH"�=���ݙ�<KܔRb�7@/b��n�3FTZ�9�eMQdNGI^��� �a�Y����;�����y��m���8���x��:�\�b��͸e�dvK��@:(ި��m�6�	�{>3i�Y,�5:�'k�jЛ�\�����i\�(��y���o���ܩ+���3�imo8�׀�cd@yu%E��߸��pk�)2O���{8���{���19Q�Y���0tKӓ�k�k@*���ɴqpԉ'�c�9?D��h��~v�$�p��T�l�Z���ޛKX�u�W�;��<�GNtl/��N<��p&�Xޞ2�XSsbv`�p�-dv>���I؉�<�?X9��E	�k$�}�ѭ�ޠ�+x�#	;_��,��,���FW�Ѽ
/�-��í���o�x�ǒ>��$�ҋF�zcm\-��eF>y�j"R�0�3�攷�ogv�ik��^{�f0Ijg�m���߃��@�5�A�43�˔��h|��-�I�j�R�awI3��w%=�"�m�<�ѷF�˕T]�3mFd����(�?��N�bn��^�Q7��+�����n��uڹ3��G��n}
�x�~��0��S���梤V�K�:X��Nf
 ������w>9�� �;�Lv�7�/��8	���|��ܨ��-���oh����~iy��˱�&2F�.�-G"�K:��r���^䴠���u��%��;�h�s$~3 l,2�!k&����S�zL�+[<���B�iss�'Y�)NG�b
E��V�߾�?�rlp���,��r����Ύ� ]�]�$s,o����R�įp$�V6٪`M`��=��������>DnT{��.���#��|R眷_w�S�i���8�R{�De���V�N ����y���~�NG?����#��"�O�Bkp�U�}3��`��zż������������13ïGwԉ"�v�h���*��w�r��/U�kW��!,�c�<*����f��n��>
?#��({WXo�b��FdHW��%>��bt�^i	����#���"G����7R=m.x�i�4���?�ʹ?���8����o⪻�����:���ڋ7�ɖ�wK��j���|�Z��C�cUd�����%���rY��m��z-���D߼%����?[���s�*��bɦ���)7V�C�O��9��<�p�/�ݎ���B���Pp�/����ݏ��� ��Z�e����W[4��w���fR�Q#~,����#�&^S�%<��5��E��V,iT�շ�>�In�.��Ϣ�N<��r�Tq�TI~mf�@/2�HM��������r���z'n�M�J*��U&iZ�c�2?���~G�J�J�����㾐+%��\N��&��&�rV-�{\͞��7���5�vC����yĥls����a��UƠh��/�=8�\��?�H|��`�@Ȫ��.Å�S.Oj��L�ܕ�Ò�z���y��Y���_<"�6�#�BN����^4���b�����d3.���a�U]��A�~h�)�#�R N����/O6۴I��	E�ke*g���R&�aMc��B\��f�$�?��q"�l�`+��m�L`=��D�~w��˰�FY��5��F�(>.������X�u�?���#�?�HC%=�{��p/��(��0{B[�˳���v��b�Q(B����6��9�E�*�߁���sV��Tg�tw�O��t�'˰=�O���=T��#DYB0:��E@�᭑V�]�y(o�~cv>��<p�6"�N�)�x��#ؗ�
���a�}|�d�gN�����
^q��X�ob~^�x:�oMA�&i2�z��`�'W5����F6����6t�T��W�m_��L�l��M�u�*����/4���N�<���X��ca�Ϡ#�&b�O��A#t�2�`�4tu�7Ŋ�~e���K��O`lnJU|�4æ��[����d�\o�0���Ij�BP�Yuj�ϰ.~uf�����o����u]�!���%m_�Rk�D��L��߃�q$Ɖ�_�_�OH
^�SL����y�]j�GN�ԗs�(�>6mNi�Y"�f@��O�� ��ik�gs���1�~8�Z�̚� }ĳ������6�Ek�����@?j|�`�m|�@�fRu�_�1K.d�a�?o����ߔ&�H\K�����a���&��hק��,k�z.�%��1i���֙�e�E�d��Q�)��C%̀���[i��2$�p����x�����|��hc��U^
����8���z#��H���K(uD��ո�C���ʐE*W���5:�=̓�������A����?2���h Oֻ��a�(
Y��Y ����Z"�]��1)Eu+�wJ���)Ұ�?�jx��P���C���Ef�Bv�Kb9����5H���΢L�jJ��/���P���N�"?ڽu����
�	��\؟&�Ka�:�C4Jj�kYZ��HG�yK���ǧ�rl�v��a�����8kBs���l�&%B�zl��@%�R8M��|~8;�d|Ȗ�Ż���L��0�L��� ��\4�U-2Q?[B�; {h(UH-nm���w�b,T^���Fmf�FRn��M4��wl�~�����߁��Q;�#��EBj~c��W�˱�:���M<�Ś�k�EZ;�{w��<���PעA��4%+�@�MDIU�� f�?F�k��PN��k���a�(�6B�~",Ϲ�����y�:���t��\X}�g'v��Nz׋־B���)E�����y}���{}�����0l�6 �X,�q�
�V)̋�U���De�Y5`ӱ�e�9���d�3mBi�K�0�1T���~1l�Y�!$W���5�r�Mn��"�~������ǚ�3s�����`^��}�4�m̾��UnF�^�AMYk�pvm3sV�&Wk"��w3%�s����3�s��W!���o�9tD[���x����!6����r�����MB�
!C;l����ו�#:���
�������	A����Ԅ��#���f��H�>��M��
%��[�w�*�F0��eՌUs���^wضf��xDFO�+?^ږ����p�@Ȅ�;��4StN��EnpٯK9ͺ�ˑ/��\B��}0�[/G�{��s`���T�!3�<��x� �3�ڀ�0|�g����K���?�ic����o�(�3f��U�`�P��r��'�V��|`�e�t�Y�P\�]Qy.�Li�`)�7���b���ahX�c&ar�Sz$W�?�,��{�A]TԴ�[G���Ѣ�ˉ�!"�^��Q�L���Y'��Fw�',x0��f2�m;�_�|��t},K�^�S
��[�G�&��ڡ2��� �w.��P��P[-4ݟ9�EK% N4k ���KL0��x�\���5L�����,Ho��{;jx?w�:�Gb�m��[`õ�[���뵼٬	�"Tڢ�7��ݫ��N�ʭ��$f7?)��*_y�}�#�kc�5�tY�o���Y_[��g�
f˟�"";XTG���h�,��t���v7*o�a6a�H��i~�,B$�5�˽
L���X�֝Q;����<�lm�M��p�-8B��]K��� =���V���jM�}��rj�3�hw}��6d�0�֦�����s��m���D�B�)�4�$�A��|t�@ʝ�C�r������&�V�~:WM{ւ��LCU�	��
�ؔ�BX�Ӱ������}�0���w�Fm��Fэ1��}��"�2e�(�&--W��4��P�V$�7��t:�PD骶UK��U×˟S�\fp,H�
�s�$��b/zǬ__2�u�? T�͹�L�F�n7��n8}��,��U�����\�;��o�3�/�KI�jw2�\���5���������Cx���V��4��9�$.)/�YlP½�I���fܖ�V���U?�݊���ҍ9�8�)"��
��9f�ͥf�/ �A?�8BT��G�������uS��)����Y�M�Ry���soY{g{xZ,��"Y9ّ+������e�E}�s�V�-���°\��RFhM��Vb_������P9�B}���z�OZ>���|s�$��b�Lґ�T(l�OS]'jH,��ss�>�K+=�C��Y�`�q�w�1˂Z��|0����æ�w�=��q�$�U�m�60߳?�U��${���?D{͘ȅ|6I>k���-GZ��f"ĕ�@�}�j����הr��/���F\xttqì�p�9�v�w���$G�)��8�O��p>>���A�I�Y�F]�D1 �aSՔgLuo��4i.<*N�������m���*���o+q8�y �������Ϗhk%:�U^��V�Ki3Hfp���e��G��B�}��
� |��˝#;�|,:����0_O\���{/1�ܩ� ؅�%+Q�Q��P�����:aj���
�/��+k.,��w���#�������3�<�޴xX��Z����9(]V~�BJ �������(xÁ,���b�e ���~�H~[���}~Z��G�C����:B/����5?�nQ(�gJX-�]krK���p��m��"G�� �eo��/t�gs���q���܇�rc�%1�o�9ҭtH�й�mx��S��ӹ�(��`��BM��XS�����p,��9C�d��V|�ӎ۲�I�g�k@��)��g�n�?��Oڋ���"H�qុ��
���Jad���^5K刵'|Gt%�1�!��8�a��c��l|���z����d�KY���T�W?�+�ݴcG��c�G����[�w�d�+�5��C %D.{�UÛ���[��#�L�d-���v���`�\�ӛ^G�_����߻��"K�\/O������X����R[W�[�iڛ)%�N� ږTժnab^w�ΰ��\}���Y��^��/t������-W'�vb�R�aOP�s�y�n�A.�"~3wF�hAr�p\_�ֻ���A�<
A'�Y��N���F�Y����_u�y�I4$cV�e��wA�=�Ϗ��v�?3u��Ώh�>:-o�kV�hZ��j"�u�5��-hsΏ��߅ڌx���إ,Y	��$(Z��E��Ц�ɳMƁ[���D;R?E������xȇ$Fw���U�AP8�ܕJx�-5g�]g�I/�G���!���F�B�G_���Rj&�����2��M^m_�zU��WU�d[h�s�?��H/���yťm/X��~'Q�֐�v.�o���Qg�����W��r��[�o�C�wgP���Zd%ǰ>�y�[2=�^��+���x�S�8ՋP o�gP���7�b��OK+{?e������)����X1�Z�Q��M."b�[�n�56�zWG������_3���$c��5�ҳYՔ���O;�����,�U��s�^M��ߘf���87U�?�V������8h�c�����H᱊�-sj�F��Y�D����í_������k��h��(5�õ��e:�zz<�.r�>���R�SzP�ꞻ>��崦��
"��%}W���~YB��:B�Y�6ݏ����l�y��$��[�c��~��.I/��0Od�Iɪ��|���z��u��ز���c�'Os��$�Jr��_����	�n�4$Z��\0�z��ג����}��s���Wl����~5�xr�/Y;�_w3I^1�$��c��̲ݜ���Z�ϕ�@�3�r�1�]5�m;ٙ��8�@G5�kOL�����(砸 �g���q����C�k���Y��Q�.Z���!+ʲ^0�\�/�F�N�(yɹ@���0~���qM�1�~$?�htɯ���q�������Q<����6��H�����"}3�ɣ	�(�:��`�����K=��B[p��a�g�c�3Cf���Xv� s��c��]�&+d����ש��wJ�.ڲ[6.��y�r��g�C/g��U���;5%��:[��e��Y���FF�X2M�s�G��W�����GN��lg�O%�,��ݘXL�)����*��#�\�$�粿2WA��/w�wޢ�	ytƧ���=���&�6�#���{3*F\��@7�co*:�_�أ��'l}���j����2�8�L� �m#N�{l��\�6ۂ�-IL��&��'����PS%+^Fo���2 �SP�-z����x��\��}Sx������̃����1�����Ǳ�|m�몯ޓ��7�����f�j��J��~(��f����)&��p\;p����r���KS�֥���!�x{i컐Dț_��ٗ��y"1RbO���s�G�_�Y��E�v�EM���l�D�>/	Ր&Ge�-�I��^�hCϱ��gwp{��T���.7KD�)��buǷ��\�1���������$������ju�]�3I���N 3��@���l_g<ӛ��*���߿�bޓ���{��`:���
">�0����Jo���D���$��o֠�NFQ�T�11t�n.z'{�P1W/6*��$��5�T���љ�;c�ׯ \q��������_;o�㿊D�U�4����m��F�]&����_�Z���5N)�s�V'E!P�b���?Y�i���=
��a���K![
x����~��0~��O�*��ƫAEf�eL��.x���P�DRŹ��O�
�q*,:���=��űb�+3���� �Q���G�;��7GĈ���gm���.s��%Ot=$���{Bk�zR������]���I�������):D晨-yW"B��M�7UD�Q.6���V��P`��.B���(��k� ��������� F���nb������4��L��z�2�O�l#�Z�z�i���E��<�e�T�;=.����n_H����;,��l��HAzj�ں�&�O�Uxe���ea��NI�@�uN� �"�@�t|O��y*2��q���Ĥ"Q�0sA�w��?�C�%Eܞ�jv���V�2�V^^!aا`\��'�>0þ��Uf6�̌2k�Dj�������ם.->�,�/��7�0mS�vƖY����g����Q���y�Go�ѭ�R�+؝�Z[~�1�y@S<
���p�O��W��R�Sɥ8F߮γ8ph{Vj����!��*VR���K.�Ԥ��J��p��nY�Mt�_���h!r���onZ?��H�%�I<k�.�j��-`L9�:������
teo����T<6ߎ2U[]@E&q�����4�8�o�d�V�O�>�H!w����Ŝ˾�Ѻ�MKTJ��Z�@�U7Υ(�"ʈ�����Yc��ӘJ�$Q�
���p�&�y���Ο��$l��9�c3��<��ٗ'
�9�w��#���n�Y+nt!+�T���j�*�,Z)�.��IDgXK1��g8����e�O���8�շ5��P��5���k���UO:De�J�g��$��?"���3�!Q��^��5����\�U��%A�)���R�\�F-�eԃ�j�� b=��=S���8���`�@�����~;Qa�,������!̬���&xd\�cE*+#Դ_LU_�f_L6�dd�{(��Yb�e_�E�r������tN��y��'4���K+[x.ﷃO��`�}�������+
����U��i Σ�*�s�0��"]+8~ɹ���2�,^\PB�QCO��R��Tx��pKq�u]H�3���D���\-M�m��#�=��):p��eq�4�9���,,�~xmi�r3�Q3xk�
r)4����\I�Zll�� 9���)�w9	:s�W���V@�AQ}5Nʕv�3�����i�?S(q4\�d��/m@�0�9-�����)����l�|V����'-�4�� ��^���i1��g`e����+����蝜r<)��9i
A��"�a�I	;]j�M���_Iaf�C�$s#�;kSP�!������L�Y^��l'@�E�il��l���F� �;։�Wڬ���[q��RՓ�8�r�O�b���*yI���<������p}V�I[��Hu_���u�W���b�#�"Ȫ�~IxzN��3��E��W��I�dӝt%n���Kv|�dܱq�n��x���'5�_.��w)��U5����zπ������x��)���WA��M���I;cۣ�W1�}ߛ��R`�J�!@��s�rHʢ흛����b3:��s�٧�Һ�a�r���b҉i��}����R�K91��E��]�e���#�!{�e�,]���+cO�_e>�_����sx�<G����_ �?D��M���F��v�6H3*�����8��e�_�o3�`��򭴗65�!�+�w�#r�/%!��L�Y���֖��W�އ�f�X8�=�W�3�LҜn���N���O�ȗC��U���C�X���}�������u����a.��K�KCJ-��uơ����)�wbk��:M���,Qjﮢ�O�H8.�C,�ZM<�MT}�*\��aaq"���b�B��dK���0R��$$x�g��%_�r�θ�s�Dv!d�r���ŗ���ø���
�e�D�����������Ώ�y��3$����To����(�pV��5B��tQ�o�ڛ�7
�J3��~W����VE�=:zC"m�,]��g�?1��*+�k��s��1�����B(���G��7�l��M��iԏ���xߝag��m�|��xȗJ<�$�0I�Rc�1h��GN���5!.D�-��>��)�;��+RA#��l�L1#c�{��ٲ�5�O� (|�6��ص�b��|��<ʪFD��c�c9�f��y��EQXLQ7n��"
6�8��Ռ.�=*�����Ԝ/*&�m^\ku����������.&1��}:�:�V �g�IS5���98$I��[aO�9yoo��|�����<�Jʾ��̰sB��L��n
��_T�I���9���\�q�Vt�Ql��_� �2n9E�U�,~�͟)��!j#f�?��熔�k�I������ps�g;8������%z��`�#�9� ;��N�t�_=%���<V	i��ƻ;�;x�Zt�I!˹�l�t*ɔo�X��`�2���U�RE5���ZCӟ0�xyٌ��xK/�^���<w�`�$nd�8�-0���[ZL�~b��H�����N�~ܠ��.jj�����|֨g:UI�Q�3��J��+xg^�C�5��:�|�6��`R���J+G��c7w����R@0�q���y�82��:gʼ���sG[Ӥn��'E!�9/c��?PK2�N�L������mo�tj�*W�ֱ���}�B,~d� �M�3=x^2'?�Z~�^��4,h��Z�'���k�}]a�K�g�e��\y�z�K��ō�� �oc�Ǭ]��y���oVِv$�.�{����9:2fq�홖�����=�K]e�������.n(ݜg�].�g��.�A�bv��װe	���d�oux9l�	��]�Y��o=�F�nqIQ��036��H��ٽ,����U�FK~7�m>�C1����+�.i�a��[���<�h(�X.i:B�1$H�IY ����z���>u=��M&�n��;�N�Ԙ�5Ʒ�����j�I�6�_ �$�.��3]Z�B]���D���q��_�1=��
�e�F���wo�,9)���9&����;���XRtl9���sʬ��4*��d�iD������aݸ&Ua�3�D�������9_�}���G2J䜊ai����P���c�Y��J\���:�z�����N������Fk��J�c��B��鼩�OM���g����@G���j�a-�ݹ���9k��b�R��RF:�^�����9u��%�#r2�t3_�Hw�[�M>��g�j@N��P���Rْ(�ͽ���JV>t���t�I�z��P��A
JY�ջ.x�<��0�z�,�ș�̸��x�	9�د�\���WҐ*�3aZ��D3����C�;n,1rIU�O�rh�c�>d:U�Vt������`-�ģ:�E-��(ǲr׫@ݷ'zg
_ڬ�L�\��~����.�y���+�]���K۳��`�s����訍���Wo)5L���+.s;`
��bՖ�M�*��C>U.%�%�m0�Q�IQ��}�����i
��]R���o� ��jZ��f�aWO����Ww.'���1Fh���H%ϣ!�� �҅���!`�U���t�i� �Jɗ������V��:����R�~^?�D_�ꙫ� ��]��<��;��Mq���j�;hb�5 xY�U��x��Ñ������,��6�J!��q����RK�C�G�^e������L�pD@��+��ubl���� �~��lC0��-�˩G�;z�3�)1����1*dr�O�;��y����nL	��~�C�d��	��\�丨��t��ۇ�� az)�2F�F�'���ƸE�*�����*;r�c���j�����a�Ȱ@��X��]�P�����#�v��.1+�;Q$�$-���	���+}������XE���-������������_��?��h������,�diu"�,>�3%zQ#�vM�q{�73����;���_����������gT���H�����?�Jζ!ٹ&1CT���F�Xp���r���*�?l�����lt��W�*������	�kjQpGϜ�-,w�d�eg<հ���i���)�
��{���+�[r9]��k�i=���n�y�p�m>dZ�fY��{��g�	������=j��uÇ@���<Co��\U;���@�Ol=���G_/4>|ގ"�֟��<����9˘$Y����*�?�'�����4��V�h7�x9���R:��AP>���/�s��J����l~
vg�L�vNJ7���4;^�C싫:*����{����~����
�џ{�\���)��6Kp���?���S���&+,i�c�H4��K��ժk45M�{�Y�q9�VQe�q���	���w���w���3;&���]q�	�'�:-�Q��9��ǀg��
� ��xe��/��j���P�X��)�cE�оo��̓�g�[�$'����H�ų����~>}ɜaI��;1��I,���ao��`�����T��	~YC,(�|���6SU�Ψ�t(�����a;U����숇���R[,{��1�����ԋ�$��op
��,�}���i��LA5t+�s�I�X�c�#_-[):�5�k�ӧ��1�]J�?��W���|I��"���7o�²��h����e��G@>����Nx=�������M�(G�|���p�����O�)�7^p?)�ֿ��'3��Q겒-|I,��� H��:O�����3T?�8w�.�Ϫʼ:�l�3c%�W��3NC���:� ��QWf��l�AT�y�����e��XT��y�禐P�w��X`�礉�����I�(y�@�	�:3�R�6��<�DA)�!����,p��I%[�+���`���:��t�ZdH;��axç%���](B�t׀Vl�k���u:Z�]����'������`�J�V3G����0� ����v�H���"����b�n��_�����AX4�&2䵎�|���7�Π���(��<�OQ�܇1Q~@�<���0~ה;y�y����#��O/�Rq���j�����ed�;�jޥ~����60@�"S%h ��k�D}i��I�޶t![��w'�@�k{?���R�@��gZI_���<�[��,��|�Y�5R��7s��9�L�dx.�e�v-~��YA��!n�1���e����.���3��]P�A*��jN�U�O}�Q���
���2T:�N�h��dz �+
�G���y��NM8~��G��@˨bY=1d�H�}�:K�x�j
�HٙNDT�<��%}s�̌��v�d�t�e�3xv�%��d��1��b��:�֙2�U�b�Ն_Ʋf?�v꿝"�%n�J�-c�j�0�b=l�o��B�>R���4�v�&�=���2E.�o5��#c3�S�����뜇�NM��&�[*)�צhf��,����T�Z��!sp���P�"sF���׮��p�:9U����MA��li�8�c��$�B�&���(��X�_Ď�ݝ�&)oK.�LS�f��;�8���LT50h>�=ʳ�L�	+m3��h����VDK�-�J̀��Rkn梯ް�H��g[^�$�.�����l0��FK�j�Vk�UTmQ#��5jՖ"�jｪ�6��VK[[�-�&b��b�����������{ν>���P<J��Ew�֪H�b�1M��2R�)<�bݢ�{1g9�T��v���X�5<��e���C�����4�A�`���	r�Za�Ya�nۨ��]j�R+��_����O6@&�uɶSGcR�[ݼ��.|u�A�#XI�u�<����ߢL�M"Fm�R�ې��E����X��{}��?��p��}���&^:����e��z/vچ��a�w|y�����X&�nW���2�'d�=5j��[�VƓ�ʿ��l�+�
 5�#���U;��,>�󞭧�YV����� G��6����{*o��vr`3����	����Ǎ/��6,�Eș�^�m(�-\Hg���A3X�\�)t�	O8��>�'�=����KYGFǍ '8 T����)Dc�"���ꉣvIĽq�XZ��&��*��o{H\R�w�R5��HhPk	u��j%֐��n]+��b/�\����J/�` o��ol�=cD�k~	��� F'�F��y�+��}fV��+��Cm��7dX�F��ڬW{�MB���V;�����fR~L0`
�X�*�#+��&q��V��ΪOQ��ʂW�瀖Һ����>'5�f�V��������ܵo�ۙ����:��B� y�,�W)���fU�سۯ��;^%:ۏ�mK_�^˴�,ϡk�Սvm�{۴g˰VY"�����`�νJd���\���{䌔mA�ƖG�Yl�2��T�5z���������w���8ˏM���K��zR&��B�����RJG�N(��=��B�Ǵ�rN�Q<J_e��Oܒ��뤖��QĠp�XX�_n��NhDt��������RN���崙 �əuE��\�_�Y/2�x}�Dݷ1?�G�6콷��?Bl����Ŕ�cov�!\�is/�����p +߁��5��coo8�@�����|A*�*H D!Rܿ��U�U.2�[��9�CcP��oc=̈߶��Y����.1HaƓCW�j�b��I��>"Z�>�i�%<����<��+�� cz>ŋ��ʦZ�^�He�l�9�v���F�ꦿEk��$���W-/� lG=X-}J������jT5�Y8��Mw�wU;�-���h��45 ćR�i���M���Z`7�l�x+s�s!���*M�K6D�D�[z�7�w�U��A.��Ɇrw�vf{i|��&�/�B���2=U+����a����˳�d�j#H����8�+rKxͶU6kzs�jCd����/�<IV����z#Hh�^�rM�����{�D>��V�V����\�d��W�'�m��`�����.0׼��5��o��i��d5��r��s�S��4�Xds�彶��Y'�`?z�.���䧔�����{J�ҤM�x-����qo��d�}#�8Cc��W(N����9V�~6t�:oT��S��gh�\�~K9�;��y�KW����]I���Й9�Dӛ^iە����&w�a`z��T�9�hǹZ��*i�ɝ_�:�(_�m|��Q��1,�at�d&�9�̬��n�총�GƇR&�z KL�қ��,�O�X@���BD��o�����Y9��>��U���j����C�iDs��}�9�#������vAJh:N�Z.5T�r��(�����+�p��f�DV��p/�p
�fQNMqg0�v���c����_<\hP�y��g�LDW��,�l�Rp��1V(�:�nH��fu��p$R�YW֎�J�c0^����{ڲ�
�ɤ��5B����1�&!����>U΋�-�]�<c���ʕ��Ю��K`��Gj�ox���Ĉxj3�1�_�?�hK���H%ܘ)s&�S�t�l�!���<��#9eF��������}F�8_�rr����p���� ���'�c"��{��`�ܝ6�:�C]�o|+�4Y-�?hM�[։�-Yу\x�������*~��zx�pb���� ���'5zcbU8�-������_'�e7������)&���I��O��U���^+�1܀�+*
Ä�0�\Sf���H�Rj���L=��W��'2�>ڼsC�>��H<��~w�s����K��Ϛ�zZ��W�;��y���{W��U�L^�X���{S�2d�,µP���{{#�T䚱2۞]�"��|�w�)�:!�8۴Ha�6w�;� P����!\=z1H���if~Q�t�r3��z���ɆZp����^ ��X�gZm3H?Kz��QEdv��,�Y��ƍ�p�g��;�^_ܩ��L�����&^����q�Dz;��xb�A�⾫y���ڳ�T��d�"i0� ����&ȒLaE�I���+C�!gqxb� Rg��S�6�~Ϸ�{]�\n({��
���NM����?q%tBȖ�4�l*GwL�)'��1�c��R�3t��Y�!r��C�	I�@��2d*��O���sD����e��(�b��#���ƴq�%^�-k��swn��w�!W�̬��/�����$ѥ5����J::]yN��,�U�����z!2��A.A���m﷙���^t+x,�"3�6n�:��P��;'�L��bz��'B_4����2�v[+�ʣI�Z1�v�C׭�h�x�拌���Qb/�q*�S�����!O����!B��`�O�e���4���tw+̬IT,�d��[��N;��[M�/���X"Gz��Z�d��+8U���Զ�a�Z�xjf]#���g�BAU%�O~�#G�4g��P��J;�z�	GN';���m�\��gp�m��!rsx���<1�H�w��_��ׅ�v�nN�XJ���$Z�K�+���G,�^�K��KSBT3S�����K�*�_��{nHs�y�)��]H2}��[�ݾ���[�a�{�3ϗ�t�|��k�j0���ۀ�-j���\I ��@��-����[kb�L�Z+��۫А��ţ�УZ����ҹ���U:��P��'�KY��s�ۆW*��K��;�0"ak�~������B�c���ٱÙRl�W 9����`�R�n�jq�L�p	x}�5ǘ����}�ձ�O��>���D�if�`#`C���w6^l�X_{2���ճ%�����Lh쩼kc%7�q�(ݍZ��Z���<��%<&��%���ۗ2xQ*�J��J�ƃ�!��E��o>k��7"G$Uoл��X�x�Ѡ,�5��HZ���#t��m�^}.�\������:8%&~�*ݗ�+v�)���q\Pr��x����Q[R��ny���7]���N��MU��B��Y͡a��z��4�y'�#���fv���������l��T;��vM����H�4��n�Y<zvI��)ϣ�;SD'k�+�F\�� �H_2#��
W+k84q;�B�6ʝBK�n$�_��P��L8�=x	3v�'A��[�"��M*�e Qq,��ݴ,�����h�9iG�z�	�O����,2��o��	�	��*Ո%A�Ԥ�3h��d�]zN�"��Z�_W�NG쳘$�Ñ�z9J!E��nj+ِ�W�+��nT\��[�fF�z���I��\�Ǘ��G���(�-������{p�m8XuP�!ysD��s*|8ZMY�R��+P(�$���;��Z����J�.1��_��`k��R���v7��F* GZUG��l������l���,�\�콐�/-��=���l�zY��èF��K�(&o��s!�KA�֮]$��"��k���T����L]]X��n"�,��B$�->/��{;Sx9Y��B1FC7�G�����^�s���#�J�m��ɢ͚��������5	N:"k�Ի��6U��9�!9�$�"�/֠P�~ʾ��j�{�9�r�J�v��4�t�t�Wᠬ�b��M��E�$
)��p���P���%�o34=��u��b�Ӊ��o��VP��o��W��e7�<fyQ�Td	���	}�U8�rӞk:f悒W9���	^�jaɭ���_�W��zȁ�aMV<Mdg��,%�������V�э��rmJ��~@L��y�1����x��܋!�݃�ao���P�ߵ��g%t�%�-����gs���i��D�&W����Tx��t-����7�s���2;H��Ρ�z�Jn��Ouwf)��h���>����7��E��U\i0����E��B�:w�m�fN�:���`����r8�*r�Z���I�����S���]��	'�A�	��cgNC�Ww�xڐv�8�ހ73�`Z�+�3d�Tc����bV�����Ķ@�ٱ��xl��>��<u�xo臁F�]���ƘlJ��_*c�~�5o�.�� VM�8��J]p�����ҋ������j��T��b���dY�稹^&�fb�&["�Li��v���v�HL�<Ϙ�8-H#68dm<s#�N)����<?(s�e�2(��?�#y�L�H�(w;��\Z�װ�|y�b�{tW�- p½���PT8�C\ϝ�ژ�j�JQ�R0
��SLЉw�tϙ�3��s&�|�ŀ[ʐ�L�6v�=�������|yP\-�\��bA}L3n�F}}?�}]��:أ9�ːX�H�4�on{�[�a;�Нo��m{qN3�.�@�0���/�m;���7�-��q�4���l<�����3�xb�`�d���x$�
�������ތ���� �4�<�~v�,�#{.�N��\e��X��Z��y$�0�]�K�,*��o!�"�Ұ*l	������E�D�ha4���м)1�[%���_�ѿ:��g�P����ٔ�\FL� �LT��'1_������J�mr�\�=$W���,
��,�}Q�@��E6�uscI��-��y5�~���t��I�\)���&%��_N�Cl�F���wJ��zv�����m�SjU}����ȷ �DM�z1ǿ�����vC4Y�t/�5�^�)�n���+,l��|��l6�jv����KG���hOĒ$�f�"CC,v&�/s%%~�S�(|gyH뮣�u�F:z`?"��ہ�.��o���~r� ��ºږ�D�ˊ�{�N�}�Kߛ5�� R�fZ�Ν-J5/G�%�׍(����fK8><Ť���X��*/!oC�C��#<=_|�U��Y��Hv;�'���y�J/O�.�
��G\	�u��藩��w��E�e���㗦4�ւ���@���߁�����9c�~�#QO�����S�˩�m_0�G|K��<���, D�\�}��[c��g��`��o"�rI�"��%�|0ecr���D���0p��}�؛��l��7o��ڴ����xZ��Pr��SL	>�K��bw����r����R�}��ГS������ ����i<խ�%A(����2?=:����� ��Ǘ��ť�	�k�%7���E�/��ǖO���#w�5���=�k+>�0��P�}e7A�ug�>l���yEhF�s�|��x��v�_��z���x�p)��ňl�/@Pn���p�+S�����kd�I�m�{�4r��Ն <i��xs�"9G0ۚA�b����"��h�' ��2\Z��;ח��?f�Ǐ9�]q�~�>'�i���_]l����e+O�j�0=}V�|!d�.���i~>|�V��~�9q�؅�I�>��X�I�.g/��4ߟv�UЈ�&ca����-m׏�B)C6U�p���f��ud����C��-,�w+|'a��*�����Ś	uIuryb�P$��w�6�9��������7�m�#s/��~|��e����E����Ev���=5�F�G�N��B��*���P�L��J��yNo�:�ЂM��!�dp:,��6�v�]�0Pu���͌���_��(��uve�<P\G��|�������)��M?z��yw�>B�g��tN/9�/��=BV�3(�5WLz�R,;�y#��X��"�"6�*�v���M5}!�ߑ�X�+� �v�c�FYX�Q��z@D�L������ ܳ����'%����!s�$)�q�Mt��
��l�����I�L�u��1�A�C���\�-��r�1������R{\'�u;�k�:��YM
~��O���8�o|�s����Z�v,\A]1t`�v�Iy���Ī�5��Wa/�����FT��}�RE�DZI��i�Θ�Wv3�
&
�>�!��W���	!���ve'�����ݲJu ! �0E"�&�Z�q��{F~K�Z����?L���7��Đ"���т��%h��Y��_�Wa˨rmC���%;3PuF"�zJbV|�a[뙆���<��^a�]�RagR�ũ2�ϡ�ю6a�f.N�?�)v�K�^a�
��>��8���Q������R����?��:N��쳂gK�M�l�G�:B7,��E���#!���f���2mѥ9Jҿ���I��ɿ�#FO^�I�^�o{�W"����
��x��ae`w�#�B%�7�������$��9�C���_����o8~ �b8���f��M���Ki?���W��N.��Z�� �_�B:��O�Tt�Ԅu�Uc�맾���
Q��&U�Oq(��
OC%�v�ITs���/\�����/^�0
}j��n��HuZNEe�˳�4�'�YLs�WݓRb�=��|�������}�K�^~���U�k<
3rQR#0ϩ� Jz��]yw����I�v�Q� #�>��|����d���A����AF�H�m8ƍ}�|�/%{0?Ʊ�C�sI/����~� �����rO<�z���+Sٶ�xD��FD���t��Mff}��h4�;��G����	��
��\�J}���X�#�<�<7�{Q[�5�!T@s��6��	q7t_���Q������+�c��5&�\x	V�	2��>�L�H�L�$e�4G����EW3x��)�K��D�ȗn�6����Q`�Ӷѓ'�"m=B2���@t���m�H�^�FYa��LOu��l��0�ib^��4�[pZ�0���2�$ӿ��د�5���'�1��ǈ���li�z �v�T[wq��.]H3ʾ�ޗ���[K��ȭ�y�~���sߜ	^�W&����V!6l�;������������IGV��m�}l�{M�,�^�at`�욣�K��A��p�E����DYH˲P�v�7��,���
�X�}���^������"Y���5���A��d�/Ke�)c�T�����<vQSQw�_�`�qW��� _��q�e�d;�C�K��}�?����Ys����&�~��j���0�].�����~�lw��(��M�r��	Z�0�9\+��d�4�齺�g��
�o��"Rբ�s�▅[��;SO��$_e�X�����Ѥ��Ȧ��U��&{��ԕ���{]rXE$���͚��o�}\nl�;~W��䀓��:�j�V�u�À�x�a.�ݠ��~���>;�I��Յ0�e�yL�g����K7�0R�r����G��� ���N�N5�
���t�N�\�l�ҍ:��h�
UU��Zt|U5^$���9N6m�픁;��<ந��n��N����\�K)���'41��X(M�m�V�h`�5,����Q�X���.��x�ӯ8��> ��K�R���|��pN��/.�;NMP��I4P%��IU��VJ~�g&Vk�����%~QY\l0�	"�OӞ���U�K��x6w��ˢ=j�e��Z|�6��C��x'��J��%�6��`Q�\d���߈L��ΠK������>SF�"�@"$ͅ��r@�h������/�z/���6?��>4��	���l�œ�$g|j�-3��T��x0m�����l�ٻ��JDw*n��а�[����S���J�5�� ���oe�I�F�Y�H���t�4��:ES0����\5��>!�?��"���:��F+Q (E�?I���NK�/����x�#=Ӿ�V3�(���I-8���93<��&M	Zfy�S��$������}M@�
Z��u%�3����pe��,�,*�,߼����8C7�O������٘ LP��yF46��)�U ��0u����4V6�e��"��Zm����*��P�"-d�a���:*\�h����M!!����:�C�9!��������S�C�t3*�.ju���֓BM.cmM�*h%�����ʟ8�x33,o�K�8��.��ᤢ�XЁ��7����8
=��������>\�I���K��<d�}���n���׉�L��E>�~e �ɖ���j�����q�9�)B{�]�~��|���穉kf�e�b�*A((C��#�2�m MҨ0tR�׀�ʠ��y�hl��`�dʐ�����U?��:�ʻ��Յ��]R=%֙��S3$�-v�\�On��sf]Ι�g�d=}_(�m�l�⫪
��|�]%��~�7At��h��y¾N��X����mX�k����Wߩ���og43� �dK��Ԏ*��Am��%��=v���N�4X������A�8���8��q�1���0g��)�D���Rфd�@O�
��2����';3a9WTK� c��s��N�>��`m,w6��\���Uؙ�e`�S:�|/~�ȧ�=�<��vF��62�����-� ��Y�y��}(�	�g�� ���l�{��&w���Y`��~=~0�X�����JdD����hb�ΐ)�V��A>+���72�����Cl
��#9W�2/�ԅ_9z���2�OL���5���`\P�QÎ>g=��4���==�$��1k~d�).�)�����'�t��Z�A�u�F6m��Tx�)�<bZ�W	e@%�~��;0�M�L�J�Z�%�4S�業v���+-�RV
��h����>����xXZ� �F]����{���f�J& �/؊Y�d��$n^ p�kM���vT���!"\<�x1�L]��b�t�J�>5Ե�������k 填���!�6���hì�Ć���red�����'��2u��߯�g(?����1ŗ�
��.f�������.Cx�z*�d��x�0V�x��X����m��G�;����)o�'k�$���j�Z^��+�.	Z�U���AI����d��5���!��JOb/ܔS��G�}8���*���h�kiq������j��g��g X��4��.��Ϣ�{16�@�X������|���ZR�zHS�� DS�|R�������;�\�yh{�c�8'�P��j�2w��B!�`��p�i�fK��� ��l5�/��ά���X����؛����HL��[���5I|��v(�e��J��V8�Y�ʩ���gw2�S�,9�E	<��=qp��wԚ�)w4�X[V8���Ze���&�s�	H�M�ꩩ�>=v��o1Wa�g�/����|����<����{�+�2l���}�l5Z��:�C��kd������0%��Z��7�"_�N�4z�
}����X�"&W�!ӧ%���==��
�}lg�J�`.~��iCf�v�}Zzu���8��8�/�)��D���զQ��|���PcVGdƎoYp�M�x@B�c؍��d�����z�{����N�Q��K��T@�Jvv徹�P��軑Z�N5��j$�5���o4��KFX��'�8���W��\H ��T��vK�f#y�.ʎv��M�����?�a�d��݈�N����~TJvS���u#,l"w���M52WM����
��1�-�*�i"��:�qC��Ƨ�~Az��l�\}jR �~�3*Tn���>��/M�Nˎ�y���s.��*x�9򄢗IB���&BRiL���E�՗^��3�P���.�|O9/���������;ρ(�z�j�n4��#Q;�_'3���P	��F}��3�YEm�ť��Z*�e�݋����]�z�͵H���0(��4ñ�,֞Hzn`�O��`��l�F���Ac��h���L�\}��sӨ�Φ��Pm�b���-a�Mg��H��U��,��s0�>'��T�T
Iݓ}m��ּ�*P����v����\��'	�d8��m��
��m�R��ܳD��v�g>��_��?��@ʡ�8�9��[�}��9
4k*)�v|��0��&���1�yi�
2�������܄<8�	ď%�z{��W�e����[�.������T�O���t��!Y֑Tw��
p���v{~��i+���A9��lCv��cW�:�@�	��m�hi.��w�~
(C��<h�pp��M6�+�m�=5{L�EU5ϋ�
�MZ������c� u/\?��pc�$7��'Cw8�ƪ�C�:U�=]�u~�1~�X㣃j;�n�Ic��q�,ϑ��ى(H��)�/���с�`\�p��v�s**[�V�%RKR��8��n�3\%�:��O���)q��'(OۤF��e�6�]gj��FF��5L�P7%�Pd�\/�]+�&�nwB9��jj`�
�o�6x؋��k�k�mP/H�z�`��̞8�i�2�iJ7^m9\�	�g#ԅ�}�N��=N�y�٭p˫�р�R��)�E]�$i���?���O�,���<x���B�؋���˨!$�e+ȟ��0�s����.צ���AX��D���8r������o�E�f�69�B�5��~s�ne6L�j�d�C4���n �,������T�C�ɯH��-��C5�6�\|�v�0c���ל�²W���Һ+�Ѵb���͏�2oqik���Q=��ol1�G,��p����k�J�/����go��ٵ3����1�>I�Ed&yW5o����LV�6�Ͻؿ��)~�\$dANae��jں��z�z�]�x�#-�x�tiF�ͭ5.)��p/���*�q�.סk�~�ĶGd¼V!p-������+(�BW�>�?��jP�����zAH��v�	h�.�_s{p-u}���=�k��9��ݰ:��W�>��x�!]���p�P�x&�~�B�-x�&�r/�����v��A���k���F�Q����`��]7�:aQu��b�G�f���H櫷+���� �7k�|�uҞ{7���;��	E����R�k�.�^<�]C��S�?�bǫ�����~A�k�n�S�c�L��$�.�*P�)�s��a�̀1�;.���O���5G��po��n��y�W�������R�/�h6;k�]�]X,�l�Q��?r����e9?h\¶��J��q+�DCǈCD��	��nϧU��F��ʰ����3S�~���=�VʎT��(F�@ȫ�p��A�Tl��0$ �0�9��yѯ�D��^?�E�(!�ܷ���zņn�>��'fS�a7!����qi�x��l��u�93}���or
^�:�/��z�Ô��œ�r�<�H�Q/./GN�lv�J��w����zb}��
��0[���g}�q���<�[����}�s��]�����4�v�n�v�w�a|��@�u���I���  �uX�EH��x�JU�G�z�H���=����1�W�:�c�F��n��[$��\o�kf��P�o��k���y� %�8�
�{�w&��Z�oj��+4�>=?�Ǉ�d��Kݼ���
X���E-Ɖ���Q�pHrﯺ.[�����C�ޗ'X,!9�����
�d%�,qeK.{���hN,"^rRrA�q�8A�|A�hj��F�>kZ\��'t��4�X�̵Ӽ�lĬ��:<����Q���:#�7/!�����˳���΃�[�>î��2\=2��?&'Ǹ�i�>?�љ��Q\�읡�a�R�I�sN��(֎(��vT/���.�)�:�x\PWzJ�Q������PDIPI��ڑ׽�G�)R��2HN�UqoL��]��`N�Z����X��d�"W�(���h�`��臾��U��ow��������PŤۻ�F`�������d�QBн��y��/#�)�l�cR^=uaW�Su�ͩ�;�S����{i�h0�%�4��B���A�\��ײn�̬\#��:���,����b�#A�A����"����}Sа@x�Zx�{nl�D��.^���g�ۣ	z?[c��^ ��®0�@���?�D��Y�$�p�:_6Y�݆0��$��~6�[6Q���������^�w �e�|G 0�Ι���E�J$@U��9��Ń��PH)b��5��[��!��D��(�w�ȇ���	I��<����'f�Fvo�h�N����o�;�TsL��i��$�k~��[ )���}���V5�$[D�e��T�v�O{��}��"�;�wC�d��Û��٥F��Սc,�go.(�K���9�u��XkAU&(F��1K��	�q;o䃋F��恆o�rN̝��Lk<�za�����6�Dޣ��UF��ӱ^�_�l����
����$џX�к�ŻM�>u��O~���n����ό3��M�5�"�z���iX�bZ�d���8|B�gtb3�	X�hE���~���)����~�ᮢ����Me�������	v�9�A)�%�b��ώ��y\��/��l���*~��8���'�v�m�ߙi���������\�}�(�+ry	٤5j)����B�ua
�*vY()K���a�P=_ٹ��!��~��ۯ�0����;#ص����r��r?���WĒ���:��Nz]����D��g6s������I�a��CK�;`9�ǪڰΏ|G���8,�� -!�R��e-3�uD#�����H+^��ղi՛3E�:1X�$�|�*?$�:aG�s��զ��~ʶ�D�z���76��?�RX��RY��S�
���B�LY�&̐�Bʏ�������Vo�7Ju9�yuH ������A::(`������Z�
�A<����ضV8l~��k�����u��R��6��ʧ��WЏ�²A@|ӝ�<䖴�
)gQCH(U�^v����
�#K����kKc�q��S�7p��-�B�hF�+��dFG�"/����"�~�ݰ��彣}��z��Գ�e�<��g�}���)�K�E �K������m�7�4|V9�$�^Z���������í�����Ty�
�兿�G@\	�e�?�ejs������+i^���()F���7$o��zҫHq��6_�F<}������?KͦTR;%U�筬��`�Gg'�̥拯����[7A���;d�6R�I�=���a��:o�����˷���I�r�����܄�ԥ��/)�� ���/�N4��R?�g���-N��<���=`���n`fN���Q��(����	��Q���su2c!�Ƨ�lu��!��Κt�.P#��|��R���j@z������{#̑�L%�t6��"������[*�\�F}_㋄�C
����g��I�*���Y9g�=]�c�JK5
j��˦��PQ��I�w���~	���|W��Π۞��=��s��5�0�͓�C�+M/A>����+�h����۽��9���Mo6�Z���=�Q��vKO�{�(��dd߇�����Qe�i�����Iy�D���y���d���_R���I�n�L63B�����0�0�iB�[��<�����͓��bn���ɟ���CKlș��>6�
��Ѧ{���]���֛
4���-է{��Y�ۛ�*�f�O�H�g;H�����p��GgT ���
7E��Y��C��M��b�A4=�yk��˂�ǉ9����>Y���p�B̓r<��tY�<�h��΍�fk�n�\��L�\������˶�\��׵G��R���4P�L�����l�Vl1��[T��/�_��ʪ�Q�j�������坱�� ���*�kQ.�r�Kf�� �Uh�-Uj��v�D	�tC#M���9R���=�d~+�S�0	O��Y�m=�<S|cL60��vt(�Hs��ցty�r�Uϵ�����ĩ�'��?�|��}��	�<C���@ +�0�o+�f��: �o[✬� �4d��1_lTPԥQ�H��:X�AQ��;��vAK)�X���I`o��ȏh<�N�:a�p ���t9O�6}�}I��Ɯ�>�zvw������pN���\O��}�ɟCb0���ٱ��ߞM�{��Ir6���=�����|%"a	�+b��������(ׁ�S}G�eu���[ʹ��6�f~�=�]->Dlㆩ@��9/ְeBr8>�Az�Tmr��c�N���>&�V=	3-�*��Ӹz��q�ݬ>'���h�@��U$O|�Xyf>�ܹ�����~Eh�����|�K����<��ܫz��T�3�
h�=q�d����w��k��&��b����⚺Y�V�� �,���"��`�ðE���(�	�9eX���i}�g�c��q��0@�霢��Tsk�*	�D/Kt1�H��ܨ/�V��t=�cc���m�m9%](^��_�t ���A�J;�=(����6J�6�{ͳ��S*��IJt��^�Y��E{I�?e�\���f����s�L��{K���g`uؚ�3�{���0
`,���6��X��Z| ��/])���m�7u��߱��`�:ś*�������8<IE�>ߌ�������p Y����Qz#�� ��z��Uv���_���;���me��[��r�����!ڂn}6�H��PH.rý�T�Z��@���	%�s�Y�c!\�� ��r�Q���G4-�OIjdl�%�t�3�7���]=�mɗq�B��!���_l��i�Y����f�� �CV�"��B|ޖ '��d�[-�_����p�I=���ުCr��w,eҘ�#o�Sp�`\Z�����-�<�,�����^�k��yl�,�I&*hi��!�p�s�ayŋm�߼̔�Jx�q�sA�US������ӠS�������>���v_4�wSk��lfK�v��V��&��B�A"
?�.ߟ6���T�>����Y~�"�/͚@csN��t�UQ�|CHJ9;4bI֜L`(�D����s� �wEs���x��5(9�1� ����
�T�;�߆�U3� J{����P�6�;��(n錳�[a�}�w�ͩ � �v�ҋ���iY]�t &b����2��'�7=m\a4��dW���b�&z���$��=r���Wz�R�X��x5XKG[��g�L\�������G�ߤ��������d���7��!6<�'�|�zc��p��p���U|�Д߬E�)��^x���!�5�VR+=��O�`�%��G��4����y2��O?�n�zH�h)�X�����S��{lٳŚy��@�K\�dȒ�g��B�	�jǿ�鳻!���c��]N�M�T��Լ����G��$�N�:I�:X��&.i<�M`0���O�
���A�'�lӫf����

�~.�!Q޵��K�4�����O8�i���΅('�B�y�4EM5��Y���y�J�(����@L����\�VCv�tQ�2+�}S�ѐN��w�&
�Ɂ�y��
��A����.��A�_! �,���w���`xu�w}�4i������,���S����ɗ�����u�*��y�f���r���f�RT�";������RxZ�;� �P�jr���ܬ���/��h'H��I.�G��º�{ܜ��@5"��(���E$����Oj�Mu�s����gt����I�_�:mp��#���"���x_ ��r�]���ϗ��w�now�N�RuC�'4�,����\��7����ҿ]�%ڿ(� ׿�����t�����<�R�K�8������˭�H�
ɳ&�Q�aNFC��:�H7$�ky�]S~I�4nm�1�4o��	���a��S=BO5�|��x�t�P�`�H�k��~8��P���!��!�l!s��*' �<U$�$~�H� ���)��sm(�y*c>!�(xg0�0���ٺ�1���j�`z\�9�Z^ѻ��Bq�e5����'C������6v����<E���Q�z��v���t��J���h	|ǲ��0'����I�C/�����z��m{��i����qX�A6��q95D�p1�w��]M�TS�����e6 �Q���)�NhU���6a~��e2�
�Z�Qr6OH�����{C����ޱC�<L7_,�T��t,>�#~K�o�����������B���c����x��ZdB-��л�w�pP�3���1�18�{�s��qa|�Gr�N��N�B��	<��=��)���"������;:w
M���DeT��θ�O���,u,EbK����t~֩�i�K���n��?�¯	�{�������H

c�����JIIL���0]�D���1�a6z����y>���8���:�}&�����Q��_�h�R�� �r ����c/xk��,�~­0�r$A��=�tk+5{)r;~F����)�������[h�B<H�B-�xC���/#]-��0�5�~U�yX��w����t�i����N���gt֙F��M�p�*���B�)�n��=I������S u�~^��*�?I��]Z��5:'L�7����E<Ǝ��pF��m[w��Ml���S|��V���`��ě��_�O��l����T���gT�)�Ĭ̂��ˁ��^�H&�ã~�V8�*x�s�b��îlnO�.�=�1��q}��{���W�P�T+�5�_��U֙�D?3�]�r��T"�)&�P���q�t��6��f��uu���5�ia������%(�C��j�,�pm���贼R'��?�Mm�[�	�h�i��2]�	GU�����8�7mD�g`���L�x��q�d�~}I\E�<�S�H<�_7OE�4�9���s_�7��E���-�
�6YT���k�#:�Z�~j6�K���}� ��oof"��}Vʺ�;�mI܎�KF�ŭ���B�֊���Z��T����S#N���!+E���F�	��Ŗ��c�Հ��cQ< PQ�f
��d���e�����Sv������|hQ{R� ���qg?�)F,%��־;�FfLӱ�r*�5q�L����a���!xP��\���uy�Y��Yb���n�P��{�²�����
�f�/� o0g}#�W���\ᴥ�>k1g�#���X_
���@��7N-zk׫���[�[���^I@�q��,U�3�w���#�2��(��,��FBy���OA���*��]�Q����f-��>�������2_Χ,�螻����1Pp;m�v��l����(ϐ�Ih]�'��R_t?���0�(�HN>�֛{q^s��g��1��2?��d�k��wO%�2g����~�	�ԺjӺ���к��ɹ��tcC�)�s:��:ѧ��~�.2Mǃ�g(y���x4�q-����v];-�W��Jl�[q���Ty�NIA��S7��G�U�G���!.[�Ry��0.��,7��6���t@��a%�R,̗H�s��ٕdH�l��a�Ą��͇bN�H�Y�ֲUz������̀�\�[���ڄ	7(<���������m�*aU�0S:�AF&���n:w���~F]<\Z�<�2^�u,�ڿ6�i/�l����I�;�OD�-=�Ľ�i�T��=o�-KLb���`����K�Ř>K�T��B߀��ܖ�w�� �
�M-�xڔ���w�p�LH�d랂�`�e�3OK�}{ny����Gy�L����EL��F�f�ȠHu%X
�pч����-b�f��!e�7�U�
R�8�tx''7��s��>޷��ݛZq��'�{�(ʸt���C�:��Y���}��Z�������6�eg����-p�7}tf����To�z��b�Cg��!�����{+X�:����V��{3V��o�g�J/�fj	F�e&*D�;cZ#;�C��b��	���w��]��1�u�+A��8�7亷�Rf|�r�K����J�j�홐���χ�1g�ȯ��>Yg~J\�]^�&�	��,>�=�z� J<w3������Qۄ���T���i6����6����j�V�������5��a�	6c�mzB8��MrT4�4H�7��i1�֬�卣�_�F�/ο���k�����rIj��0��f��9��h)���zv.w}��'���YA�̞�R{�}]$E�F5�fN���ڍ���#B�Ͳ�������LB>N3 �����kZ����d�����o�7���U7��y��S���Ʊ=�ނݬ��_%
�)�:����nsE�O>��[��f�O¼6ܑNi�s֞�U_��g�-iV̨1.,��A-b���fq]�9���#����^�#�őZ���&'�W��ʜ1=+�d5��K��C����W�]	������ַZ��.����W��Vdb-8�Q�����%&�l �+�l��c�v�*}p��M�oyf-�8�������s ���1��rF[�����O��گE��7�=$T ������vPdIٹ�ƈ�!�|l�}��c��E��!f¿c.ɞ� X�����
6�3�[�t'�}��Mn�ҙ�@��<��T��[�P"5��.B�OZ�e%�ET@/�?]�3݆�FYv�w�o��V��s��G�,�!f��s����Z�� <�x�8�����w�r~� _Y#�.S�q?��'X�4硰dJ���%o�A��줟Zf���4N{��\?:V*�4@͢0����5Z^��Rj)�ˢU�x�'�Ɇ^���:�ϔ����|�R���B#L��?�<\��x���;f�"HS�=f��6��Zw��Iv�����F���{�ǆEa8���շ�R����OK6iٰn�u���&Ѫ�ɛ���l��`@�:FZp�	�UcDO��Ϭ��Q<��m�����h�S)ߵ�gʮ�ro���~]�OP~Ex�ް��*�3�r��;�
X�jMV/�[}���}3�b���(}�c���Bѡ=��q�}�{�J��D��K�PTy_�@�/o�9��v��11�	a&�>��ƥ(0�����*����j''�H�P��>�:�>Av	��LUD�^��7n������8���=x�̲�h��Y��TKr6���Q,�$�'���U������x�ĒT�2��+=a+7@5����EV�+?}��WSʹ�L������?��zƧy~���p` �xv*&�4�'��7��2�����֔���UZ��C�|����;-� mmYm��0{��6z�e��F�mm����k305	����>��W��4H�^��* ��7O�=�����$��͊��C����N��
��hۣʊ̷�����LR����M�ۄ�Ҝ��Wj������'�pN3 ��Cuk���ּ^Y��_�j�OǱ�gI�tx2�8#�e�����d!�{`��u�Celc�x�l�Y���	ǁĹ�K`�s��堘�?]�_��aԉ�,�|�̪l�e{�29Ƥ����@�t5$L������ý�	d�t?��pl�9�D+/ �£߫38�)S�,c?�����n`2KW�e}2�F�<o�x���a��e����4�]�/�S�Ai����_�q��nh���$V�h9Ha�1]>e�C��՚a(����s_��\�b)w*�M��m�������m�κǙa����X��@�iV�)�j�*����h������=����wH������I$Q��h;��n�il̶Y�dR��Gϑ4�q����m���:��kǑ�@5}��� Tm	Y�|&��o1���������N��1SC�ͯ��^B׭�*M���m>����s�F�zW��r����|����؃<)�W[=e"�]��%k9�k��,Ju�I}�?�W3�'v��7'g��,&�jL(�m��Xr��A�42\+w�h��7�H�����O𹀒���=$�7�I���o2MbB𫕢N�E�=dE\���)��9d0�OH@�i��tfBL��c�e@�}i�_,��4��n�c-�36o�F6�4A������Ǜ*L`�^�6���Z��g5�r����r�]n��5��f�O�E4ݰc��3�wi��:0̉�������/�x>�U�:49�?�@�rה�cNՓ~�����|���V�\[�H;��w#�ɕ�ivi��Eu�ަy�%@F35�1��ǭ
/��O��<����j��m�i7q�v�E�[;�QP� ��x�ƌ�#'�F�B�XJ>�>���-xB���@�<Y_��SX*m8Xnß_�� !#��<��T}/�LV?�b��1��2i3��*��^N�z���3��6{��J�U`�b�{U�&`��TE"�Z���q�,g;�fS�Dz���e�H7'n��^��#D\�J�o\���Ĕ2�K�6tn�����^�P�Q�p���FD����xHm�&�����_@�h{�3�{�º�I4��������i�5E��r���\����DƋ!����k�GV�(�9��V���NZ��[����^i��_�����nI��m������nT��*8���Z�\���IWՕh�'�ϨD��G���Ii l��}8��M�ُ\ �"Tqͻ>��;!�+<��iآ�֔eU�l�T;���jY+r,�yc�}��?���ܾ>��8AƓ�:�d#��N���C��t>"��=]"�4�q�X-��q�Dk7�va� �� ,�)��i���v,���Ч��w�z��s�[R#��"\�e^�x5��g���/�t�kٹ��mx��_�f�e���$���ɢ�; e��H��ep2�nd��4��#��7�(��{^0������M�`�f��A6��y� A=�Q+(5���N�ܨ�V�=��'��dr��p:6��&�Q����o�+����Z9e+���en������M�����$��$��\yԏ��O��$g+��ߏ*��9I/#=�H%���c%2N�2��p����s�Me�"|��ON��N��)�0I/�l�!$1�:��;�6a��-V�Ks�4#��M��7��	��O�TE�us���f֒G&b�)
�?�փ��O"*��ϸv��7]�JQl����8G����{�湘
�z�i��b��*/B�G�L��x�7�WdVFCxg>�̐�6��v����lu�-� ޥ�',�K��]/@�����]Ē��H��u~V��ʇ�2�!{�6�;{s�m�bM��#Q��:�������w�YD��.5a!�v��������aЉF'ހWnyP��h@_��0���4b]��_Km�F�԰2�^K`fI����OVH҅��˃\{��4�[��{��>�%l��;뇿i�G,H��m!? c���tU��$2�NcK|	�O\뵦DUyu~��8�ag�;�"�O�y3�ld��ޑ,  ~"� ����Uy�5�D����G�Zyߝ(�\Ѫ�1�MAu�GG�%���
,8Z�����W
,k��ԅ@���R�i�(�c����菘κpAmrJU��{��4Ҥ�1&�^+9����HtV�,oZ��"
~�_i�Ų�h��u{]�rE��yTu\���$�1�O�����n��/W�G(�o�B�/0��鎡���=�&��-����ש= ���ONy��o��۫\�jq�3�_��D�]�=�,~��G$���QBā��|2����s�6Lxf���|�J�R��Y;忥8���VE��hWǚ���z:NLx��9f��w�8�	f�Ǐ�y[�JݧF:]���%NU����ҰZ�I�l�`w'��Z�����2�;���EKrW��1z��/��|�VM�)�ߗ��')�o�V�gr���c09	��JX����>.K�?��V�TM��:���ϳ��`Ҟ%����cĪ��$(�//Oʕ��ݸ7>�������ث��oL�<������K���d;Dd0�ZĩG$����Ĩ<�D�*w_ec�N��e�E�����v�-Ը�8#�6t����P��<҃�������H"y��&��Ӂ��i�Ql�:7N�m��Uɝ�?^W!#�A{�U"��[������'�V)]o��O�O�{�0_�-]X����7"��C�B�����"�R��S�q�3���%��\����^#ұԫ��D���Ez5���#��Md��C],��f2^����)��<�fm��[�D)Z2P��`�����������g��"�K!xL��D�.�w-Ŝo#���=���.5��b��&�Q�(�x���8_�a�j6��Ǻ��}S��T�IMT�Zp�5i�#q�^L�]t SF50�L�w��%���{���d!�X%�r�躺Ԥ4>��e�z\Z+cQ=�+9���5Seh|a'�a�L5�k�Yaֲ�-4�~���c���k����kA���0By�y��^��W��<]Af�D͠�¹�w�2��ȑ�6�]t��5_l	>Ku@/��� �����D���%!�O&��]m�-�MЍ~�ʭxi�eu>�uE�Q�q�I��X�Pޓ�����d�������6�FS=��*�ݻ%]%�L��Y�d�cy�v���?�'��`�t�K/����Y���+"��f�EW!��?��n1�Uv_�iM�a�C".��Y��nzSH*eo'i�� �@��z" �X�zX2򦔊qW�giVsUq��mbM�$�N/87^�of�2(�Wiy�}��yj��%9��\ƺJ���k[�RV�����nc�o喵���1mr�ج{9���=D3|`kwt����	Sh�e-�5\M�{W��%�Y���������Rt�%wA�8��T)'��� �OX�O�h|�!��[6k�w�[H5E��o�7pB'-(d��E��^���)=��fmI%,ʄ��@"A?�䅾��ʴ�q�MK<.�	��X���R�+��=���7.��˴�K�|�s�����ݪ6)��-W\+4}[�w�s��ߝN��CG�/c�l�����t��S�~z]�	�\���~���p�^���Jʥc�"�"��:UD�;��!�����z��9]1�qz��E�}��4U�|Dq�6�ٳ�l�W��5l��*�����?�b��$*��n�z=�:��J�2N �P��������*(��A��Qj�5����m���}�M��i⸘g>�K�t��긏�t�c����0`4�b�>?XM�w�5|.�5|��^��Y���,]:�C�3�\豮24��T#���0g8���7��sQ-,}A+�)��m��Pq��#�}���-�a��t�HZ��(9�PI�z����%j)f�5����q5�Cj\�0Bxh������9K�aaMT����v"h�6w~ӻItcW�P!�Ȃ]x��nY�F9�~�1�����̐���a�2[�g������f�J_��f��+���b���ھ��܁q����0~�g����
Us�M���w��x�o������E������j!�T����Ώ�s�/"�w��ځ�+M�
<�^bq_cі;LR�A�	�l�=�hՍ,n&rDc�]9.�8p�M��0��]38mc>�h�ͮ>U?aP/����cC�3�"�5�c~K*�c�+��Z#�Py���R�`�v�])�g�����i�?O���i�6U�ᙬ歇���ǳ�X��.�=����1���.�9��pYZ�$����Y_�[bA[x��1��A�E��r��c�T�b��ư����Y�?���<�*�w��8Iw�V1��F۹��l{��"�L�SXy�K�	�E3�情��J����J��1�y��V;�U��!����s\���x� tF�
u#�@���,����V��B��gCx/�V��-��8��&�!�����:{��ZjʎD��U�z'����8�Mh�2���VO�9�EŬ�U<^�N7
W(��$1W=)qz�;��0W���Y�ȗ@<)�M���U�g�R�-�f P����;^��̫:��� ���~�G�����x}�0 �hY�D�`X4q��%cǐx��)PA��򑖿�6�E�����X=��:Ǫ��
���>����NẂ�f���S�Y��������կ,�.4���{�~� ��E�пx����PB��J���CzDP����s�uЇ��{�[�x�v�!hd�������<�o�����҇oeNgi���z;1E�NwD��t��˿��̌���|J��YP���x��i�B�m4n,40���4d���"�L-㬈�xB/�s�}���l*R�d�ŝ)@8�U��$��=��ho-�Ey��[���-�����Q������З�ι�[B�*Y��	�ӊS�N&U4���O0�;�<D��F�2P<� XM����1��4�WpŠ��'����bz�K=��_�P���{w��x�߹���<C.����#2bOT�藦W&��S�'�v$Z�i�,��C�X�K1��y�tQ���pq���u˲����1��ţmbY
��ptL'sf��_�b�����ݩk��5}}#�ֹ;%ə0�����������}N><�ܝ?���OQT&����Vyf�ͻ%ר<}&_я?hj�ŏݿ��fz��Ĥ�sL�G��^�r�Op�D�6?PU^-���d~}�����e�,;)D�_�xo>0�����V�֔��,����ݽ�K���2���iJi>�~+��KH��1��%X
)���m)Ƒ��� �!Y��Ó�nOR�b���r�i���/�u%#��NnNI��BC�]��9�k�]�M|�Rn�7�\?�X�;�?WQ�6����׶��8�6P�v��T�%�0�
*a�y��C]t��v䧿��j��x:��R�m�}�hY O]��:���(�R�_Sn�p���N�d,��d�zt5��x#v��ȓ�C�1��kf�[����kEύ��*Ƭ�2�<F�΅MJ���n^3��w�)������Uq:~UfR"�:l���$��}��C��s�����F�������"��kۃ�l���݀gz��pB�V8�Yp�^�H��<� ��֬�q+����I���z��u�R�s�R�G�5zY��}"�m���TF��E>�2�	q6@E����v]H$�vm��Y܇����CG�<��I��,x��'Oɧ�_���9�$d��2f��N`��,/�U^O�rAR��6X���ѹ}U�[���M��OQ{��8F�cH��)�,���:���çi�&Ý�2�|D0�����*�:������WA�"��l�M�&�X���c����(l>���fk�_�����E�������}�A󐾸Ǒ�5������9��5��4!��C�eW���(��^��(�>�_��֣G&Dy\����y����{��/l1�|�/�Ӏ�Ќ���	���3��\*����o%���4��_M�,���N���Ok����X�K��b����Us���+ є��f�ufv��)�#f7�ٮ����4�@chⲝ�T�Gw�K�~���Ew�Tt�������@"s��#gJ/{d[���N�+�+Q[7W�lݮ���}-h�!�')�ǒ�߸^���k��8u	��?�'�Hme�"g�ͶQ�<�nuG+=�O��ΰM���/�R*Ř���O~��4_�~�)�~�l"=W@�w�T�M����g��v�k�u�>W���r}�bљtי&���3�sw��y��m�&N��]w��^!�Y�x���`��o8��E�a��XJ�0?�Q�^���%'G�bz��-c ��s�>f�6Z$�]7���+����˔Kf*�~3�������d�&Lu�V���|���e=w_�a|�����}���n#��vE�U���O%o�$? �kW����Y� ,oݓJ�UX=#�{Q���꬈J��h�����A�'�c(���K��Zd!՘�.�~PF�
��F�sUF�uB���!C��iu#ڞeuf���51'��R�iDB��;�����fOZ�l�11�xài���m뻙K|u�#��:| :IҋK̔|DH�cR�c��ۂZs�~
�4��Ǳ�u�:��V�A}u���&w���>�����*�_���SS"�F{K��Ih��/?Rǃ\�_���rh <�&��z���ٚ�Ҙ�K(��\��N�eR�1ޏ�еʦ�M5C�	��2W���:	�xx�#��I�l9�BQ��zΩ�y�ك>2O��&4Y	S~�GB�Q֣I�(?M�ۯS�踁$� ��j�"����տ&e��������ݘP#��������
��*Ȫ�C[�~�Y�R.
�g����w'�ǬA­����0����y:���w����؏��v*j3?<$m�ە�f��vQu�s2"ŉ4]o��/�]$������Yk~r�^��f��:ö�o�u�4�6�����+:S�]6I���<�\� ���y�Pz޻^��E���U:�G�����^�0�?U����K��43OW�{�
�� Θ��nu���}/�����yv~D�Y�2N5��ij98V��rH˳@�I�{l'�GMs�Սˠc���77�TlAWݯ8#�3�C���)F�j�P��ۣ�$��2�6����/��9�N��|�c�����2�:4�@��%��f�|�V�,6�3g2��Z����_L5b�]��
��Lj&�Wi�='P˫��?V��W��s��B".BJXE<��kT.�L�z_j�=��K�)%��4j����5�7�������/yR�H�d�w$'WW�)`a�Gk�7_g�f*��J���6�Y͠�<�!,��y�N6��\�;q���K��x�\��5�c��R��}1�3���ʺ�zG'�����Ňi(����Y"섓��Io����d>�AP-pKa9���������m|�v}Gn�u� ��]�&wWuҁ�%�=7*��GZ�b�̝�|�� w�9��( p�Ic��n���Q9z)��S�kA�WZ��6��:��)Lm���:<x{�����Q�7�>GΎ)ս�+�����M�׸xɷx�Sj7�q�uO������̝TjۤP\��k�<�g�sm������6����c�/�[�p�U,����~���������ʴ����s��{;w�7������iO/�I� z[��G���v��d���,��t�sVxX���ge>wBN�N;Ur�j�P-Nxr�����|�
}:|���G�t�\�7+	�mU���?E,NG��P��>�1��+��,e�d�N�q�i��i��S��A2��P��O�1�������.W�hR*͐Kb�5.uj�We_֒ܨ��V��7���4�]R��$(Ŭ��?bn�+�&P:O��a����`Q��qH�DsHCc!�lg?�%0&�0�k:���Y>/ޑ���d���w�9���(!S9�����tMW�N���Ì}
Su��ٍ���J�����9��u��@�WdgW�?��V[*�9dܦ��`�P��#���&�:�	^���͆coJj�1���M��i:�6���c��W�c�� ��큩lih"AU�v��I��kb�Ή8���1�nt�\�q�!��?b������y�x����kӠ����B�>��;]�!y\��v�C�Wx����1���yxU?�k�gQ"�h�1u�!�ـ�zoPQ��W�5�-���(^[��f(��!�-"����\�/�F�;��a��|�<�J��W�`�G����B7/�
��>�����o<+����k���%�x�x&��%xѮ#�e��Մ��-�Օ7�?��?>�0��R�����,�>P�8�_0ܑ�C��Nv����m�L����N�M䬹���9�ng�T߇�m��z�He�	��,p_��mNr.�=h@!�[����h�ӹ2h��
N� \��O���8�?���ʓ���?���D1'���-�&W�M���+ڵ/�xaz9HG���)|�v��hC�|I�p���7��*o.�Ē1�V@��1���}�]�,�g]�lflWM� ��ݽ�[���5)�ȔZSGrq_�F�ˮ�p��y�5�b��j��.dO�O�۶�<�����xm���uO�S�2�jn�n�+H���]f��&�) \n�z�Q�#�J����z���<���&���ߎ�S��B��/���Z�a�WrmnN4�2[��_u:X���K�O�|�L����̒	��{��5������g��2�@�'��
UX��0G�Ve�=��/�ߐr��i*\ݔ�N'E��j7O��M=c��8,5C1��6v��������5LR<ks�,1VM�Z��?Պ'�I�
����(q��q����ës��t[A�%�k��c�+�|&�]��u��X1��_��EQ!z#���`+��_9+�����o�V)t$���Se�`0l�VN�W^�Bq�|��,0�8z�rD����-
�3-���a}��}�wc��7�]���Pq��W��L����4�#7r;��yR�bb7��{���b���VG�\�S����f�S��L͟��TP5������؉��=�W��'5�U6�UeH5�4�yMI�P��G�l��?�w�{x��l�ZXq��k�lpP��Ӏx�v&��4b�$|vfbl&h���a�������},�ś���k�&���.��j|��\���[Z	L�%�5Bu�]��M?���1�!<	9��y-b����g��VG~��L�H���o���s[bQ$X�
��C��A���$�)�m+�:�����GSk���Ld�չ����G��*o���R��9�FxH�!1g�T�aוe�fC�(O1+����,z�Ҭ��ۉ� ��n�l�ohK��=��X`�Fu��hn���W�1 $m��۲�-���1mu�hw,a�p�kt���+5ċa��+�4����ՖS��փ�Qe��\���
gO�Namsb�����;�Mg[��H��^;a#�u��ᛴ?��U�i�$�"���Ƥg�r��]��%���kKR��
^O�'%�D�KyϏRs�x����`%�|,(a�C�r�3E!j%ƨo��$��}����;,G����T)To�~ �V18bۢ�<��V[z?�C���e�R�EBe���a'�?���k��e$������� �֬{��u�{)�c�d�sP��a�i�us26�M%��Cs�O���t�>ߋ14/a4��ʤg�Y�!���J�'�!�U"q�2	�R��w~S�)����~])��z��*9/�=2	�����ny�;�#V �y��P�W�LD��d�le��X'��7p�������^�>�X��;�z��W$t3��W��G��o�b�W�7����Ӛ{���'h}�b�8�߈&kz&��E�R��P�O��{�&���gB��4s������]�	�!��,�r���i���SIP���i�q�M�ž�s�b�=9��n�:�яyN�\W �����:�ǒ߭��|�w%f�!��",�h�w|�o��p�u�ZE?@�JT3����<!)Y��3������.A�yE�㯓���t!E���o��l�)O;�j�i~�j���q�\�6�q�����e�9ox���Զ]5�ɳ���8�R�*Q���-�D� (��1�M�����;f_���/�e�N`Sf��$�J��;���
C������@!����Sc&�׀�"YG�ZHC����Ι�{%�D����\g��.���3�pPC��W�3PZ)�s�3��`��s)Z�怑1x�V���w�aJ�ڻ��g�un�!��h���h��g�ѯ:5��*�#P[�!��� �syC�C��5 B�L�i.�R�I׭���>������}��v^������E�c�������F��Ҋ�mK�^:�@��۲3�rE@�=݆��iH)����[��Rwj��q@,aJx�����/Ο�Ȉ�m����{ضVG�U��?o]��Q�b6gp��p�ω\=ظ5��g���ɞ"����'BK�ŬY�O�D��U琸2gd�T���֍���4��ի�մ �ni��������b�x������b�$]��;MsΔk�6�Of�L9�&�W�hӥ���J��{�̙��b1�3@��?dTT�x�Q����UeV,��_[�/�s��(�c~�\�W�:V ?p��˔���t�C��'�����$Z�W�Wi�J��^�����d��Eo���Kb�A?�wV�t������e[�Mj�[�8BfC���2ĈC��0����%t�f|��Q�+����s*]�#UϨ�v��=����j߿љJ����
%����Ժ��z�R�(�X�C��D�9Z�gLT��X�E�(�#�m�#���Q���gw�2t�D��~R�ݴ���FF
9���
K�q7��v�q*JKwy�����wk�<1���qh95��|�0�v���μ_�[1o���8^#�\���x�O%scd����w�lnͬ��K�UE��6+��^�Ҷ8�h5���2T�R�?�t�8�����^�Y���`�C�O̗���F:��X���ߗ�
���9n��#��Gu�vcLh۳z=��IO�[����0�5�
�ю3�!t/L�d�Z��X��b3P;2�|X4^�;��(�\�m���[�*mP�be~���l�`W�>�7��^ȁ�nÏe���M
ImR���+����.�A`z�~sNN�QT���;����*���|�m`�+٦��Ih��Kqzk����BPA��z(��T������t�D�B�n�d?,�i��m>���2�|�ʳ��h�C�����~�t��b��*�Q���=�vr���9���o����5	3|9O 9�K�~߬��y��I��n ��`�Ϛb�3Oy#��m&{�S� �y��7�1f�*�tHH2���8)�]��G���H5���	�N62	�!ɵ��/y�k֚,F�/
*�i�ټO�҃�i>f��\C�����wϜ�����h���g^ֲ(]�p��SM�l�#��j�欸�Y�G�;�����F!?�=���`i�.뷿�'��I�B�F�����*�.�L��p�؜R���@ũ �D�Ǩ���m:�	/�
�	E�,�����=�ۥ)�k\�5jd@�\�2y�n��-��
��)�# ��WjCc��K��R�p�?��t�_-,@�	l{�{Q_��U�w'(�~Ԝ+�{���nj�-��)u�!��86�x �ځ��CtX��rJ��h'v�[����'�J-�l2_��
�?jU�L�U�j�0�"'�J�T[����x��޶�Y���x����s͂ҮxKTb?O����i��K�_�n�v�L���O����D��?�qeş�y)|��$�)`0s��7�>Y��ȒO�����z�N�V3�����}�t��3�Q��h��Gl�Jwܠ��pַ����l�!�b�o��Y�q��p��<G﹁�˯�ڢ�7g�����K���d��eP��p�eY��O�ky:��O}��p���Z����It�����]�K�b��܏.��jHf=tGH6��� .X�r���X�/��_(���Q��Ƞ�l�庂�i0�g>g�>a��H5�'l�Pٔ?��X�np�8����5�Uf��@[����rUS��$�|y��P�c}|~�����U�8X�|�Y�|<=�����8�}fЄ��~L��P����n�3��Yy�9Hd$�t�k1N���j 3�t���N)<X��fz�&�ش'] �˺�ʊFD��ۡf�}�I%�H��z]��"}����3�d�û����F�>�շ<��0Q�b�Q��KQ�$�	3�F����1�VA=��|(A��"�.s~ތ��}��]�}��L���*��>Y�wK�Z�����+VIoE�7��㿬N�7�������fԕN
��z�B�>�;�g^�;d�dv�L�&6D�"�ά��y'��*�b��S=���_'E[X��s�M�31���m�Z��/Wt�"���4QY�����9>W8-i4�;pW1�ɓbYZF+�>tZ�8�`�|f���	kJ��F�?$�4]��f���]��V�+�>\(jE�!�_�P���=��;�CJD���>�;�WL�s�1;N����3>�e'Nr�5%{x�H��|�UW��j}Y�s?wݖx!�3�s����$��tpE�?�����ӛo�乶`��$0r-���T9�K�`#�}�Ҧ\�o�D�k|ptH�!됱W����
/��Zu7f3>o:�d�l~u����a4Z@�s��'6����B��m��+n77ʜ�s�aV 5Cl;�8.U�Ye�վd��2��G�Cn�5� ��E��_^�J�G�������=VÒү�"�sd���I�~��$sm ����3������*�:�-�?� ��h�k?<��*���$E�z|�iJ�z7�8�%ն_N2^ ���'���W�#W4��K���MO�	���-~t8˙�p�:��U�'���2����#0�H�k]>/��
�z�,ʬE%0]�sa%{�V9��(3�~ӏ{��V��n
P�� ]@��:��eL��K�vΤ��8u�x��4Hٵ��7N�4��� ����K�̀�[��@G�h��_�+ ��������<��7_X�?qt\򧽼���A���e-W���;3�>��iW� *�0��D7�8�7����?+��{��l	��
Biz����ԣ��}9e�L<��Y�xۏ�}�9��`�엏����!sC
.�9���~+��@�)\bK���.ti������߾��;���&���>dz����*p�]�1[f7L�z����ī�oa9�0����o�ܢ�Y[�*�H��k~o���r��<�6l윝>rIkH���eɅ�]o�C+��Zwѣ�x�I�0o�z�ef��,_��#m���Qe�Z025��p�Y.n����hX��%�k�g��_6���Sx�l���y�w>CA~�K��I�|�[U�=KC�������z���T�P`:.��w��m�pċ������5?�յ�: -����� 	������m���=+�	�X�ۍ~C��g���{��_�g�-߃�x�VZ��in���Q,0�.��t\�K�]����^�*�63;��%y�g�~���D��u��mIN	�9/�3���Xn��7��8�����vt����w2�!�����/R���֯�NN��C=�{?��W��������?^bi��d����t��6><aC��Q����t��pG���s`�0�����X��M������AY[�K��u����캶ٝ ]�w����/�;8�ej��岿͛�(s���LD6h�hC$�|q���L: q�}vz��I��SiΖ�\2��zf;	�x3��Vw�u1�9A���϶f�I�D��OF�����K�[�r�����?�rD�!����	��{
�08E�줼g^�厀֙3s��=$Qw�րǥ��ꅾ�%XU7�4�����&g����|4��^拫��ͺTg�p|��g���
�����=���J�,���c���ߤ�M;k#e�0��`[q�w�h���gYRz��R���gy0��ǥN:�
�#N/���nO�m+���|D���he��_�u�ѻ���C�}��M���:�/���:udC�����s;�\U��)#C�8�dV����'���F�S6,8ef�I�������ַ4�7m��0���=���e�p�S.]�7���4�S�!\����V���Z"��|�U�ɴL�ut��7nsc�g�o��&�k/��w�1S&�F|"���c~�����Y��1�ڿ�Uy��3�Sz�W����C���K�~^U�h��Iy8�8c2�5���܎�+��i��� l��j�U	|o߳��x��W�=�2���s���<���*��pz�~2�ߦ�y�O���Ptϲ4���Wv�v�l� ��4O����5�q��3A^�x�A��X�v�AЎx��}��������k��1����#����^RK�OC^����{��a�����g&�γ���ˡ���3��FZ�^k˲�U�t�'�g�t>�3ؐ�u`�"m�v��iig�o�l��f��2@����q�uPqj�_�Y"H�%=d�'gE��1�Ɠ�u��c�������8��Kw�ލ�<�TI�� u�saM��@�ٗ��v�
;&���*�Ϊ���8�k{��V�cX�
���H�s4Zv{r�o���$�y�[�E�:�.��u$��{V�J�U���3������A�4>���Ih��;�%��v�!?���n����V�Q�Fց62��`�'�	Ƅ3`�H�M}��<�R��7�ͥiY�$��B�)�����,���G7�s�v��`L�A'm#��%��)p��F�B@��|GM���C�?��,���̊{��֡�L��߾k��w�+;S8����G~����[D6>(/�32*C�'�����p���e���s��OJ�n����ڲ��v���8��@�NR:�x���`�Ю������֛x��]�IhJJ��Fn�1#�3��[�%2�KW�X�����zZ���3e9ԍT��+x�z��A;?�$M���Iܞ��)��W��T|s.�:�:����\^H�tR&���A��K����A������y�)�������a_��}9���$\���}+}�2}�"�̢>��_X}�>쯁? ���������`�yp�3ւ^��O���w���o�y��Sn��t�Sg�j����βy��3������5;W�9��:0jqd�m ��'}1܎<E�Kޖy�|z�}?���g��7ny�+n����(~I�`1P9���|��������O�t�N�;2��V�Kӣlm0����XwXbWhĞeS4���O���9�V��`�X��À��l��16O�^���f]��e�4Znp����)�ݑ@Ȁ�'�ݡV�ȩ�J@5۰��Oi��� KO&X����tfI��t�������Q%3-Y6�=XT��jVJ�ٹ33�gB���1�	["2m`��9��W�<������l��p=x������k3�*Jڸ�D剠�:"����ä�N�yV.`3{�9�pڴ�|���pFg������<��N��X��/=i��-���Й��"ߺL�_rZ��ay;KD����@̀8��[ݤm��O�Uml��PWi _��W.*��@�>���9�7�=���n`�u��>����8d���>�П܉�w�ķ.f�ȯ�Cv�l%����g?���-7���ČwP���e�-m��<�-Fq��~��65*O����E+�O�h�H�s��\�?����g4��I�m}��oJ�RՖ��
�ߣ�8���D��^�>��!�6��Ƞ��"=�{?z�O�O8i{�\�Y`h`=
��,��Ӏ#��hD��l��8�{�(˄Wi)��ʟ��a��+O��W�Ko�M^�[�I���
ֳ��N��oe��Rx�O�q>g�KEo���KYk0v��:�������}��Gߴ?m�eM�Xv�L��`9����3<0�K6��"��n��'Aca���[�����g���KG&��?��������?�cl�C����q����N N��wu�n��Ș��I:{�>��#�qfhI���ڵ��"�~���|g� �9�m�b��0�N|ݎ��ya�<y��ɽ����{��{��߰�mo{���`=@��&/*1P8Bq�[����@�֎]�,�/����̶���ͧ=�����K��W[��r����sw�c�������ɡ�{&|js��xh�"�Z�Ҟ��N,O6�ٌ�6MN������kؕi���M�&�6��=6��q4��b�%��X�#ʜ99=y���7�k�m\φ:^�|���wR':5|dv#N�R-��rF'k��gҥ��DY��v־_�Lr�l8�Bcz��sv�2�aޙ�Sl�������A>H�k�Ó�o�yr�������Q1 ���/KCt��T;��tf���!w�������32.�\Ipᬋ�:�L�dF0�3E?<�UN��A�S��U��'<�Qsx�uh�ȻTqΐp|�e��TV0"=��uR��zs8�0˜��6�Ӷ-�Ao�,I_x�~�;|g�2�w��)gM��6m��ofh�Wynr���g��ɑcG3s�es[~��~:�ܭ�lF>�f��4�'�A�A�̭;e�*�\��x��'<�V�|k4��@ƀ�߶ѭlV�~=8�����v�w�Yt��}pħ駙�b���a�^O�������c'&雎�p�傛i?����7��'>>y9[�k��̬>�\�4+'A��ýɁ:�z��+kUO������:(�Ծ*喉#��0����E�k����AG�����)����Y�^���=[����e�f�U���A.ީ$�ݜ�wr�.�v�Y^��a9��!ӇB�&�Wiy�än��\�=*��/�	�A�Nc�	�	�����{� M��@33믻����Fw��q���I"A�%JK���ٗ}�����]3i^��f;k��c��ՌvW;6:F#��F�AB"@� ����U]�]Y�}���L��V �GwV�������qy���l9�0��|x�Gw}Hߴ�{ %������7-�����e�.��,cN�.�ug�� �]�{�#ðN�Q�����G��??�<Ҋ��t��H�g�-/��̏yL3�_z��[�q�o�Cp��i	~�˟��?F����Q�ޟ���I�g\��*��[\57?3��0�`�,O*KY��5_��TU��W�Ay�C����b��A����T]�� �`�W��ɞxU��\zF�y�C<�q|1�>�b�uϑ#Go����_�r���$W�23�A����?}�����u(㛇�x������������ś��.��}ꩽ���7���L=ti�8���b�Z,�����X���;[c���{�'�O�d�}K�8��0�j�`U��˩�k�TK|5�)��˺�0�'64?�a�z���̎�!��G5�f�[�v cICU�;��4��J�u�@*�����9�Z�l��H5�m+�:��=;�5���~�Kg)�e:|�pq;k*��=z����e�i(9Òۊ�Q����0^�>�[>�CQa�>'	���`4>��a��Sn[&7ϔ��V���GBM;�v*N�F��vVF���"��2ۿ4UD�0є�٫ N���d&f�4�4����p�|k䨛�|����8+:�j`zO�W(y�ҙyj�eYF�3j�uVʰ���Pa�ɻ3A^��:��!�]�x�CwCDx�2����]4�t��l[�2��5�Sv��PsVEŶ�- ��˜9�i�>EA�NY��〇��br�U�ʙlk��k�v�����e͝�G.>����]��Tq�ȑ(��0P�m[Jm
Z(�xӤ|MA��e��
$W��g������}NYoHx�P�eϳ۴w:Qhd�sp�L�8���x��}t��NH&���!�]pK�5�նi�W�<)��rC�4���%/�˗�o��<|&Ļ�+�B�} �5�.��8��g8�rZ��n�AS�lʏ�����k�ؕ'�#{|d�e�.^����Yz��u!��t����~���&eXq�<�[ތw�=~�?�a2qo��b��Y+Bx�.�_�s������}3��:.:�����ߠ?�}�k�j�%t3�{�I�'��z��߮*6]5�bv�s;{�N�x��`�|-����U,���a�~���d'�:~:a�s7_>U@=��ցBʯ�(m� [����訅C���q���o�N���ճ�>�0��n�=�UXsV3���N�~�L�y�'��gn~�����۱s{�;�޻��v�-�֖����>ګ@��z��N��}�{O>��7���O������l�G�}��z��ߨ����~ç�~�5��Ж���TՇº���-S�1�4��4�>π����0F�K�V(23
�YJ�0bX�G�5����6������
}���0�4J��j�%}쒢nT \����YC,�dk�=��K�z��S��v��]�۷��_�\�R���qЯ���*�V��o�_םm:|�pɒ�[�����mgW���Ҡ!�cl����⏥rkk���}{c�'=�K���]Ng���i*
��y�K�B���=��~�,�6Ae;E����:��i��fy
E=~����}�Sc���,��/���Cс��,��ԃ��N,ߕߩ�9�U`���������� �O��T��i��^G�9�~�Wg��A#YZ�^����f�x�a�Ci�>�#:x�*]�T�72T!n���;�;q	�;��)/�NZ(���F���+�Z���w�k�tD�L��^Zİ �� ���s�'����g*ϲ��ݟ:u�����~��>!�/����EHq�;�P�o�S����%��6�p����LZ�䌖�8�����ܡZ��!�%\*W��<�Ɓ@emSz��֭���'Ƀ����@�y�G�Cϱ���KFy���L~˓�!{iˇua�ּ)O�\^Rޠ!�L�2���ێg��~�3����`^���D&/�M|��ֿ8���gZ�ٮ�?�o����i�J������-x����đ�I������q\-o�Mpm��Q˙�������;�	�Y?!i�|�F���}K��m�X=�w��s��9�!��{�I�'��q����M:ϋt���F8�X�EG��n�R�X6������^�|�˝�d}�J]�|c p�WQv�J���e6:n�n��C�S�����A��|𝩋�x���z��ʃ��v���A�,��I����K/��eΚ���?�����u���<]mݶ�8{�l}�����}��>p��gn��L�����e��/���_��?��7�u���ߙ�G���'?�<��8t�kT�G�V{���4�����͇��w�\켶^�Y�f.���٫_�6ا��P� p|���o�%����ptVņ���AG4�S�`�2�1�?8\Ln�^��mEA�-:��S���:r�	�n�q'��U���	���uO�ʲ��T(P&���C�u�CC��rv�A�A���dU���3�r&��9���mqدyš3��J�s�Zy�b����1��@����<0�dj��n�h�@�nyQ	�"dE(�P\�ok^&+�*�7�y����&ӥ/MD����w���?e%�˯��rrO�ƙ=��Fd2��+��A_�'+�b�Tƾ�Ki!�w0��a�d���/��J�r�W'��f�ٙ&�Zcؼ���c�-�(g.x��}�_�+��,�k4}As ��KU�t�Nѹ�>g8��RɎ��f���B(r�=.if��=}e$@�����:��Z���g�X}�+���[�p;���ҷ�,�_�+,��=ee5�/�̶�q����h�i>���e���@Z\��1c�+i�^�2�n ��&�"&hE~F�U^֑A\>w���>��h���5�W�/������w��]8��)��<���[�LO�	��J=�<�r�"�<�t��x|��&�$�AOX�r��?���LZ�^��82iX��G��4�hȴ��|�����+}.i�@�x3���<���-�_�|���Ӡ�/�n��im�ˋ8-���7���?���bO�/~���c�瀟��ޟ�z�@K�g\�-�%�i�����`_���4���1��:C@� ��q6��4Qb��웛/�t�v�ѩ��c�&�
YV�f�J���4��y4T
��_�Ur谣N����r�'Nv���S��������;�����^�?P"��s���ַ����O>��^x��q9�Q֣[�UK�+믽�V��s�i6�2�]\��c��v�y_�_�Q�w�a���|���}��S��C���c?Y�v��ͥ���ۊ��7��գ����z�g�.�/��7=���ط�8��N==;Wq,.�J1�@;��{ܐ���2U�T.���s�u���˞��27��i��h�����õ��(�8�pL��cIZ�l��J~���莡����/��3C'O�`}N��D���./*�ֵ,�a�a ��g�`�+f�4&�����,�V[��0�I��$��h3>�>l���P֢9+M����OC�6i;�Nh� ����g�Z����[����>�C�6/��I��9�
���i����:e��Î0R5b�;��M�FC�r��ф��]4ɛ`Rc�P�,���i�)�<�'>�y�������Jg!�Al���0�4�,�t���cF�(.���GCQk���(_#�h��D
� G���(jfi��:��< x��jg[U�Æw������]"���d�`��iXq80m���9�R9o��2�ef��������9\�/�}����k�������53�Ay��UJ���
�m�UP)�{�X��͓�c�Y��鹭r�x���������e�;G���V��7��q�O��>#{zW��h�߉�x}��&2�v���%��m�l��K��vnے>W�Y��a"�r����e���n�y���KZ����q��>)?�G�/^��B��,��N���h�+N��O���=̅l�Cz�� �.<�w.��}/�~�5�����x	�Hj��~�W<�%~��N�.��/=e��?��M?����G�i�W�d����s~�=�
!�BO?
h{�f��y��/�<Ǘ��p��G^y������33�>g2�{�c^^F��(
���ƕC>����n��Xޤ�7��l�����3��v w�m��Ƌ�2��%�[XB�}F	\G9�<�W�>�~���|��뮻�w9��E�bg�g�w0��}����}�;�QΏ��bG�L��-�Pz]���3�j8����@a����g(��o�����~uF���Ϟ7N������~�ŧ���λ����{��=ۊE4�m��/|��b��k�'��o'��D��}�Lqb���Ł�>^�޻�:5����b�jK��=�S�h쵪����>�Q���˻���,a�-Z�"ʤƊL�k8� bf�͘M0��#g*mڱ�<;�"�Al���lR�~��`B�*�|�ֳ�?�Ӊ~�ig����a�����Ƙ�����0�,�m�<Κ�[&�_޼��������f`�0��Ԙ _(N�β�~����L�*^�ȣ��C�<6J�i�_��)max%�x�G�ȿm�!���K�|6�WC��W�ViL�u7f�L�<p�R>��0��o0�F�0ȡ5�4r����cǎx�����}K��0n��u�WCz���8F�c��bv��922����Lf�8X\�%�]�K�͙,i�Ƣ_���_ִ���04Je��Y�k�����������'��O����y5���YGU�����j���w³����s����[����?�l�ri���W�Zy���'4�C��m���AT�,'�P���	<�Oċːqzϸr��'�m�%r��o��V�X>��.�{���62U�MyX�泞�������]�8y�|4�G|,�uH|(�-�̓�G�-�;�ŕ�E1Mxs�w�e�ķ�i��3�ƥ���iuÚ'��,��/����ƢrK��:��u�侪���}��#��Y��%�oD]9O���]�ڸLG����۶��q�Wۍ4r��g���|A醆�O������Y�~���O�D��-\ ���I�'��z��߲:��֙�?��|ua��]�}���c�&�q��B䞧��&]��W��X��q��1;X;t�Z��rʔ
��p؋A�N�,f(\���)��r�7xWV>�K�tq���Z����#�b��`z��i6�~��}�&�������7��ѧ�z��S�N���N��:�?�hwTB��*.\8�y�WWQt�l߱����w�/m�4�{Հ@�L�ll����3ǿ�����G�}��>���>��O�n����|�tG �[��m�ٹ��/V�{��wo=�[��:�ƹ`Ͻ^�9=��������_��:���C�A��W��	�!�я}+%g]��m��Ie9�xzc�_,70f\N9���(��S�Z�������QA��҄��xl����W:PX�k��Sg1��d����UC�nv*�
�Kլ3�afݩ|X��1܁; �.Š��!/.Pr�E�¯�zjk�Zl�*�T~5.��-�L?�.T ���ź����s(Z���~�5^>�#�{�뫮����@B|�SE")�.n��!'��I֢|�#�iV/��Y.��Fa�e�}S���#���ʪ��L��,����=\�s�n�w)Z���X񎱤���l�Ҳ�b�5s�k��c�e(������'y M��2�<)#����/J��6h��-�)��T#9�3�u�׺�����7h��n��#��[f5�Yg���e�ï���>@Ώð�!�8�H�<��������OT�?p��p}���J�K�Y�ͬJ~�?��`>�^���1�2�����m��9�5�<4Ddh .�nZ�����͏&�E4Ƙ�HY*7y����.�qM����L�tI�H�gӉ�y#k�#��=ɱ-�@�p�|^��Y�^�f��iֻ�2>�	Q��Q5����,�('�-MaR�(�mzo��ۙ�L�H�N�!���y��*���=�����n2�V��Ắ�c��y�I�3o��<Ֆ�빅O�	\��~8Ѹ�R�m������U�>�Uf�W����������w�=�e�ZL�Г@Ox	���*��[���cc�E���'�}����o�����3��
%&��� �N��D����� � b竒�fbЧ����4:���Qf�7�v��tE^�;�:Hy��71;k��H�ge�(�o�r���;Μ9�s�޹���)���(�S
×.�����w���x`�X�c�%Z�h�{�U��͊ٚ><"�����^8z���S���sK!V7Ƽ��e�hoKkk��.������~������?3��,�6V;��.�0p�N_g���y��Z=���}��zlb�z�%K�~�����Ǌ�gf�����+�šO�WؾW�|�'�NPf�8�´7�#�x`�\�8uG�U?e�`ph0u�����Js��)	�/��0�CYg��C�^�2�{7�PC�TM�mxȥ~�F
���Y�P�\���u�r�=��&4��w��mmݺc*��1�03+*�33�°b�`�%�r�6����u5����d�M��f4m?�i�1+F��gӺC�i~��0���c(��]�i�QN� ʃF�������Q83�	Ȁ�k�(�F�ʌyY�|��e|�	CL�J�a���_�S�������F��3Y���t�ag3�c0ɯ�y�3���rX��3��r��uf�U�\ڔ�3��f%�PBD�p�t+��j�ʋ��r�_���$4��Kaݎo��e�<�w�^A=H.��{4� ��XDQo�[���Z��hg=�P���>�g�����A�L9,�x��_�*��(H��a�e��m7]!�!\���"����p&�Z��h6B�	<ևy�7�T�Ǡ�����j 6x�]6m�1�l3���U�	�U�<H��K��
���ֿ�L?�K�/�)=hX^�q�2�yB��b�wk�d|�E"�#n/��$M�(k�Hr	~şh�x�	WN'�!;�5�z0C�+��}F1.���s��E>�K4�A��5���Nl�Qi�_:ޥ�C���`��"g���-��� U3����?�I�,OW��K�Ò�}�9޻?fI���O��Y�x�ޏ�z� K�km���o��K���˿��+|ɽ|;���ҝo��N_��:�8K]4;�9۔?|�	���ɫ�с��1z����	;���A���X�dO[(����s)�|�_��R�*�䳎����|t�k�\ZZb9�KSSw��-|����յ�|���{�{����/N�h�A�m[���?j7j���9����M�_�F���k^������y�{����qv"X��=��V��$��"�ۗ����}��?~b���������t�)/�O���/��o�-,�n�2峊'������r��=��v]�9�Y�'_z��/ף�������:F{Z��,�^���0����#�Ln���C�A>.���E�@`�,G8t-^�,�!��5J<{[�Q<�V,�a�a���Q��4X��K�o�>�yY�,�$�Q��d<�� 걩�f٠�wR�C������j1��>�� �^�R>m�3�n[ضm����"Mz��>�N�Q�˥"BTcxX�|���N}4k#�O��̊�y�g�ϖ�4g����Y7/i�����x,�FKc��1�˙�M�R���(p��F<�[�X�#�i)��K�  @ IDATq�WJ�4���,��Cci>�5�o��Ӹ2?uKy+�ڔ.d�Y����ϴruIz���<�[�V<��z��ȅ(�>��z^����SXye�{��6)#QQ��~��,ڕg%ɷ��l�=0�g[���~�����0�=��ٹ9��RF�]�W�����C���b��ug6ӗ��ȏ|[�>K7��>!������?�K�Y��0��|�W��o��k���|�'����P\���9N���G��^5���m��,�������x
��' �����z����,�l��͇���!r����?��3��pl�[+}Ox����\�s9�8��8s��3^p]����9d9%�
"��D#�[۴���Ee���δ�W���6_�v.?7�^�e{ )�y�L�8������i����r��CW˫��\W��Ϻ֨��K�n�_���+�c�-/�`7���N�>�N��{���7�|���>��3g��{�I�GB�h�#���I;Y�\_��w�m����D�]�U�>Ϭ �x��B����>������,�Q챢�u���E�ۯ��``��Pi��`�����c1<�׸�qK7/GA��T)ҥ��W^~� {��Q�יŨ�.Ou�x���,¢^����%�T c|�� �zl��Т�����{q�0<2z˱�'6^x���p�}��w�ݷgǵ�sS��=�ʞ��u䓷�۹������*pD.��Z^(X�ĸ�xX�]���i���p���}��7��2R��ïV;N�)v���G���Oή;?�^��~[�e��塨�pΓ�%����l�ɞ�>��Z>v��m`y-m,Gݰ�&f(����(o��¥^�N���d�f����:.�c�,8O˳�t�<���L̊ƌKx��$�;i�}5�.ҌӮpT�RlP)�8PA�����D^�����̎N3�c��/}�����G}2�8:�6��<?�'�[�����?�'��l�mڻ0��l0ݶo�,�%�V;%}�W,1��(y�5ʬ!�ac�-Ų;�N�(����ku3��8��3�ΰ�[�L�=DI�t��xg��P��t�[xil�R*LSS�#��a«��S���=l.�����<��?�h�[GI�R)g�69�MY����j5��/?�L�tk���)0w*�x�laxp�eX��%��ٹf���#�R8�XY[��:�Ξ�z���K?���_|����1r/�����T,��P�#}y�,F�:߶# ��i��M���)p�xSZ�-�縀�~�C�W#?��M�i��۶*�O��j��SK߲�z�Y�X~B�%:M���wӒ�M곑A��������-��2=d~�/��#hxE�R�d|/L��~}�C�d<�"�w��J?�\�'�4�-����CT�G��邉���J�>�|)-�S��oYRy�.�������]z)]<�۸RZ'>B�V���[�C���2����1vGy��bF�I���|��]���bp�	���)T�w�I�'��z��E��i:]������e�
� _wc鍊$S(��%�Y�H�>ub}����#�����,�!�G�O������dC�A�.)��ۯ��@	>�T�� o*����|͟����
�|��p�� h�y�T�=��R�FcY� AY+>\����:l�-ffg���x�f�t_����O�?wq�Ж���SǪg�y~����}?�3�fc^]�XL�0�1�c[�-�;3V+���}k8��;���t}��n���}�M����\�4�)N����OT;���l����b����~���f_1����9fs�9�j�e`�.(�`Fָ�����A��9��Q�$֋3S!0�j�f�X�)6�7��MJ���1;B��b�s� o�+o��!���r4��:��]���N��P�T̼�O��aP��;��6¬����'ڍ��u%�E�<�7���-5�q�M�����^S�VQ����T��W��'���,�^�[ے4��*a�a�T`��(r鞳I�R��_��D�$�'ih	'�!:!?�KD�TCHy��)�c/��7Mͫ|u�.]�F�btlK�kװJ,�G��Y��ĝeh�)���BqpՃC4����3y��\~��r���w����\��"<..��4g_����Om���+�y��R&�A��C��e�z	�螝�����e�-���+?�����������i�ϋ/��Uu�!���e}��)KԿ9���3���@w��~�y�;t��o�������� �|��Ms����m�9�\)���8m��B��t�m�%-��e�>3�RnO����m��S���w�g�GZЋ��O�_��z��x��yz�����i��
gz�-�-�t	��n���Oy�3_�9��	�y��և���B/���2���{����޶�Uy2\���r薅I�0iH_�����M����I��y���w]g=q43�5Go��v�k,q�C�g�r�w�I�'������������_�O�r;������8r䭑�G���0uU�l���_~��ott<?/�x:�|C�/�{XP;w;i/;p:n��3]�Үr�}e�x#�U�T]���;z;x�u���¦�v��Q�D��d:K�R�8X��a��[��p��]�K|'ǸҰB���ŧ>���u���-[7�9��L���7���e���;��}����o~�Y�JlT�̠�p���֡��ckhM��m�ξ����@�ml�Ek"�s�J8.G��;�+ X�q�T�15Wl��/\*.��b��e�֢�D1�WE�ř˱����/\����9a8��EK�C���ff�p�Y�/�5�`�Us����1�J�"�.��X*��PV�a�Z�8a�]O�֛��`�2�%nQ�[2��k�b���J���Y��"a��^l�;`�qH�F�uJ���F^�(����?�p�4�H����YN�{�����Ls��϶I�K����b�2R��ݱD5Δ�6n����,�����������Ò��h��&/����$-gd|74��!=��'F�^g��k�I�8��C�K���G#K�0a)���
[yG԰�=>ڌ3O^�r�:2�m$�O�2s�,�~�����=c_�0mQ�#��:�hC�B_����f},/2�Zs�e�we��ߖy����^��a�f��
���].�����_�r��'8f���:���>J�����#�Y�ӣ��bk�yOr�t�F@w�F�n���n�pQv˓ww��h7.�]�\�����W8a��3ۻ��x�����+=p����f�J�9������L\����$[�����y��y��8i�s���ϸ̟C«p�����m2p�x�P[��_���.�4���"����9����o�\Q~��o�u_m��e�pݗ�-�y3���w0��ۇ�/�w�'Oз�1�o��~�B�o��Vɇ�?Ã���ꑯӇ�0^d���I�'�9	�f�~UƢ�ͅ��w.]���/�t�~�
��>�% �U���Φf�E:�|U�*N~e�æ����v�e�(�
k~;t�P��5�@��猁Az8�kf	H�Y,�@�7�u{� �y]�M�gy�p9B�l>�N�/Pj�T'O�*N�>ͬ�˲&��F�b�l�í�0J�Յbbx�z�׋o~�k����M��L���;�q�qQ�����
"�_]�ͬ�k�0|��}��\�0���kv�~�s�k����o�7N�K�ѽ|�xku�x�}|��zd�n�[pv��R�?�G=�b�[?��(��Th��DP{ӳ���A�[Ƈq���G�J��!��?�2FƌF�R1�����Y���=P�o��O����0��8ə�M�v��4��Խiֿ��P�+��a}��h�s��zV�0�_��v���cY�xD7���|��L�0~�{�m3)Ѯ��t�/��a���&f�l�Љ�#�m�^.T1!Ĭ�p旧l,_����������e6�\�#n+�pJAZ�7��u�1�o��]���
��L�����B��(i �',PW����~�L-�<�|��QN��|�sV�:����q:��F#K8��?\Z���|���F�:o��OC61IyF��2B��i�K�F���L,��jhK�>�6u����/|����D�9��Y.(���1����x�<����� ��GQڼFMZc��O��)>�e�W`�|���G����o�V^�ogxl�0�S&޻�rU�W��Ƀwa��4��C��<,"!�t� ݹ���H#)� J�t���%-�)K-�H�Ұ�������Ώs�3�L�w�mhA��O�	ɶrE#r���d��d�!�3�'���eX�5xB����C�Ts�x9�?�\D�K��i��r$�m�<����K�i4�/�w�ӝ6���u���`4���Yܓ�SA��5��Y��#���;�W㯕�{���wL]�.����VF$����K/��G����<�z�K&ށ�YU�I���:�T~El!��������׭R߮�*�[��XyR9�����Վ����U�s��)Kr���v�_%��%xj����|��~5T�U��QF���U�W�{zA��EN�?p[�� ��)�;#���|,��TEe��&~D�k{��7�u�N(����$�nIrl�b��?�����/�<�p	>�����[�H4��A��Z�'0��w�Aq���j�\C��hi�~MMc�r�������F�����uVoO9ϟ׊!nf��9`��n����豮��W�&�����d��6d ���VO�n�;nH�>�Al�j= �Mq[�����ƃ�i|�_ө��&�x�+½#�*��u�mb)��:7�gY*dC�ǳ��݄ *'���v������Q�x�y6��n^ xnpR�������3�:9�7�������v'J?.��=�+-���?u2>��#�r.ˢ6�A_%�<tӽ|�&���p�`�z�6�|.��ż���\��)&v��T��Md��|�gbN��Nԝ�����#���cÁ����خ���l�a��M����l���!���K�d���#)����"Sl��&�dh��yB&���y�5�{���ӷ��o�T�����6��g�7�)~�>��/-O�3=�lk��,@iÑJ<����1���flB��T=DT�d�������2���d��B�^Tf0HJH���n�$�˯��1ɖ�5S��1ieL�~:a�#��N�!RTJFO�Od�����bTH�4��eߕ��̹d{
�d{�J���a���%2W�ka�qS�f(5�He��v�{�6�X��+�J'���k���E5Jp���}�1jʹ���9Y�4Eq�rs��x�¨�5L��cd�I/����Y�V�z`)�T$t���a�^��w��)vߕ�����}
QA;J�}���N�������A���5�fY��7Wm�>�	�k�v��"bf�LD�:[��ɒNgig����h��K�>�w�<����n�L���6�nE�W�L�[@�������!5��EӼ�rZ�/��X :�>*N�V�}.���|��\�ː��gG�� �����HaM����/��H2t��7�u��n�ȅ�<7�o��|~!Bi_C���bϼ7L�ԝ�"5ɣ���mB�h�	
݅uz�[v��M?��#��7WKKG�U6Y���+�͇�MnrӀ�m͆�������y�Um���n��77�)�X⥯D�L��R��Hs侢no�=��T��u��^�����Dx��*�O|ʒp��ֳx��;M���G�.��M�ba��aҐ�Ogp/F�Ч� F�.��o��ayc�>�ś��߯��y�L�^߶1<�$�)%���@\�F�C�҃�9V��j����J�tǟ/��S���۾+~�"o`���C�,
�q'M�{&e���k�*��#l6-�����*'bUm�εyc"�����~P�~Q���ʖ�`�X*�7�MI�R�AK1v��;�D�Sz�"�Ñ��|w`�df
A3��D��k�#���8��H��9٠E��j�ѓ ���,V��Q�0�˒fr����o>���kyfN��Fj<}p�^�p���;m�c�l��M#C
��RR]��4cN�"SWի��ڸ><���#ҳ����7Ze����7_�2�do-��m�N��K^&�8Q�w􇆐�nb{�V_g#��l��ɮ#�^O�|�ߢS�Qv��$��r��j����;��Idv��o4"��a�u��j�\Ϫ|*>�݃m׮{]��؆��fAz��B��A��=��<?d´\n�팘����>�U7���Խy���;F	�q��`Ɲ��Hꮞ��b�G{&y�"2��G#�b�`J~7�~Ϥ��P�N��[�KPH
�)į?bU'����᧫?�x@�tR:}aA�������z�s���E8�s�z�h"���/�ͷ�r��;��K�ir|b���x]�rR�|�\d�aai��a�G+��kE�,y�8� �h�XM,�
z�c��[;��;�fH��A�����*$h�!ǅÅG)�?��. ���z� GD4A��U �H�GK1�7�È�-݉EM��f!�#?>4c&{0 ����ϲ�]�O�-��3{U������8�Mx��B�'-��akZN`���E;;��]��iw��"�����#Tdsy��
!��M��Jׄvd��ii�x���{�g�@_�!���_ݏ�iny��3Tu�$�Ԏh�h��y�K��[0�=�'
�^7�S����w�C��[��G�� a�gC6�2sRƆo׺[�h��d�|4^"W������L��4��R첾(��í%��D��b&+&4���{D��C۱�r<�܀"}Z*p[>Lx���>��kA�!^���7��_m�2^�궯����H����.BdO�tL'ߧ��. �ɲ��/�:"*��`�<�SD��r�y.Gz+�ƃ's2�94^Ǐi�ؔ�	zo)� ��o�j$w~���E��U��w��0�41M��]��f���'ְmԟ���*�,��Yp��tn��
D��Q�ݳ�jgv�
��Vo� |����x��1;dl���O���D���a��-�tڢ��N3�˲LR(I�ÆЙ˓�c
�?#�ȇ]~Ji���l�����{����^��
�|��R�y��m��e^zS����	ό:x�>]���ܚ\�_fg����ܮz�ک��ǘ���_�(�񂝰�p1�Q��ΣX��Q�A3-�Am�l<�l`����ϗ��>�O��z�VXæ�"jp{ �࿽3�:8�4<	���#��ר���{���W��f�;��v����"[&�����o��C~=컀ܢqH����7����������oҜH%@/w�M���.�4�����4���M��n��֡��,����p��|�2�&z^�W�c1�KM����E��f9c�#���q�)�4;B����7�tb'�"o������"r��Ԝ@�K[�[���'{ ��9��b������d�
�s���<�p���'������iy��?��o5�Q�	)��Ϧ�<{�M�Y&�4�9k��>#����C�8d��.yX�[�Aω�$F�h�3 I�Yt���8tD��.,[�XT>`k��	�B�Ҵuf-�I��(�==H,3�l�o�7�@ة�8�@s.�c�o�����7�hW�,��CJqSc�O"/�Ds���ܭs�p�}N[p �jJ���pץs��Z4�����hz�J��ŭL��eu�!�y1�J�"�l���}�� ~|Y�Ov�K�:�n[#�ȭQGL �(�)����ܵG�k����D�gxўҹ3��~_{N�q��β!w�T���k��ؗ��|���<��%��������e�[���3���/Iؿ�H��5�HB�}�k+��LVf��~���=�A���*h��������<IW<C�o�'����'��'��ۏo�ï�뾠���L	�W���L������ѦO{f�6�д���d���_�$O�<�a4\����P�3ݥS3��YE��A\R��n���쥰
�H�� a�5v�A�;���"X�ݏ5Em�9���8$��C���yP�m�g�gu����c�T���,�jF�D�O�9��M�?����1w��y�9���6��e}�L����C7m|t�Z�u0A�o.�7�<��\1�c'�@.2��}���g'�S��L��W��jR�9c+d�'��Y�S`/3��S�<Q�tG��$�/�0��ԻW���.V:vH#��]�� )EmT��{�A��!B�<c�3I��&1������J��=9��d�qWZ���e��e�.��,�6KS����R�8i?z_�t/�������Q��VmX�o�^h*����x����e&�7���Aѽ���R��ұ���m���r�}:x��y8��+_�B��ȣ�����'��?����^�а�&2j�=GR��oFme���03��-{��cLa�ݙyr�6��,�p��l�-�T$�9��n����un$V����!D���
�z�A���9�di�9��o�0o�'�Po�S�b��G�Yr��7�w3�~yD~�/`NW�x�9�D�'�q�j�{��ն�3�'i$��X����Vv�ZR��7��ԣ�Z]�ȕ����_ �|�EҦ��*UR�G��촢䣶?�8'�+��.5�f��4�w[�`@,:?`
�vmQ�~��Xʬ.yo��0�c�q�q�G��m*k �N��rE��=�	�`ZQ�&uj�E��b��R�6�p&����]��'��/�K��b�9+��G:��~t"-�}\�Ob���0vS_����Q�"X+�Aa��L����	>R� %����Ī����׻L%Z���,v薇�]�,N��×�mZsǦ�V�aB{\&;J��Ƕ���VY�J���g�y{�9����
�7v�i�at��j�k�3.ǩ"DP�	���jR5o���j�*�Ag��f)��p3xT�OsN����0	�0�߻��].��7Տ�����&�hi�9���o�������|�. ʅ�ɴ�bI��Y��Ő�l#���ţ
�9�<�-���a�#�����f�yM�(��{�E\kN�jV����&D��L�d���Ĩ�3Aq����3��"�A�|��K�D�4(J���p�9���m K[�՚��8�b"��Mo3/��_�^39yL1^fE��۷8��_t��体������(wK���?��<��{����-��no?5��B<C�	�w(ҍ�!��#?5 mϒW5�c�����N_��^�����Zd�a���Z�����>ȶ�?��������y�-�o'����r]�Mb{�2�������	��R�E��s@���w�&��P�(��O�(P�L�
������ ��"�<~З�M�k�C�|*>��K}ۃc��]��n����z@wWR���ŋ���\$cV�l��w������e��~��F��f:K��%��9.I0}�e/�T��$`�Vexce�Pl��߿c�����i_�&
�:�4r����nq+�6����a�e��C�n���)%*T�
��
pEe4�=!�;d�;Ap������q,�OZ����_�F\Xy�Q�������u��3
��aE��ue���)����S􃿝��Ŵ�G�Q��vpc�k6��1֣�~��Bi
xYx�N�V,�	�j���QE�v�,��\�*��ҍ�Jh/R��Ww�Iw��(��ѧ��,�!5��
hY����i�@L�?-���]�O���[-��������;�����6!�V����;s�t!My
2��6�(jS�׭�P��q6褡�]���^h>�Q�@�ց_K��])/5,{l�V>B��z#=_�������~I�]�V�]T]�Fl;JA?<%H�G�������Tw����o�@$ݺ��q]���ne�U�S��z0�&��p���2��*g��Pנ�I�Pܠ6��ӭ���~FMS�>����ܧ�r��9t��,6t�e�|��8����~x�̕���PÍ�خ�zLarS1Z�����biĐmC#��X����lH��b3��ך��4��B�M��2Z>��	U��1g�T
�DG��a\+�;��^��&��v��=+�8xl2��Ԭ3k�A����mP1�yf��ݶ�4��e��*k�K�afڒ��m-��'�]!?��h5�MB���غ�F�r0%�s���i�*z��Lػ� ]_��O�H�ɺ��2�|j�e_�m��l�8cҢ���~x/���j<��qP�~8#p�j�{�Q�����R5sxք�|��_l���ꞎ� KauIjN˝�KSFnW?nO�����������eN}耴5/��^rs�����A-Ȧ}Ɗ��<<�r sϝ��)��".0��Ť���FO��š��JIE�:p��$-��0�ԗ�`X�����DI��ı�U�@�F��}C��R�Όٮ��9(�|0�v��I���	���&\�2��&���G;y��v�2�U�V��o6���t�z��`xraV6ߋ����(�Kh:ɶ��փDŝ����$)��&��~!���vax��Voy?�D�\-�?�׉���W~s�-!�$����H��C�����bF�[͘u떷M�6"�b������ �t�:����I�xll������od��V�L*&	x�6�`B-L>�,+s~Z��'�CФ\)ϡh6+_$�Mm�%�*�q^P���5�.S�M��1��WP��{�հ�j5�{Un_�r���8/|6�H�Jgh3�y5	�0s�����jtwC5V5�kL_��B���>[8c�L��1~�Z�?��j��-}�ԈU ?x����R��t?�����g����'�x�ЏC׼�4�m��߷�.H` XS�PCVY'6ssM§q��xښ	!���ܸ�ЇWK)M{S�S�m�����i'��ʰ&��T�bhm
><>�b�{�����v�H�^@����b�'���۞�l}H�豼��A�]bYɚi�J�!�X#G�r�.��Ѩ�EP�[�
I�-,ȯ�ߍ�vw�y�ˉ]w�:�Fa���2V|�Ͳ���x��jg=�Wo�����\�`q^6_�3��$��O���^?���2��sj�)���#}T�ZB��j���H��sv3(��]��7ٌ̬ëz�`ܫ��ݽ�?����/�a�M"Y�{u�F��Lױ}�]z0�)( ����۱�
~����L���ܯ�\8�0�� ���얁�׮����.��	D�7��U�0I�����&��9>g�B��O�ա�`M��_�}���,�j6Q��5��8�t]�hy���z���u,Z�)���j�:�D���s�I�s�7x���m�ؑB͵�!��>>�!�v�^,���q�C���n^��4��c�*�AP�r;e�����8��54�roi#%�\�ߘ�q�:��l�s�7����?�*n�����I��+Ϋ-N6��m��6�@D�\�E/�}�&$m�!B�������z3��m�<��j�$�w7B�>���m�Z5]�Ť�mXi4�ħ���S`XI�|Gֿ�X��G�����>bM��P��A4���)�)*��lll�zc����,�$�,;#�9�	m#
��Z���&���	s!�/43&p$T2��0���x���Zyn��)8	<�L�a�<�9{�՜�����;�2	���*������ު��p�t��C�dsK'�+��7��na���B2�2A�F����`�LC�@�LvH�D��)�H�MC�����K%�+v�ɘ�y��.���nl�얝����N�h�c<`v䲂S��<�fĒ� o2�q[*�S�蝭����<��߹ٝ�B�	!��w�G���y�r+.����8\O��wp���oT?Eac����A���.�Lq�	�6�S~�����U럶��x,	�vd�(������y��],���׍�(~D[�����mtxHv���ac��ّ|'�{�O7lh"g҃���Of̃��pS��[��^B���A����1���rY.Fls�=�Sɥ�� �+�6�\lT��c	��0���g�kH��!�M�Gt1(It�/��t"��->��O!��՘�J�%J�~�M��|DO�J�[�1�
:���m�z7�
�tއ��N �;Q ����*Hβ�v^_�Fa�B�p׫�79�c^M�8R�B�.�9��,��������1'��W�����wr[�r1]�~�,#�c�k����1A���&�!]lW+��GQSb��@
�Z\�.U+����Jl���I&yYWQ1����k��]Ă��~F�7 �F��b12Y���jf@�����&Y�A?ȷ�m0r���S��%��Ut�)��42�p��0w��� /y�j/ުM��缸���.w��>��J��5d[��Ԗm��iQ�(L�'�#��\*0�}����P�hh�\o���6�F}w'J��,A��"�)2�,�d�k�{mZ~�g_;FW*GU���_ݺΉ{Cf��a�d;[�ab�k=���%��4���X���ÿiz^��$�H��
���%�_U�v�.�VAak���.%�!�Q_²��e	G�*�c�G�;-�/K�@55�j�%�c�qu��&ҥ:�u�p<��"8zޯ�,�RAr�t��ѭ�c�h���[%���Dr�tc���jt�$Z�<��*7��P
[yyCʏ|������W��U��C�@Г�L�ɪ\��=�ljmgP"�/P��SonV!Ŝz�l�v�.a �]����R�mS:�?b$���jްiP��3��e���z $PIp�
��}/���
��6H�4嶈�ڭ�\�a� �/�2E�ӷ�)�x�� K� �9W]N���޳����8�h-�X�)I9�.GN�D?E�?L=�8(CG�h��[%[;�������㭟͢�o}�O\$PΓ=X���)m�2��W�k��t{�}��$u6?���c�T�J|!��%p��.�[���ۗ�L�EEs!W8���d�Sh\Wp<I�����q��OW�7��R��^X�g�qO��8��fC'xſ�c9�Vې���Fo��30X>1��("�46"�y��T��� ��m�s�V�WG��ӈ�fg��	�z=���.L���;b1'Ů3+{�+%0C�5���s��]�+�/k����"SB��K7�#�ݭ����Ѥ���ݭ��!�e����lP��|�Y�����F�*Hă�R�p�n���L�0��_:lk��^���)~:,���i��m��_D�r;sFq#�1�����w���sJҚ��;~��>�Bҁ����w����)B�y��������hl�d4���dJW����?�r�v�q�{�̸{��6:U�i����,-7k-;��~m��v���C@y�
X�9���ic����Y���9U]2V>�Uqv�ρ�G�0�%Ɯ��Mn���P�������ȯ��6i�}-�m��E��/!�1��k>B\"��/���+~�>�����o���3�~�f�2巊as+�*-�����;;�ȷ�M#d��9�*.`?���O3��6�
��+}�����I<sy��}6 ����Z�Č�m;�s<�EŲm@�L��<55֜H4M;�|�Ձ~><U#f(c�ώ^�_�R��;\�������J�b[+,X��9�(N1�~{Ue�K���eE�
��}*Ս4b֧��\|ɯ(_.L��t�Ij�-�D�쀜D(��$��-���S���e(�b��sV���\�H�!�ϹU�A�l��NV�Vw�B_��:
�L�|�Jթ��;���T�|�G*��i�f%N�<f0H�z�cM	���_	m<�Sޞ߹d^��i���dv������������X�ps���:R�F`��3��L>�����O�Y1�+��S�{�nI7�5�^�G4|g��=^�����+�,ۯ��p�_W�2���숭m���z��K<i���۔�2�Ռ�}���<�M|(��+L�2���b��nwb�P��D���z����]łH<�ywÕ��)wj9��$X.��y%����o�Jl06U۸�kw,���Z��$aq���-k���������,R���%kI�+Ex��,7�-U:�I��89�yz��i>�	?�@��%�%m�?b���f��e�c��=�;�~]t�p-�e���L)��=��St@Ѣ��k-~ͩ<D/�����ozo�Yp6���Hs�gc�+Y�KQ�ɣD�d6�����îQ�X���>������<�L��];�;���Tɍ`�-�z��zq��vc|z�Ϲ&��wq�;OJ2&�=S;�-]���.�ݔ̇kk:��:�j[��sa�
 �Z�<�E��W�;�v��K3�V1J�'u�]�zI��R!�,]c�S��� �t)��+��CëO�X~��t��oxnXi���5�K_�J�cTD����&;�Y��������� ��^��)?O�����i(�~�L�Nu�G����i��1[��P��£�Ғ�$i2
��^&YM����bS{5bGʹRpm���	DL���t��L=�P�r��C�����F�[m��v�(?�����h��b�x!���ˊ����#��u������9M��[�%U�"���"g�"R�^'�@����t+Ǡ�E{H �V�pT�	��z�0ܚ���J�WV �8�6i��<	�=�wA�����B-�9����0��'^��X���#��2�_K��S;^�ǵbH�؆��0��1)2E��B�H A_��5}�ӯ?v�UP�N �������zErn|SA���U���piLi+��*�f'@ME:�D]���4�7$}�Q��E��Ƽ9�c�G�=��d�{�M�m�1����wC�<.�WT��^���O��	�ӍqJ�,f)p�"��^���k⮑g�V=���)u^��xČ���X	V�n�e��8p�����/���b��h�Z�|^p\�<��O�\��|V�����l�9�)ҕ��Q(�	����P�0���{���̮����9H�F����֬�j�Tō���,��rQ�w���+�a����Y�'�X}�b��?�?
C���*Ɏ���x!��Fc���B���,����{���<�]2ފu��]6�Ў!R	�eo=��(��W67���8�&>��v�i����>�>ab�D�UK}�N�a�S�W��}c��M�<�\��\�g�Q8�ߑu<E�4�Ie����T9۔	�����h4<���2
��@DY�����ʉ(�U�'�X�.����#�����k�5��XaS��$Z��-?����J\��8�١�������3��;7�W�I�j�]���Y0%����-ScwP���7s9��Yv�n�,�M�o�uJn�=6�]v޴������!f���B�`���r��˰���_:ʔ̜����� a�1�|W����4�c`��~�9�=Qy������VˉY�?e)�3��C�������8�2�0:{J��Ҽ����"�(�m����
��5�.�9�}> �4}��L+���1�	�O.�vehE�q���Y6��V#E^Ex+�	9�����4rm����-p��_�%;�r'Sp{��k�{��ۓS�O�a��RA%^_*�=;�FQ1έ��K�y맬]YnǛ��}h�Ń2�7�Ǚ��J����|��I,�H܃�f�{Dd���#�h�c�gA�;��j8j�jve2[�M����6�0��c��h�+4��4,�:�&�"���C�$�Yf� �Ϊ���Pe���/N�us~�yKU�ݗR�RD*H��`�� :S�	�7.��G=1��p7�NK͑�ɭ!&��=�r\���?Kr�z��^+�L݅��ŲM�G��M��/���)���h�sۅ�pK��Q���E��*/�tV>��xY.�>F�y<^��I����ǟu�����̰G�h����U�&�����-��z�����Hܤo���8�/���] �t7A=�#������ˇ:�U�Ủ��co����w����X��e��IX�fl�/xVZ��g_́���4�X2ˤUG�3~���sԛ%�E����ĺ��T�~f�Ά1-�i-��e�����3�h7��x�2�W�����i����+���>ڊ��w����~]�fi�>�R�4.d�F��f�\����;(L^C4:��������9����}K��u����0��l��a2�'�d�Y��ZאF����y6��<.� �5I������� #`If�0��/�33����g���i��������/�����ǫ��n9��/��¶� �ej�����i&K[{9�o�1�O=p�17Y��9��N��TGh�o��E��k�m����q��ӓ\�d��G�A0/ևM��V��e�+a�3i�^C��Sb���&���v����3g����G�V�vZj�V]:u���y+�Z��T�'�������z5_�!�����K��@M�/�5�znӊS��iƸkn�-�C��B+��o�$���~�j*��lUf��M�Y�oxE��Fp���Lw�6?J���j��f�h#i��C*m}S��h�b�����~�$QF��x�F�Fۣ�Eo,ԦU��{ҭg�����BG2|������?X��GP���=\#�E>���8G�$d�@�UZɐ�M��?��{���sZ����m�R��t�k��΢
����n���T�W�n����ȼ��.~q��6 ������ZsO�#l����wB�l�nF8��ډ~����)�kF�]U�`l��FПB����5���I�.��z����$�éM�@��#�F	��4~^�S^Ap��&<>�e�-�H�i#�Oc۲B}�w��>%2�Ӧ�O�(C�6m?���!�}����f�}��^�#<�� l�C!*���A�O���2���OK_���Iz�<��/��^�erUxÔ�~���|��kec����"�]�-U���<M��N!6\$�/��ɅS��� �3��݊}Tb#�نV�
�ghu���E/��+j�2���Rw ����z�@E;]�1�}�[�t�����N$�q3����X1}�� s�PL5����P��A|�\OZe6kn�0k�Z�a1�Y�zl,��,w�O�BL$cS�����"�W�7]���f���9�O:�3	�TVI�T d!˭.���d�/Hp�F�mB���]���Y� $q�����A�6@��� �o���p�'����(�&c?�n��H�{�T��O�)�$�uza�O��%<&��dzg����͸�S�eʣ���tb�zň�h�F�4�o$M�S�Ւ�Xa>��^zc��?�j��_���'�RAS��A��D�-5�k��"Ms֊q2�7zۘ�M$#�ʇ$���-c��y�諪�PT�ś���_(�n̐����~+�M�����}��j�����tj:��!�/[��8��ݻ�X��`�]�7��J��P�c���P�~�]&Ft��[1�I�`�/n1X��Ԉ!����b'���i��WRD�!��O����~Io����Y�<ě��d3n���V-^�|'�o��i��-���'�&m68��O�l:S����uf��υ��|�M�����N�b��}��>gTUq&g�舙h��r��Ǡ�?k��UrL6V�Ԙј�*���W�j�>��)Gq��"9"�~q���\+v�10f�|ZJ�
#�A׻�����$c��M�Q���^����]�2�{-�=���!����*"w�3�~lM��4ڃ��&@�q�h��W�jt��F���d$�	B�]�8�g�8��?�H\P9��4���{/���Z�������4��bhۧ���	:�6��>Vxt�S����[�>�]���6q��_6$��p���n�q�ET?��������䴷��@I�U[���뿆�0Uɣ�:wFH��O[6Wj+�<�]��)��~q�}4>�Ko�ح�Lަ��Z�l��)a0yD�n1U���2�c��r�����͗[�z>g�VCV���4U���Ȓ{9��,�?u4t��n˦[�ꇘ�{¤�ʽ7ut�i뾮/�����Z�1fn;y���^��O��Rk��`��@rv(:+ʣ���"�x��X�v���(�z}��"��w�޹@X��=��7,o`,�˳��ki,�>�B�[ǒr����T|�\ ��`:J�m��Y��!)��iq��[Be��W���[?%�,6�w�%N��*��$���ª��4��n�����j�=x�R�{���|Z��\�-/ɖ�Ct�g����2��`o�K��K�t�!j����;!�:�O���E70����3^��O�VQ%'ХgS�V3!Bx�{;��Eei�u0�����"�����/G�k��}`=�Y�X���r`������14~�}Q����'~����ʟ�5��S������0�[.��T�?��Z��RjXC��_Q4s2��&o1�Y�x(�I��_�S�k�˯:i�ج�w0nF�jٟ"�SL�妃�^�q�:�����O!D���w9c��r�,p5e׈|Za���ւ�/s���K��R�7��d�� �����p���dİ,B�`���'\���l�1��iA��tu��_���VVj���m�n��P$�k��Ft�)k� Y�pˏr6�l}�YϏ�v{��\����8e����a5Jh��1#�E�~�� �bv���K���Z�9,�O ��n����>�,�����*�AJҴ���C��G�1]b��������#����ˡ0
츜>}���
(T��6�O�z���5ո?�?�Щy+����W�ca�ȫG���/=�ev��%��=πg�[����^��8n�wy%�$�n}_�v����O��c�s���b^RUo"LA�;�%��N���|9Ë����ż�i�T�������I�*�dOnr�y��7K��OS��8*��4���.p�e�&����Z��m<a ��NӜ��1������*`(nY����Q����&�F�Ē�JS�x��#}��k>zt�h�3���&�9��o��������#�u��#�C v�֡����?2��G�M��g�15}P������`"P�g�SA�>��� 7��k
�J�Y�@a�C�O*{<z�}��<j�!�g�jK�y��>ϟ�#_��}�;�t�2H�59y��h/���6�՞�X*?���R$��_���e���b��-������3D�!����R�ӓi�������L��*5��Yָ������Q/|Q�w_�X�2�"s��!N�'��H���!�Z:�l���`�����C�O�A�>��l��Ԕj��m{vY�4�0���,��F�)�e��?�i�gݿa�1����#��J0Hv(�8�#>�B#W�b��<��������:��=��;M��"w��^��8�ǳ�������ְ��V���'�Xd��z%zB^��/���-�.�z�s�6ױ��/ }��«�T0ǰ�^�#�4׊����4�3���o,���
9���¤G�<�O~�Rv[e�P�	����h��!������fwW)I:v���'��n�E�Y,X�$��2u�0������(�X��$��%���!�fU��	3�7SJ3��ϯo���
�zy�đ�1�v��*���n��v������>���Ʈk�)�kn��oj���ni�Yi>��4�I�Zd.F^Z��%��?�H�������6�[ѭ�Ե����G2h=9�
������}�5���-`��E�n���FqL��eg�*S��� S�'@D^�<F�e	�ݛ�]n�)wwn�۩,d揻�WY�Я#�͞]��=#�<�@���B���KC�G1��@>q�;o����grk��}]b���x���$\�������Y��)�Ӕ�g��؜���d�t�[����}c��\�������$)�ĺ����Z�rp�ՖB�aB NmG�p����y�M).odd�[�� �E���jxT��*4�F 4z�2]F����X�j��<���g$�w���oz�i�����D�`����HsL>��;�)���?z��t���I�_�V�~F���8�j�+=�DM7���C\KrY�n�Օ�8�dL�_Aղ"I����͍Y�lGo����f*�,��ݴ�^�����Ѫ���5��2��h7���g�.:Ҕc��A�bRr��(JΟ(�X�eC2Y�.g|�co�����^�aF�>U��6�/)�� K�FB��y��ׯ�ѯ�L�7���q;�j��q��ӎ.�1#����/�1�O*f�Jd�b������?�޲�`��.��S�@�
��(�������]K) �����PR���=�����`>̳��{�����*ߴ��]b�n��?�}lޟg�ɢ��w�Rz�b�L8`���5��:
ݔT�dz<F���i�Bɓ�}4�ădП|=lM3"�A�J[yJ�N��m ���;�S�WgA���c'Nc��.�^ 	�ZA�c��x0�ͅ��9�����f�`@� ��C��X$>����@�b�w���.��<��C[[_a�q�}&��+_}5�Ȉ� ��5�����fRV��c��-���)��͉���u�@����v����j+�3���(_k�N�H�j��E'w��8>�'95��*��^�K��	;��ž[�v��) `�s��]�Vr�T��R�@t�c��@o�!����d�oԣ�E��R��I���m���?��������4�5�O`�K�i$�g�	@���`�Cu���d�P-B���O�hV:�='xj���ewٕ��v��۶N�ֳ̎0��'^�s� ΃]��^�����T�x�#%�����z�Ԅ�t������(�ݏ�@^�����r��R���݅b"�:k}<M����S�X�u|8?8_�M��S�cR�")S����#daa��
��S3�󷳎z���!H_���zy��杔�{�b�a�@v�n|�X7Z�	Ӈ��7'r1�N��b:��9�}�E��XW'��Z`�75;f�����R�����q�T#�PF"�E�)��V��~�&�O�h�v��e����=�O�}��JV�q�nGDa$���M�68��$4ƹ�UM�2H+��_���X���1Y+��WKzY�j�-{[�X�Ud��a�{OZnwzϠ�H�ҽ>��#i��3���D�yqW$���M1(Q�l�	�&�M���zxN,?!Y�S=���Q�:5f��-;�4�{��*��Z.)/�u�^zp��dF���92�d)1�NL%�4�����;�x��Y(2@�'��G:�':}���%7���ھ�K��?Ǫ�:�Q,��7�E� �!_?����	�d�m���#��Gq�ZԔ�Wm%HE��?N��&Z��ks�H)�(y����U{�'O�kz��E^z�,!���L����g+6��D�����/�4>Y�̀~dЍλ�4��A[����8(�^���Ϊ�yu�ǰE�X.t�0^̻��IVI��&	=�=�xs�fƬ��xd�y�!ɩ�~�S��&�b�L�ׯd=���ۙ�߇�2%�?��y����g�|~��3��Lf�Eh+�nX�B�8�siOw:��m�S4�9>���Rl�Xhv�	>!�{�ʖi֤����!>���*�\���K9t���$�H�p����Ǘ�ᣛuG0˅�߂�[���-�z%��g]�CA�y����-ތ(�9E�\��sg������ޙ���"<Ј�D�Y�n3��.`�{��b������{y�ޞ�پ����w�u��:�'�Y�x)���y������,��ި<�=l:	݄�o����F��C��a �Fg�Z�Z@������I������~\,��p3����7G��&~q굒rZ��e�p��������Wf��K�b&���Wi�c��e[�����| R�d�E��r�p�Di�,�3�.ڊ��f&��"��<�Oh\4q�+�oHr�R��8�:��M�&����t$ ����C��{eT�n�x�;|�x�O9��9ޡ1Ѷ5��Lr�e���>2�^�AD^��t&�cN"_	�a��3���_б,L�t��e� 	.o/|�?JN�����1̈́>o&,���+{���G�h�{2����0�v6��<j˾��2f��R��ɭ�+~�|sߓ���8�#���D����S��*̜�zz�7������J���\�pK��/ �����6�Nb�`Ƞ�}y�w?��0�m6�5ɽ"ytV��J�Ҙq:�D���Ɖ�B���8�=��S�nT��&�# ���E*��o�M,9lVwj��o2]--ֈ�1�±�6�/w"yYη�v�`�VeV�g&V�y��֐�X�'�Э� >5����w�������ϋ2?�y��\����:��E-������E�g4�����Wߌ��ޙL{�ә�[�S���m+ә�Z|��u�Sj�/�ȀA%K�ߛd��XѲ���1O[�����g�>��:��9L)�_2�NlU&,�Yt�#۱���}x[
K�A���bDկ�G�A����S؇/�6ͽ>���h*5�psU��tï�f��:�A3�M�x��j�����:��_��&�w0F�/|^�:�U��
;k���+)���%.�	�+>���L�L0�~_q�ݵ�g�6Pڅ)�x�0o!i��/0�C�2Q�>�e��v�v�G�����q�߈]n�һ��n�f/�ַ(�b��&�SW.�ފ�eբ��+�`gGX�g�ЫQ�[��4@���^�?��O�ox{t�O�}���n��>���Z%@�f�F�ݾ�/�嗸�Ӿ��m�M��7���xʳ�L�C@l�����͌x3��	m��3�3��X@�*�_�pi"K�k)JM�O��@�LM��� L�A��4�(ҵx]�U_�[�؟#����̐�HP��yE�Aΰ���t$g@E�vI�m� �~������	|q1���o�f��<)̰BKn�H�Vou��c�>`j(P�7�<������p�b�883��u�ZX��B���8�!/[I�!�oo���X�KC�˞���!Dd���H�O�� ZJ�3~�[�t�G�.�7B�X*���e�]�������a��\BwC^͡v�S�O�]�shN�7V)A��R��#���D�m4o�Ȫ8���Cy�V�R�7�M�"��"^�������w���F�@t.�73>�Z���4#�{�zF����嵓D1��]���<m2Pvs�<�M4��86s�M��&�#��u��4�c���]�TO��E�$�?�K��أY ���7���J�����p��Q�L*�9��5�����k �d���q��)�P�ێ:a��ɟ�MR*���b�������D�?�O�zW�QN��c3lJ��O����4ǰN�^�uq7�1|	΁�Q�^i����F�P�������Œ�=NB��x�a��T���7PIU�Y2�8C�� c�ȹ�R�`��~�/��x'�s�.��$�4mh@��X��u������ե��R��\}9AQ�܀Lk���`������ݻ8����@`�畛�{��an�8��$d��A�������*/@:������6_�JgtC�K6�yHiE7���9ad���B�M��"��W.�����1;5姮¾�\��\;��I��/�}zf5��K�8;Zu����V����}��M���u��	�x�������$�%����@co;�:}���ᵙvO�� Ͱ�wI���ؾs�"�	4�����c.����>�]��FG+�?]���Uw���쟙(�8^S�Ug�yu�>p��:d@�2�ą3�]m��A X �ѻ_ݤ֩��S�=�>,h\��ʜ�0�	��+���+D<�m�/�/��!��%~X�M�|���_�ݹwil�(�]�j�	�Ǽ����0
��W���d��`��n����	TnN<rO��� ��G}�&��%�%��R't��2�hp���(���|��2�0�C�ii�� a��{���d�Ʊ�[ۢa{D|�4�2g䀜\}� w7:,�acW��\)Y!3eqq�KcX�~�V��8�s����,�Aa��|�:��a��(?��ˇ�m���FR*K��M���l�3��a�8�l�E�t�Q��Ƈ���A��ρd��e�)�?�v�y(�|����nFk�Bܸ�íա��f(.�ޥ�I�1���Ь0d�RM����$m,&�,����k|���`?��P��e�u�z9��T*��4��$�W��w��̫t������7���k����i쉯D�7fhK����:)��uu��G3��S�F�C���vI�
 �C�be�W�c�������L�$�*�;���r���t��U��f�#g�"2L����͐E����a�����אZOo�i���,����,���m���?�O
�a�X��k���n/}�L���D�7���3�]�/��־�Ճ�'�+GS�'=�6"pw1��$���S�����@�����w<s�>�C��|�'/p�@��Z]�O�<~�����	�?���k���o4m[L)�| 5Z�����f���,��;%�3���-o).��o.i�Pw�H����h��mJc��⽬b�I\�������}@��^��Ӱt�֛�3N�k�;�=�>�������]\�.�P�M�p�A����A`O�|A-�?�������!��Q���^N8R�fR\�aq�A/��+����?�o�_�/l\f�<�mm��/��[:�7�]�ii�ώ�@Z �1�fVu�� 0H�{T�_~5�g�V�xꋾ���kA4�.����'��Į˲O�0G���������F'�ܦ誣$֕�v�gޟ��F��w�f���#�9�q����(�zS��7�Eݩh�=ֽ��&va�_l�=���a����Y����W��bU�M�o��_r�Y�M��=����s��yC�S�Hp1<�kR���ovę=!�FF; ��;	����R���E��� ~U�^�,��i��6K������z�AsD�ޘ^���=zF����$��]�\n�k�f����p����6;���:L�ԱPo]�yƹ�#&E��G�#w��))���o_�Nm��@�S(9Դ����������T����eH�7�= �
��Tk�(�8�q�!�oP>RS1�Rb:���W�h-��O���Y�?�6H]���H�Ҹ�k^@F�<95	��z(�jB�ώ_U;O���1oPJ}�(�S��T����\Kt�D�:�MMM����,��a�X�L�S_��D���Fͦ	L{��s��K>O~ew����E��q����(|��:);i�8&QYNs"q����V�E$)J"�'�"=�K��)��Bu�q۱�"q=��q��夓�y�P%=3����I���K��>��q��.şY~���A,q��2���-�H��LiN�]���
6�]#�
Y%�U�{DF�r�?����,�]��v���@��77��Mx(J�W��J1~��m��^��{��Z�P��ޮ���>*K��k��JB/�z��+��0L�6��Vй�%��,�x2�۝6�����h�y��¹{�����2:6��Z�$<�`��wS��׎)NDn !Zf�/������Jߜ0%����lă�D}���9��y����=́u�99T��2��p��9��6�z��J��3�!Z5�cK��!@i���5�[v�k��2�b��a����:KQ�#���|]۠��y�c�-	�pȽ��?ĉ�$�	��BS�ʀ/��+��u�|oH:jC�\�w|,���E�<r���I�O�Dޖ�l]���՘�$pİ�_iq9��6���p��?9	eu�<΍͸nZ�@�6�;&q=7ؚ��B����A�^H�"�3ƴ�������������gge ��IX����A�x�T�	��:���5"����]ʨ;6����>#[+i֕I<~�[�����%O����h5�H EM�MD��kL-|s?{x�*FSp��U�A�wͣz�tM��fٙ���7�Ư��pSf��Zꁽ��5��%��a�`;l;�$�Z%��p!n ��������UdY7�������
7lEJ&t�D^�DI�9>p=��Q��Cc�g�M�,��<jR� T.g80zl͓��Jk���d;S�g5�)��/U�ݽ������oh؀��
+�ͺ���R�;"�%m^�`����.Lg���1�*�V;��\��8������d�a~��?��ob��^4��h���w�Y�@.x�1�ͭ���&�O+l\t�,�1���1"���)՚:e�ɭ���d�p�(R�=�&?����)n3�1?��������R?�UZk꼮�<k�8%C��nx<�°�z�{�c��� X�mE5C�,�|����A��$Q�.>���4�bUiS��UX�)���+Aȭ�}�X��e��K3j[�Y6�s&"Z)=�^�Y7���3F��O����n�x�)���='�Y4q�M���b���������yܴ3�)�x�Yy�r�/��Ŷ�P^�I�鼖X��J_���+���m_��Y;/�|z�x�(�FlWZr2��|}�ӿ�S��s�Л�����z�.8�:�/+=.��I�'����pkS�z�OvE�x�K���|�s�� y��璾�b!�?�MpLqbB�@�wq�w�/O]��Tؗ���y�YZv�t�O���@ �	���!�]3��雷����|�Y��0�8�U�RfHT���{=Z{r�qy�3�m9g�+��E5n�>����X}��N����<�{U�^e��<����ͥ����@�1���d$:z�� ��L�<�}� �?{��2�����H��1�m(��p�jw��>�᥹�VĆ�C� 'd,�K�\��Ǌ%)�M7�MpZӛF�+�"�EV9ȹ?@{���'|Ƃ~��{��BD'�t�g��[XT,u��m_2��^Loy�jvPp��u�9{��&���v�������VĵJ{RF��0�/�A�����v�a���W��"���V�qy�]~t ��%R�.��a����17��*M����q�4T���U����c}����q����G�MNB��w\wr�B���#�-N���%	ʑ?���XW.�!�Ro���EH��-�Ǧ/p�-�i��D˂���Go6�jw܌�,I��G/T�I>�'I�!�H�D3�J���`��������P,���2� �޷��ぴد+���;���{7-�S^�4	�9f'��^+h�����Jy�(�'�GK����g���ß�0��/D��st��ٻ~Z13������������~s�Y|:�=L7fъ���_��ϴ8u��3�h���t��Ĵ,wDx�>��.Y���k��E6{�Я�=�t.ޫ{��bv�]��m+ᖝ�_a��Acf��gn�nѶ���>W0`h��ض�k�fſӄ|M3 �0T��ඇ��KSm? ��25��O@YOy5��i�(�����Y���e��mݮ[.�z��<������F������?e �FD�	�wDb�<<�(�̲�Rn,��s�9�]K����8燎;>�<�ҿ0՟va�R����k����[���`����.�+ � ���ف9�
)c^�`� �~����D��x�Fiă�0��!\T�=P��}�e�#�gBo�*'h�9�AEKD�43�a����8��Y�zËho�h�O�<C���S��B7��G������ݢ��V�~;��k5��urT�;��I� H��I�#�Ǽ�tK^;�L�H�&�J�G��6癀"�EMJ% !B�=g��}�������)ߝ�ؔ@��cn�Ś�q]ݪ�!�_�;[��̫����~��!h@�P���7��+�G��ܵ�T��~��ѹ\�/��&;�u��܌�U��c�WG��K�#��S��q?��ebX0�x���o +t���s4��K峍 ��o�c�(")��a�v�dN���/,;k�J]ƕ_O�(�R���W��&��x8�K)�R���R�������T�W��xbX��3� �v������?�UJ��`P��RQK�I�(�K���S���+*%{l����tΞ�t�'�ܝW���p$#�ձ$&�$��Eó�"��9N������bb������D�1280P��0iY�C̌�?5A}z��9,�t�*�qG���X�]9���zC�t�L����h	+~Z�)��
�\P��Ӄe)������0f!λ�k�H����E �]�+��!� �>w���A��vg�'�	|te>�������u�|�� J�)�9R���Q&��
�J�05�V�vR�����I_�^����h�+�0��*�6$��"����<eX���П���4���L�Il0:ܳ\Q�?&�ί��^r����
cx�˺�o����]?�g��B�E}k���r�A��H��W
�����_T ��;3����.(oVcZJ��6��S�������CԺ��0Og?��:����[v?���u�C���bfvI��d�;� qr�Jݖ�g:`2�n8���K~T���Y���������PcXW�!�.F`+'+#O2�Mq�*s)͸����:�
l��o���vv���uĈ�us+����U葋�joyK�91-�����f����H\E�����i����/�#�����
V��#���ݪ腡�槄����F���E�r=�U�C"X\�B,5T���4�1�t2�94m�b/^�"f�B���$��!|�gԪE-T:�M�^f&/X�&V
��6
l^|)������[u�u(�Ad�vdb||�Β��i��)�v|�O�ph�8���3�:v�t5����*��))��%�>T^�LLolݙm\W؀f�cuI����P���ةj�E���x���X�a_iZH�~ӑ���8��G��?�nj�6? �o�����E��V\�� ��
�Oѵ\���R�ҳ	c\E�R�H�vF�����H�{�.��O��RCb���J�`(�xb���C�Kv���,�

[K*Y��uh�r,�k'����L���j�����5a�iV�1D3�
~c���@а0�����=�8���!��AO�$���i��e`�JC3o����� M���`gϦ�Wڞ����������>%hZ�2�.�|[��^��zV�R}��7��Y���l� #qM�N���=Y�4�r�.���ێS���,yx��S~{�kݣ@z&�܏>������an��p�	�[J�i�A�����:?�=���̉+�3��=���E7��Ê���4T�3�&�zc¯g58T�i/;�Lz
R���E�fX���$Ƹ8Fd���?�|���wL8����f��0/#�M�j>{}����|��E�P�OJ=�� F��G�u���}	*�X�uQ��sA���m}�|~q�xUB}J���:�������b#.�3�ҳ�ʻ������j���+��Oq�s���)!�׉AdA��=
�sі�Np��'qO�ϙ5�������5�+J�)ȓ��G���EY~�_�=�]"�"/��Cb^��ǵ�J�eC峵�<e]��+:�����On�.^jY����W��F���7�i�|�_��̃�89W/?kw�8O��)�Ey3y��b)���߭9�+3\x�?�؎��3ԛ˺��Vy"��Gy�'݆�%R���<����X���9,������&{@���Wt .�i�#������?O�a�+W��"�>�{���mi�l�fd}:�<C�E��<Bw$��c+\����o�u��,fj����HCǨ�[�&`��OƗ��A�Ḻ�pŚ�J�S�!�i�8v�*���U�KB-�Di�[��/����Qѷ��=�h�uUvn�an5)e�ڴ׈��dFۜ���� j�0��]oHMC��ؗ��j��d����E��/��<�ql��[��G(i�,�٩�\n�39T�A���������T��tf�v��:�X_��̈́�5��A��m�"�zz�x�=M��&����$VT7��?|�O�]�~U�3���F���%��?C�n����,��`��&y_u���kJrބU��%e�ln	Aj=R�w������l�(��|qT�
�5Fd)㤱�rv�~'+�^>[�����w���?[�b�EwNi�L�[�p�Y�}��x�'�t�hC�z?�x�Ő��[z�T6*���� FpM�����/P��Y�ͫ/67*R����(w�$���#�Z�J�B�������b�Cl�6���9��u�a��pD#�>�
��7r4�n���r�Jd2p�Bp����eGb�G��O&�8��^��&;tP�
��I|6Eaވ}�X�����&��8���baʍ�`&�ވf����4�
�Bu�#��ԝU÷���fś}we]�9������H�,�d'��P��ɱ�Odp������֟O$<�;�8�w@��MG�`����V����x�~(k���E��+l�k������^�"{�x��8D�/aذ�v3o%��ylO�o�|H��|	�c�@�L=T�ML�Dq�|~7a��hf�g|?���N�1����5wQ#0O.�UC.KV��r
w`�M+�{ۇ�6��S"�e�%?��Ќ���I�yB��|��`�,��rK����a��R��g6B�Cf���"���	6��Onc����8urbem��!��:���uO�{ �k��w=}Q'Xc�7f��֊��^�h�F@��O�ͮLb�!X�u�]O�dX�q(����Y
�����Fq���H�bi<e��~ڲ�csG�v�b?���^�N.�1���EnqQ�6ͯ�3u)B���ɍ�� ����d -]{o�^�lEm�t��K�PX�˯�_�u��<�ӓ�w��u�<���X��[��D����	@��ܣ�a;�\��q��e%�!����M8:��(��LӼߊ�-@dsF.:��M�n�;���p	�.0-C�qZ�����4��LC�I�	��	���i1�R�?��/u��2"�.�k�X���gBh�U���˯+
���C�W���"�Ҽ�(b#&!jV�b{L'��hK���r~Wy:�-.��Ƹ�����F��*G�Ovm��K{"�(��Ni��p��h3%�	�.��!�<-�� ��^�Ӟ��X� F�,��CH6���x�~y�0�וM/M�Q:F3,�2�8�Ӿ3�Ӌ�����$�4D�X�0z�����wNsL�Z5�w>f2 |H��'bТodA�p�N3�4՜ߖ��j�6���_F�dY�����x�>qZ:ҟȿ)>O�HU����^ј�.܅�U�L�!B��S�v�K�=c�͂�E�8��%��:%YԐ��&�!V�"O���o���X��z�G\&;k������-���b����xы��}�����7k���<Z���X�c�������;�E����_�,�����(!�e���K���K?���7rPQ�ŵ�	����;x&�����ɇ��ܦ^�dm����h�W�������j�TR���4��W"�q�V��o�d�>	x-CV�gB/��$��yCE�9`�e��z!�$i���:�!�R{<%�^�h��X���Q�?ͳ~ڕn��3K��n�w����=9#֜O�d�W�D����%�� ��Й��|���Sܢ�+�A����l�`��aX�hB�8�$Z_�-tv��1覔�W9��d�=���tHT"�nP�=�M^4����+�@ ٌH3������z��)ǬgA �ͥ!n�[:��zS�X#4՞P�Sg��!v55�����^��d@�A-_���)�GG*�<����,3��|� ������>�GC��_�Ҵ'"kX�r�dP�ž��jDI�}�pzI4�5f�A���A�Z��1����01��j	R�@h$1��z�qm�E���Mɬ�M����� J{e��Ғ�-�(a4�F��Y�^ L���<tC�Է���?fȧDI� _�k9�`n��$��������z�&�YGM��!qS EDZa�y"���\��[��aB�?�j��- �ȁ���,��������Ӥ�hϺ��Mm\�q%}���t��z��+�M��<��\;u�s�j��+.��5�4";pv��D�i̅���oAm 	-�=��@}���O�bS~�7�1?/���mK!�2`C)�X����$�vo��A�7'T�!h�bH��b�E���e��^�݇�C��]�d^_R�=�+����a�-�����:�'�~�t��Sϓe�Y�TKQ�˟뙍�z��?���S���HK^�@'��Q�T�{�\;�X�@����{�%�9��r<Z�}��Lap)rs�}u������m7��l��5�q~�t�C�8<�v=�m�R��6cJ#S�����RC \����	OFf�T��5��s�}6>��fVGV�;��\�#)Qsi��׎�������H�9���r��Q�V8"U��G�`�X��'���\�d/.+.�DUR;E4�X������[Q�	��'�Pr�UD$�e�d$�,�{TX��i �غ��R���3�3�3;�LjѪ�q1��4�gd�=�G�{ҟ���8<03�ʾ��f�ĆI]Z�d~����-�F�as����eMc�t��l\Ջ�6��uD�bT��f&��
�C<�����8��-���Й����E�|K�2y�!>�\b���雇9_s�o��@hm� :���
i&�w���L2e$�#BqK�,�=Sз��D�V��:�$��Հu0yY�G�â�%L5�疈��ߤ�;ffR|/��\>��A�ciԔOg�r^�;�@�P0���9k�XJ�	=�;B��:X+��n�r��K<~�<[�B������48aX_���jm�n��0��9�޲�xJ'*7�)W#�!�1��G��e���q�|���q��-�%<��o�c�'*�QM��<�h1wY,�y��!jvǊCo�4�V��%��{���g��[�������߉����.�fA%�Q�o�9��/�Ō�����g8��t��\O%�}
�4 �	�dV����8��;�mʠh�ֹ��Ë��Hj��j�K�`�8=K�kLЖ\<x�K�B��:Fox��׾t}����Wu��՗��/]����}ż���� ���
MN�ák�<ꁳ�4�ޛ��'=����eΙ� i�r��>���g�����ٗ�G<���3}��υ�A����$}^񝜼�%v��2iO�|��^%@�R��6�M�K��AFߤ�7�T�<��?u�<����1����SOd<�zmbv���;�t�4��j��X���s���_�a�v��i���П��rٺw=fT]#�����ҷ1@)��g�5�$	$D)+F Q�G `���E�Z�J9��]is��HA�8��|�K� w!��\���	RX* ��ؼ�m]ע����ָ��#��ԙ*�~������T�G�b~�e2��uM̑V\j*	���}��o������11[]����-u�y��[�g<��!߇>�zB���</,�x� 1#NË�X9�"B�A�[�}�f��8!�J���R�.U:�
°4I���;�FQ��R�!���js�{���pZ�",n��>.��ǟ/Ts@%�������h���Mp��*_��_V�z;����w�4��p���M]�^���[Rf���w_�6��mi2����H;e��d0�k=�y#�D=c���@ V����KhE����V
�/�a!�j�b�;�ƅ�iBX�P�4���������#5��3�Ok����s� n�!G�&/�G��O�'l<��&�cE+�rEԥ����x�\�'��$y􉈆�2�CT�]�hN��9�̲��i"��ge�W��}U�y���F���G�E�:���d�5�E�Ѱ�U��q��O�(N����hf�ֺ��83U�5C�~�E�_�W����ʷ���-y0G^xk��k'xk8��AC�i��wG�N�]�.�T��qo�̸�#$g��H	>W3lx��:��[f��rP/cft�(&
�h�d��������:�t?lZ��w�Q�fH�*L�J���j��<�7�@S���]A��j����I�>s�X����U�b����է���"R���p~"��A+�Ǵ����!�7B�~☱��4h�=���H��C;��w�?.ܜ�,���>�l���-
��\rX����VFd���V
3�A���v�g=���yW��׍U�*%�D޼UJ-�@|�ю;:�y��Ѧ�����%	S���ukt���2*g��~/��G�Hs)��%����������nM���S6��uY�?.�_���w%��f���9��
�����~��#aN�f!e�`�e����j�Q�|P���zy\�7l��A��h��+Z
/��i�D��?q�?jB3�-_3Ģ��O00�ahyԗ5�p�j���<������pܪ���v�[kwA����o�ֈ��X=�����q���" �e�	�J����*C�r��%v}�� 65��7���L;�ۯ%>���\0U���������.�ե�`o���cT�?����&��/)R�./�&�em-$�WD����LФ�Мp��:}��,�E������K�P�G��)#��GwK�"����$�p73'+Z-�2�#��^EOw�*p�n�d4͆b�"e�uZ����5��k���L�X�s��s�L������a,'G< ݅ �S��`��kZ�y�S�[�2%u)F�gd���!8�������v��ơ��|����J>5���ҘO���$B`g�" ������I��}XB��k?�y}��4j1�G��Y�(]1l�Y�ru�u��c	���;�x랎��>_����J�D�U#J���{l�z�D�d��޶�v�r���\Ӯ�1O��_��Υ�
l��=�X ,M�[�N�z�X_�)�q�B��A�i������g+�b���Z��M���B{=�����S��zT�6��4͇�|ˍtJ��wi@e�[�(��Vx�ȸ�1��F�꣺K�3EFS�����<�va�&�煶�̞�5o�9v�7u�����z�1+f?�};����R��2�3i��Ż	Yx�V�gkb)�W�b������:��oi�2�E�l�@�]�b?�I-�2>=�U7|�O��EV�0����EO=��'{�]�U�6�ܪ>����{��_R�/;��OY�_އN�90t�M)�d�2Ͻ�aS��Bm�[��^N^�������W���?����d�@B9k�#陬��nڠ��)I6>^��.0��n������ډ���&U�+��xq��A�U�m�vmw+J"S�*w >���pQϗ0C@h�tv���6�o8>��;���	� �1
�r�_�ˌ6�M�	&��Q�	����L������!.;(B�Ya0����W�u1>���U��~ ���q����x~R��5�XS"��P�kt#���T=�⍵bJCw�GQ���L��E{���rL��cI�mn�i�]п��j�p��Y;h��a����{?-im����(b�;Y�K&4��@��|Y;�[�}
��섨�G�����f�&��@
j+z,���%�k���BK�o$������Rw̭"��qE�A$��I��A��``BN�*�)��O?4$�}�;ڎ��D�b�Bq�T�3<j�y�"�4�L�*�)�{%p�;U }(5�z���V\G�s�R�:o*�`��oOg��Z?��CZ���n�W؃7Ch9���?������F�C>�r0�drcP�l��i��2��J�`�7�_7I��6s��|u�5%9Д[fև-*D�������댳c��d)�R��I�],�����2��6�1wO<7#����<�����o�c��!.�m��E.+}j��%���o#��]�O���6�}��~ň�1�Uz������e���c
XSFg��V��Tk!Hb�?���N�π�̳1��W�O�
Z|���uV��*T�];�C�QD~T�^����i�C��RՋ,$�(*Mz�O¡�����~��h�#ٻ0���o?��bګv���uS��O�3>��hA�D�]�;)��0^�?��$�<�kNa���3|\RX����$���¨O��f���?�W͵5�B�3�G�~~���~}"O[��^ �UWB�Te(c��~�{�x���^�������������y�~?������<�&���e����`A�`>����R�����Cn�j��$l��ki���}S�ʪ�23,�-�:I��<�!�����bPSȚ'C�7.F}w~��} LU�T��gFW[S����hY��z��W��n�5�Oc�(}Bo�S��k�K9��e�c�}��
eg��
�9T'i�.?��$�#y?�1�1 ������GC�D��8O<1��f�fӎ���h@} eLp�e�p�o�c܃���1Y�?m%T���>�NH����ҕ���N��P�\��&�[i�XK��[c٩a���U�x��t�h]�(�;��o��=��x�ˀ(��y �;ɥD	���DJ�{��n�.E�k)��X����~?�{���yy�̜g�Ƭ��iQϏJ�z,9r#.>����~�vg����s��`)5��	l�&�h�r1�4�H�ς�l���4��fc�e�[��a@�y�?��!��)��e����F���*;�r�ZǍ�ז$�	M�m\����x�g�Q\X�z�M�o�ޛ`��������%S5x��kW\2��\i4`!�@9K7�%��4ರ������{ʹ��擶?�o�f��A�A����s�L��v���3���i�C��[�V��<����,�>�ɓ���
��ٟ�l��S�+��L�.kL�J�����0_��Ry:������F�'�V��f�,=��X�)�z�C�VI������ik��:kPZgGn�e�Xo�+[�\3�ܠ���G/��'�;i2�B��|U"�,���[u�ױ��t_j*��� ��.�l:	������G߂L�x}Հ�	>oB�����M��BF3.+�����m��ڵ�����9F?���>�����P-�������z/�)����{+�u\�c(K�ЎǼ�|Sx��)��\h�Ṛo�}�����b��q�!������R���iO�*�D�|ϳ�}���r���&��Z��S�����D^�v��D�\<���)<"w���x��q<��
��r�Q�M���#�[!b[�g��O��E����n�dn�Z�g3k��ҺRK���?�(,����_��c�o�**i�-[�B@R<2Rը����י��6U/,[�8���Q�`��Z0�3��]ܴ��;�����o�wG����)n�ˎ;O�j�O�y3��'��O{�F�|,2)�[RJ3��G�f��a�Zў:�h�4
0.�����`�?�2;�Lu��N��b`���-J�w�J�))��l�uʀ�U�Om����D^��Z�l��2z�{��Ī>�l�������0�`:�*쇻����f-�X��N��{�hr:���F�n�L��XQ����%�gsT�;�-�І��?��̑6�L)�U���(*��gzb� %�|��0���zF80s �\�qD����8�yG��{f�!��' ��jn�VՀ��l`�.�xWOЗ&��Ι�ƢwL���^D��K"?9-9�(Zo�j���D��a�G�k���+�ڟ)�u�xBa}
Dj`c-�dE���T뇳T����~�z`P��À���q�&��s�'�\Q;�T�ߌuZO*r��'��y�n���k�!����&�Eoç�Jof����n��Z��;��&0���d;W�)��`F��x[����r�!Dyl�E�t�X���2��t���~��~�`���I��X�_o"�p��U��S���q�5�>�����^�9<�coJ5A!���|iJ-_^�N�r0�S�T+v|�f����<�m-��/V}�hH��ۥ�F\�mg9���v舠t��oX?�8���0b���׾�\��*m7Ou1�q|���D��cɭ�T���7{����(�E��2���ׯj��B�j�u�<x��9s�׼���]�z|4�k�����[ZeO�Ӛ0��1_�_������2܋/�|�`���<�I��4j6��0NT&,�Ο��sN�O��l��������v��f�� !���}j��@��O�e��3E�f��R���96��p=�c�x��κy�A�<5\�����-1p��E�柤.�ׅ|��%Ah�=�1رa��.]OA:�Ni���C-eQW�˫���k��s���3��eQV�(s�&O���}�ܔ{z���֕�P�C
4U�i�f�1����U9���'u�߃���nھ,�ݩ�q{؟4A�{�`��s盅�/t#n�9��&�_Y��&w JcBnI��` >��(L[��v�Ɇ�NH9�xl�:`?�J�&�^�W�T�u|\�"Y��S5>��<���Qh,_0�Σ�\k�G���_,�q#ƥ
�S���g��5�a�������{�,+��X���w
��d�M�S�������ԁ�AzX	���̏�ԣ�H�{9ʑ�4��x!�F{�-�[��,��O��b�a�Q�rVd\"�5;��@�6/���_wQ��T�^bJe����K�J<�M�*v���,�YT٪( �y|���S��&�p������#gM��0�h�A�yT�>p� ��ϰ%Gڸ4��ʸ�\z~�[�9i#VVj�����k��\�C3ع�R�4H�w�)g`��S?k�yVl>�˧��ں?�?~f!��ٓ�����؈l�~�Ȓ�AJ��d�_��o
v�O���SO�=�2�'�~��$�����`w[�Z��V��ɾ6����m%�|�[�qx<��H�̵�M�0�V �?�;tOSW�&���%rZ#�(׊�0 ��~s��K�����4l����p���sM� ���N�Voh��L�q]+����R�ȑ�^�V��-�$�[X�_*��psH1�����͏��������{�)o���Ǣ�	�e~����!G|#����t�!w�C>����������z=	ѷ� ,xeQ�>ڿw�]����j�&'���LH
�V^��7F��������j������NO;,�8M���6���;���l$ϱ��E�����6�p�ȥ��Es�/�m�V8�+U�%�爣�yA�/V���?e���_!���ˠ�PR�^�[�H�
�?2_i��`y���,1��v[�QĘ�˵�~���<Ou2(pԲ?�Kz,�v��mb����}�������N��f����6���tz�\���[����SJ\������P[�/<Y�\�eS]��W=a�:��r�$����8~l��(�נ����1Q�J0��䰐e�>��~��?��i	��˫Q�3Ȓ�}���
��m�x^���i���n�u�^S"��m��Y�R�	0t�CC��&W��2����{1y)�;p�8����k5{ڗ�jg+@w9��P��M���)����ā`>�������fM���$�jVz�^��ҷXL�q��m����B���6q��A�N���;��Њ��j�L敿�ҭ��ʓ�Ѯ�s:��$UR�����$K��1�ѯ�U��xOF�Q~��?�������]YB��Bb��2�(�jܩ�6R�L�v4��+�i����㡹f^�f#���K��4��gʟ�g�F��� fa���ΫyL�|��8��ϸ�8�_-��h֐龶�:k-��:���w��=}oj��RB���P��>���c��5[7�!�IS����,Q����� ~;��L������Gp�#��r�Uj�f���w*���^s޼0,S8�z 5�(9Ȃ��`,�o|L�cY����Xa� KʣM������=n�0�!��Aᑳ��F�5ח,,����2��Ϧ�Q*��R�L6F�f�;�y���E�v\�0z���B���g#�u�@M�,}B���1�7�(�L}1�|tT�#&��v�QƬ3�]0��p�|���ZԷ+�/����B��a�G7����eu�s�O��H9BjuC�׻�ya�3��.�0A�g7���H���0��3���Þ������(���R��<tk�4_BKy3ғ����W�X�=�/v?��v�0����㐵�r��s�}�os+�i���n����R�;�Q��J�i��p����>��M��*�xU���E�s_1Ź��vu����-h'���ȹ��wR���u�AH�t��n��-����1�,�:���GP���3򚏍��;űx������(�&�Iot;�1�OF��K��~tF�,���6���#P% (qa������3H8�]fU�7՟%4�t4�$��`t�1�XBT:�/eQ��N�p��}7�h��U����{]M�6���_�]R�$��U���w��ז��G]������Ƅ��/�G#�iMfA��zX���Ǜ��̢a�2��"�6��y#S�O�g���S_˳[���q.7�\.)0�+Gᝊ�yQu���.9q��öP$�J�� ��g�u��$�ۖ�?�AW�fU���[_�̃C�����57R��'���\uk��f�[LwV��rG&���W����00��衡���dK�!��U��<1툽��Ma�ݨ��c�H�W�I�`�)��X�b�
��K���Dů'��މ5�ɍ�;t����m|�5�����#ߕ#Rg|���S_��H���x��h"vU���ǭ4�O�rd��hv�V1�L�w���Ԭy�O��`+��B��p$�pd��bi�Q���'0+u���wy�MX� uLp<� �_�ᇀ������ ��CV	]mf�u��|�C�k�Kru��0q�*�Ǭ�y��!�9�G9`������b}+,��!�#�%6����4PC|��E����a�2#�[GJ�t~�]s����w�rJL�a�6�`��N�UOiP(��%���tX��E�ѶʟF�eS��۫E�J����[Y���\Y�:�mN�痸cUO7�\9��:_B��6%�;>3*�3�k��w��d��n2䰦�9�c64���)u�����,cN�28������*7��CE3�O��w+.�q���9��o��������������+7�W��B���|�ѶM�5~�5�=M�����4����4�CN��Q_l�'���,����ퟡrM_��5���F29�6Q�5/�a=4Sh���8���-!z'!�-���o��!4�6'�W���FͿ���e�k���-��4�[ioX�Q,uq�Ŧ�>N�ֻ͛dԖ�9l@|�\���ѩA�M�I��&!�w�q"ɗ����(����B��A�����,L����8�j���W9��͎;S�B����Ɲh/|�����S�$��f�zƌ�O;�ϨW��V�%V�i<?Tt�ݖF'̭�̙��2E�@~Y,� U�p߶%EG��1g��I!$��tꤲ=6̤�AD���_(�daMJ4"k�))k�D��7�A��]Dz�b<օD���?�9Ţj;</����Ї��Ͻ���֮!�����P��d�5�m�с�D��~�YgҪ3���7nbˆ
A�(���3�Nt�L�C%�P�ԩ�Ͱ����wK����j�)��+�b��B]�m�ߚ��R�[�l��[?�a?ۘ�u�~a�Ɏ�~��c�Z��˦��^|{�
d�<������	 �u��6,�p9���l.��!��2��1�k59J�.�q���b��|9)�B���F��yI�:m(�gjdMx�6n�q�������s�}?�����p]%j��'5n��r���B[�5l_R�U9��ۂ|��k�%ۖ�9�f&����ݎ�@a�r���� �by�
ԍyj�,�
�]��o�u�����C��0�Ѭw��X�'�B�I�5|��F�U5��{�6�I�D���eA�2/=$Z�;���7���}�N#�\J6�S�Ne�����Y�p��M��l�X�����!g�/X������J�1�譅�X�X����܄���G�D`a,ڵ��T��9����#�at��.��4�l@]��Y��}�?�������U�t{��z��|2�^�7����������l{��l�e����p#��e��s�����rF��.�Oj���i@%��FK�V%-ÿ���/I!Dt�LY�_����u�	$�f�Z�$�	�|YP�q�;�:pS��
&iUB�4I�g�g��
2��cC̕�O�.�s��w]��� [}PJ$�!_�w��*gSo��b���ٺ@{�� ��;���=lh�O�����4+P��'Hܤ��F�X�e�WA�co��'+��5+?d.*K��sYu/u\AV�~� u�������������Ȓ����/xNEN��( �����z�x�SaqVC�M}ָ_.�U�} �ܗ��%e���i���ԩ�~T�a3|L���K����򅵼l�9ķ�ke���.D��X��uɯ�9�1M���I�q~�Li0�\��j�D�|�56C,�d?�l�s��P��z;���~���k��'xK�2��`�s	c�M�e��ZH�Gq�s�b1c�sm&���GCޥf���W&@J�}�� 3N�õ����ƿMbtIM���l� t���aNȣ'Y�5�u������#�JL����	�s2�(гn]d�0�hSn�k�j�5��޷���,"����\3u���j�][C�9u�7��V�[�d� ���a�o�F�r��2�'a��s�a��ÔViic�+�z���(��V�^\��`'��7����i�����B�����Fs�/���ECm�IOtG��|��4��'�S�.�G5�8F�-��JF�� qdom�ٙ)w�F�&+i�Pt�_����lk���tJ���fG��;���ǅ�F���욳i0?�x�6Y�
I!�c1�M��!��6y(G/ae]���1p�w�A3����ۼe�QZx�qǃd��C���ݓǨ����w?����Â����]E���v����z�����=�n|�r�e��-]�m�H�����7��?w�w�y�zrAE.�r<���.���99�lW��Y� �ࡑ�QkzŁ��i��Ԅ���$F
�F�L&�R�qsl7+��G�	�YgWV������F0�'O/E:�3�]:��(ʩPRN�j�6��uu��x��'��2ٞ2��6�M*��;�iDh
ʚ>,d�^f�,�r{/ብ�hB�Ǳ�|g~�9��v:�#�ņ[n�r{�+��V�. �p��-_v������^5<݁S�pD��	r��(5<Գ-1�����!�R���?{���W島7y�>�)g�����=I�Bw吂�������ȴ���5���7ϥc��mYj���ng�!���� "ɰ�-�'�E�i�%j<5�T����=p�}ꮻ��B�
[�P�/(�&���"	WV^�.�Klx��W�I`0����y�%0��'�;0@@&�ա�Q�&�XYQ7�M��U[�i�4������s*����ʩ�Z�ɋ���Ͼn��=}��3���6i�Ȉ�C,i���Nڭ��i��=��g
ǟ��w���������jGO� ���#����:
�s���Kc�sx��p.�]�%����b��O� �O�Og"�>gu*�K�w�U�%e�CwWg�.���fg�6��λ�e9�d�)����J1�#]C7��Z��CخmQ�d�) ��ղ8Dxq��￟�j���j���1
�h@�t:��8�^/���h�W_����o�G��t�5��.y��[�I�ɝ�BMӑ�q��|��v�ĳ]�K�hֽL^�L�O��z�7A���&Y�,���o?�
Q�h�`V���u�q$~�I[9��H���S�ȗ֞��PE��9��}Εje6��C����{'y"R�>�,�,��eӧ�x��	��dn��������Wl(3N�2�UZ�˵�h����8cc���L�,��@�Dʐ�Xڧ���'���h�k��kS�����	Yf��ü��7�ӣO��tbv���?��O����2֘dg�i��γT�m鷽�{t\�g�>�y�#��6gm�}�C#�o�b�1(�c+y�����9l:���u�S�UO��}Eyן�nwg��..��FESG����p���6��ӈA@���焀-�����lf0��lO�S0�S���7~�"z|j���{����O�����ٽ>�'���E)J� "��L�@Q�]��Ȱp�=ð�9ɂ^-�P"^
O�Q<|.z���1Y8*c7��~<݈�v(���A��mi�*ïK�S�B�ɤ�j6f�$z2�1]�u�p(aL���ָ;t��_KH��_����C��B\"0/*��Wd��ܧ�Y=�-3D�I�wY���Jx�7L/��鎞�X���i?-,\��KE;�����������<\�s��g��_�'���#`	W���W�zͯ��j���d~�1�`��h0��y��G)ջ��>)�k����7 �:'vZ"��%�e�LZb��F���~A6��ʟ��}^Tq�k.�s�LQ�M������$�
���qu���j�`��H�߃N��1[����x�~/��)�j��?�7G��}�M|Z�yΫ���Jl�j���QJ�P����ˣ�$���U�ĺ����<�}��x�!��ޤ��=�c��tÂ'ߎ�'�"�>2L_�? Wb���Y�ڷ�2 0��W���8W��W���۸�Vbu��Ĺ򮷸�f��׍�CЯU^,��y�?����_"¡o<���[B�K��uV��&7��(l>[�\^��q{�f��V۾w��~]B�I>��C�i��M:{���^^�d���[�t:��u�c݉g�]�e��eC3{��-�Td�/y�.pK	�7�"���r���ޞ2�Y�Z�er�h[�t�ˊ�����oݳhzk����l9lK��� �g�®$i��F�� �;�0L�1�ӿ+_�fij�"��AI��<�`���!�N�������P�j?'j�(R��5JC��:k����5q�|����&��e��=K��d�}����ή7���x�fMXE����)��w��J;����t�.�)0&s
?E�_�(��y�9Jõ�L�e'b�h��h�B͏om�p/~:�V	�}�����0�Z ���MK�I\�a^��ŋ����le���:[�@	<�1S.3ڼ�����R�mT��y�9:���xr�}��<O*k/�ښMr��3����pbK����|����a{��R;'of���uc��6�5ͷ�g��t�G�`���#՝��PC�C6����A0U�4+X���M��N�{u�T޸M
jA��AD]�6T)��:j)�S�g���"@����N_!N@~NZv�u���RF�+�]��->����*�7��i�m}�X7�����n��	m�B�$+���5i��q'?�#�j	�%:%'��y΄ �Еձbibn,a��Y�ss����3h�����<a�~�')��{�[�d<YA�wFY���"�������^�3/iߩws�s�}�X���T|�E��۵�J���~�VΖ�A����r�Y�Z����S�-�n��H瞐��_�>}������Կ�1�
�.|�h%b	]h�C�>t��V'|�.i��1ޑd�[ًR����#&�m�2�[ia�� ~Lɥ|m\���`Q�S���&�c40� ���D^��ߡY�ߊ�^[/OƓL%�^?�(���	�8`�%�?��A	��m�n����Sk�&G��{���[�K�DfP���Zd�G������,����f"�Ժ�D���A���!qZ���/U#�l�8�\�$��be���>~�zo()�9{�o�{s}�	��?@��h�$1��:�T�"H[Q���
=_^Zyd<>��pom�����oF6�f�9
r>�$i !�D2��lK���ʝ�("`OoH���#P�~��զϪE0�:%3/1�@�TƇ��YDD1E�j�-+���lOz��:e�|>߿��}vDsn�Rl	w��SI����!���6��%R���wvZ���5�߭=RB�u��4�;��8K����j�C����>��r�w'���QV2G6����7K�6���PmWNC8x�ɿ&�&��.�(���J,�g����kzJ[?�%�?��)��a��"c��D\l��L2@Vވ*׼�۝ͭ}C���{����&s·���*g��ͫ4����<yD�����.�b�*mh��{�Zb��:e�6���~Sd�I%�L������-lZEV�]9�׬������
$ͿtG<�L�u�������W>��+5����a���|4O��b��6�S�6��(p1��mm���n���������m���$Hч���(;����(,�Gt�t%� �`�/(�?�!�O�
|Y���2���R�ߓ��"SA�"�y�Y��H�W\�nD?s:�Uٲ��VI��}c��k<�����œx��34 �'���G���S�e	�O��:%A(�e�Ϗ�ad�����I����'��*X��Fj3��m��^$k=�DQ�
��r���#�B8V��Tj�s��ӄ�G����"��e �}s����|��:���A���_n^����g��`w�u'b�[#�]T�}.���8!LF�~�w���J?VkVY$���C��	>at�@=�?�K}����@Н�0S��u"��^.i,wY��:H�Ew����X@?7���F}S�s�����߫�j3�z!�����Cǵb^�,��Ϛ!��{ \����bQk�bCQc�?�Ρ�逥3gggm�+�6Q���O��;��}�-��0�#�u,p���NL���e�<�w~o�ogoߞ"c��4�[mx�s��(���)s��q�a��~�1O�� � )%*ҩ�jQ&<�#��'b�M~��oSԾg�S�D��O��qB�7�L�����!��%F�@�nR�$%���Y��.~z-$����
B�7�[쐜���^�w�p9s�蒗گ��?k:�h�	�"(���,R�˺�݉qSq	�����D��ڞo�#�ɏ7���~Ad�������q�H/'F?��G(� `����χ��[�{~@�݋%|[:4�I��
�e�}��1���KK؀�2C��8�%T�Zy�J�����k����Ƌ9���DV[:���dr8��+��G�f�P�����/��tBc��V�|��_���7�!� `<�T�Da��œ ���L�/��
�n�������[��Ѣ)��4��<e��Q����t'/�B�?|vz
�it��D�9�1�ݳ���C������Z�y����+8!8AU�Kq�'�1!�Զ�jX�:2]����m�y��V����g^����YfQ\�i�[���Q~C�qD�ڮ���y8�N4�JX*��[�Z�Ӆ�?v	�}���2���+wU�e�f%�,��<����;1�QI���t��t[JAG�L�����M���O�[s�Q-N�ݮk��n�3-�Vkr{]O�3��B�)��X�|�%�~l솧3������N
Ɏ���
b;��8�Q;Z5r�*P�N�L��
�X-��;��[�_n,�t
%8����.�)ά�����s[�\���"������3�����"����,UȺb_��|��5��z�zi�s�BN	�I�M�Y.J��&ѵj�@r!h<�����~��w�c�����q�����)!�8��� j��/��	��\��q��a38p�sO��c��Ïs�?��4���]���.���G���N 6�-�ٺ��8����G�}���
/����ho]��)"��r���zµo�+��Gq�ͱ��Qv�X*	4vc	\h�2�@�P�1������ ��  ����$�;Z:^��Y�����������c����"st��{na18�`O������x�8!S�Ƣ,�]�=�݆����I2A��|@�ok 2�~H?����>���1O-��Fn��=�Qh���jߵ\.�o5���ۦ�e��Nv���q�W-,<��nsd3l����C��q�]n*l'��@H�gu}�T�9��e<6yN����� "�H���^׽8�S:c��.O���1�H}�,��mE#�|��d�������]?/� �4��E��QƝ��^� ЅD;�j)�ry�!X�Z��v����0�!�+h�Em<�Y){�+�h	鯫��$�&^O
�+È3�4$p\:[��ؐ$@_�?6��6^驋����b�҈+�І�}�C�.Q'��L�w3.�I3�b����2��7��C��2%~YX1������- �C	i���`|�[�m���7�u�Dľg|��*0�8N��i-���X���]�8�q�w�;O��|���ȩ~���Gu[�d嚑�֩�˪��<4_��]�ǘ�l��D�r�B���]R���_s��V��O�O����;�Ps<���96�xQ&��J��Flk%J/6#����������֦@����W�I>��S#.�b9�K��Z���@�w�"&�"i<j6���Έ����#�_-K�e(�!<��s���+�?N\��� �Zqf��6EO:�*�*5H9����� ����c��U9�~�%K;��y�reP��&"Ey�6|�7���>�mJp~���s�E�ҥ�ќ������C\��+.���|��߼��ˋl��j��Zd`666���k��k�,@�I3՜3	9������8�l�E�~�<ٸ���m�\t~�X� �ȮϞa����e�^Y��	@��ͯ'�j�ץ�f}-��Ŕm�xz�<��АY+�CCѰ)�%����v������1�?q�a���{��аU,v��)���z�D��6���Y(������/�k���_!���K�Ֆ�K�X��e��خ4�xb������(�%�mg2l@�)zf�"= 3~�-\GL�]2
���	�MM�?U���C[;�U�V#{j*x�9D6Y����r&�K�tY��$f���C���A��j#��Κ"U-�j��>��}���°I�J֓����UB�U�ʳ�b-N�?��������eN�jZ���>ï��(W,7�s��e���v^�Z����/��<	a,5�)�KBڐ/��E+TV�S1��P�i�G�|S4�l1�����^�U��~q��zw͗Wqn��1�T�������q������K�(�~��Y�f�2D��S�g܉��yK�"O�eqpK`�kT,�����B#@܉X��
,�2��J����~�ꨜO�H���O\�����ZX����ww�ϥ��LbA���s�o��=�a�"TV��9�i��u��{46�ɥ:&��5�[s'M������B��Vv|�9%���M���T3�Cp+
�`n�y!Y#Vi����VSJY���I9�6�Jh2���i�{��R|?�R���TrY�R��+�@k@t��_~kC�����:L�x�T��Ed��$�T�6{3�"{����2��M�-F'p	p��1^��8�
�Ɲr'ދ?��į,�j�?�쇉%�[���yZ1-�n�vq�5�cG?�E���� ���O�o��c�8�J���Y�A�-��O��g�����Y-�����FO�g��3�_[ұ���-��⮱�G���5�M�D@G���+A��E�k{�\]V���]}�����ﰌA�S� ;�	�n�g�����L��l���I�5�6�=ܔ��!P0�,��zEψ�5=�r���!��B�X��V#����.�6�Ȇ?:)����N�j�9C���L�+�`â@:Mğ�勜�2'x�װF��/i�Q�%w���떫~��0#���?��x�D��C�8:L"3 pB;o�ċ�T�N�$I��l��~�����:�:	��S�/αw���U������ޝxg�9�T�M�!�eE���]t}�h���N�z@և�î�*3-ZXO��y���TR"u��+��ϲ�É�!��j�=�@�EՎ�����̴�990	o����3+����x�aR8��yIZ`YtE�C@0ʤ��	���ʖ�%�K~�N��GP����Q��L�*��>����C
%/���i�v�?}�O<GF�G�B<�6sNTK�F��g��[}�����2�1�0�pYm.*2;r&!���X��2+�A�!um���V�'�j`*�{��!����}>�/�U{�w�k�pb�Q�G�G�v�r&RG�z�bڳ����B+�E�q��G_���Ϸ�#���H�W#�w����^�[,m/�癧��΍��4��S�V��V����t?��ٴ�4�k�����
u'K�>��@��5 Ǡn4�`/YD�-k��Ӫ�'�u� ��|�[�T�}�J�c����咂x�⭰�f?�2Q�An1��m��������g2i8�[�i��%��f��e�HgX�)9匼�*a*�."�lAn�[|��µE�/Z=�B��;Z�/H�X��A(�X�}ϐ��+��|�2׹׎�T�3���{��N��\� �5%$|'�K8�����:{�tl�:e��'73��rM��
T�]�Z�'���Gxnl��c�I���>�n�@�&<�e���+�d�9�Y&c����Z ��p��<�=�v{)�0��A�:��v��i�cOw\���$ɽZ��y]ޔND�s�1��+ l)[i�s�RaAh�_ݖ�t5�;���А�Lٿc��f�'o��h<��|o}k�`�Iʑf����x�W�:��o~�M��v�'
�S��m+� ���$�V�(��o�->͵�W.���M���^��I舥�ӶT�m�E�J��{9��ύ�������(l8	�c�(���hoBD��kS1����:���QE�]0�?R�2^zbv�Y�'�,�ig���F7�x���'�%����$.Rq7Kb��X�!q�Vŭ9p����K��w�%��Vf\�g`�џ?玐}��/���"�>��+6G��28

@�Y��ͮZ���*�Z�
��7,Z�:#D��Fh5JMq�ۺ�C�]'5���)�iq
i������g�n��և��hOM_�, �BE�	(�$�~^���#f��w��?=�|�t�m]	����G؀gFa88,��!� ����'T�_.w^/�O�q�WB󆦃݃�h@?��F�sP:�b{4��i�a8�e�\�v�l6��gB.��h���&z>���Eou�����
�7����\(��|6P�r`�DcD�%|��w��b���4]���LD�e���_oXzo��Q�1���>0��*�-��;��/�8}D۠��Y�8�yi��s3�~K;���v5x����<x�o���Ѧ���s�e�^�|hv��KȬ+R�>�=��w	�7��o�����Dl����Ϋ�V~.W��\�)���8[��?���MY�Jn|���yf7��$�;ܘ��;�S�<~
��%�y�S[����l��*w����r}
t�f��L���>"������@}�����q����+b��?�L�I>����ޣ��4���������4c<�f]`��5��$0+��~7ncq��	����S_:�cz���:�wu#p�X��"�W�ܮ����P��스�Xڬ^�,��1DɓG2�M�'��y�5����J��7��8aT %��d�z����D2�b+�Ӻ.�NR�+?D0�3~��c��D;[� 5N]1E���.�ü�dz��HXl2n���`�2aС�j�����JT�Mn�/jl�#��#����&�|���-v�]�\��.V��qAi�N���[HV焸�e*�py����pp)�܎���u�k��3;������A�&a�����=��"��0E��\���} 2E��b���o�����z*���{�w�����R'���D�z�=�R���\a���"?�F�_�y�̿�[w����4	����3�������Ƴ��6��j��f-1܆L��F�b��{c���ȫ�!��I&���}�����VQ:i�y!�7��K��Pex:w�gT2׺;�u���>6�(����CY?�3T����ě������i�*�0��;����e�6�&��ˍ���H���e|�J{��?5y���PL
j36�� ��LHn�u�[����m
� d2��Ҧ׾��୐��X-<M�a��<)C��z��y�/�j�� ��͘��u��F1�K���Ӟ�r�ş�@�: �����o4&���}�ǂ֐�~����B�vŔ��{�缵��*x��!/~m+�n��Ɣ��=����"GZ\�z�c���{Z�t���(`>Z؜9��l���X'�G�g߽;����k��lz;̐��K����x���K�V�r�Ҁ{��gV9�l�mX��HR�w�uB��<N�-��sv��XS�T�'U˗vN�-)FuX��	��������L��}���@�ح��X�Y=S�	'��"]2ŧ8��|M�"����S�����R�����uX��g�[[����.�m��RS��SS)�K�,F�+lpY���&6�LCe�{��u�����nɃF\��V-)�w���I��c����Bj��;7_"��+��,��þ�s�m����]�7�J�;����bx����&��Cn����l�d;���
,�f�G��T�ΐy]]�*���ukMv0uF�#����?��I�U�"�]#�e���x\����o���i؄X�]��>5��������W�E�m_K��4��tw(�(�H7C��!�J0��tw-CwHw0�����>��7���Z{���E-��̇��B7v�,��K�)�YW&����^�1j�Xt㕃���MX��SYP�� �m2��u!�e��ǋw��ҒL�l���-��``�)Ӎ9w��?�LqI��d4�hil�Ol y=�ZP$�\�b6��Q�%9r�S�$��]��nM�Ǯ������ᙱ��A����|�ww.�h��b_њl��p�p�����D!�G����b�o��^�}��ˠ������ڍ�QWp��Ɏ�b����h��e�� �ɟa�q/S�������ɤ�nM؁��K�������;bk���ŗS7�Vi��<��z�P��֕&���:Ga}��+���T@@��<G�+V.�jgp�{����������h��٫���ƨP�o���k[�q�&z[�A�G0m�d�f����C�f�6���05?�"�5�X����u8���|]���Yێ�ZoF^�ӽk�Y����[�Bٺd�s���^���f�ٗ퀈�v��6̽�Pa�� �}�3cq���ǐA���X�J�ŀ��)v��DIn~�#�����,�xn.��ڰ���,�?3g�7	��J���L��@⡿�_�����r?��"5��y-�����t&�1�N�\4^J�����a�k��5����:�qn��Yp�T�
"s�3)���zJd�"�u0�~)���X%�θtF��]]|��ߙϭ��8�����[�h�����[��zogs���f��E�M<S�ڎX�8tĶ-�X^��v�D8�)v�t��}�>�|�˖�)�DltJ�ls+�Z�6t(�g��Os�����p)^l�P��F�/�_V�ُ)�цz����QV��);ڙv��\�Vux"4�:p�U���%4�{��O�n|��sW-�L��8v��>����-Kr�A�N`?=�ZA��[b�)����U�����U�E�깘r����:��d�ȐH?�-ϩS�"��oz͐�>R2k:�S�_&ˠ*J0Ţ��{����M����]�w-�v��dOi�BMU**=y+�.����ɗ�S���R����Ź���c����+�ִ���̆�؊(�Q��ހ���I��>��W9�V��b�F���w���Bi��m�y�٩U�*�d�]���v���u�D���x��+�Na�4黉`"��j\�mT���,���kѹz;�dsTmYaI3��k*��pQ�#��ጨ�<!��[�����������)��>��(8=�	�;���Pr�%^�݊X�w�ze��Ӭ������D9��4�[o��e]�4}ziu�I�V���.�/�3��k��u��A�\w뷞i�(Џ�O@(nq�V	,ߋ��<�y���z����"��J��� �@7#5���N�"?�%LO4qf~��P�+�?M���Kws �f�Q�񨅖��ua0�G�1�����Ywh�-e䇴���V�M_�ZG�(gs0IT��z��.�@��-nΎ9�j�_�p�ϗ�	���,��+�]G���g�����e��Z �|Q� B<6R,�;9�1�/�8��70��T�@�3��\��2�m�Y��f���lܹ+�uY��ߡ��3���>
A�^��ʨg.M��Җ#�WZ��	EW�8Ȑ����t�g���4��x-<۸ڣwA�Mj�{�62\���;\���l�{��o�)3a�H��Ǌ�)�Y��8MÛ��v"�_��O��~����|��t1������"�t��`ğ��R�v��E�$������a{�ML�Vw�w~�rc�v�,��=^n�Y�I4��4�34H���!n���#/	n���#XI�gaT�Jq\S4O4�һ]�`�"IX��zq�*�
�-�<g��@�o-fd������r���~�wP"�
�ّ-�N�
���h���eAJ��G<x����s�E�E�(�O�Sϴ��ظ/Y�%z֡M�'d��K�?��=K��ȑ��I��F��\�<r�32,҅+*�#k.~P=�G�K6�cT��΄�4��_jM1ף�V3���̋ݯ^b�u���]`�GLg���H2|Z��gy��L�.�̷��n[g�&��SY�'�;BnǠP�+1c�!�pXP���\(���ys�%qT;�k$��Q���@�6~m��B��R�J�V����ytϬa�H%
����]�֊��0L�!.��ʏ��/{�V`ex�$�hǤV�C��L]�/5�'>�]%ÉF1���?]�:��d�=g�c���>k�.��z���>�J�D�b����EM۾W+�h���P��S�Av�[+f��~k�^KYCC�_uaƾ}o�mgh�! �P���1~="�����Ԍ_��� ؇��5~d�F+ eo5�a�f낢�o��hm����+�t�L=4\=�<��B�w��i��߇�-G��2�Ձ`1'3��`g�����Ƹ�ѩyk��R}Pa�^v��i��5��n�ݙ��v���Q}݇��{���Q2��_�k�	��|��矴~Kk�}Q��3���X�D�o�Fl���6�@��!�N��Z�����]{9��e�v���u?���|�w@�|��C�ߌ���D����n�"��}v�,�$��XX*^�
g����~'u�їR�\�S:�@�c3��H�e�E����z��Fl&��զ9�G钔-�9j��/��q�c�����X��c���|�0��o
Bظj\������f
�B	�7+yh�̭��v/#�s�M{�jt�L^+E�B�����e�&e��Fo�1+�D$����l�b� �$Z���� ���d��@�^�e��D���F���_%W&)��%8^ڛ��`j�xeo��l"ȡ��l0�:ɋ_2��t
�=�X���h�m�{0,/�n�g.)fז��@�����t�d}WW_���nA_��pk��) �T+�إh�e	�T.�N�3-e�)�<���+W�\�-A�5�WM�!8�yD7`[{ɬ&�@z��/8��e�@
���6�j��kC��XF�bP��u<g���e�h���몙��<;�З<��v7��?�jZx�<�<����/�b����?�%Vrn�T�`�%��%������36Λ9�3�,� �L$&'�=ݧ��Q^�(�'F"4�_���	�0�&��c������ի�.�#,8;h�6��}W��rQu��Д<�R�6"A^�(J#��\_40E�c7�DM��eO��cRcU��t�EW-��A����+�I�`�P ���h�K����ya	�yJ�Ek��7�U�6���,tׁ��9����8*.'ПL�D�`��B��R�2d��d�[�e�5j0?gS�@�\PC�a¿ֵ9��߲��W����� � �����gI5�wb�Խ��:s��ԃ����8t�T{v��F��Q�E��+�_���."g�b���qӱ��G���U2�s�o�����I>oG��yF�{�l�Ke4�g%��1���� ]��K��������2��3�B��P����UO+�cy:D;}��3�� #dG{{��Ӏ�r7� f�g�*7iQ���ȅ�~,��J�	���	[��u�\Rg���T�E�p�L�26��/�ՄH��R��������n��L8�GΉ��^�n}B;&B֙C�ޥgh�yץRz�"BH1_�O�_[:����J"���8C{V@j���叓���D}��� ��Ӊ���~�+^�9�pa<�ϼ��]�J\�2��U G��4�i {���j^<�K; 6�"i�3�+���uQ�7n����f���3K�ތ5>�����i�5�en��xt��7�:yV�П;�Z\�Xիh`��pCIcB-!VHb�_�M�	��7)s}�1�	��i{�[_���X�a�c7gO�������ږxũO�[,��߬'�`�n�14շ'�-0b�~�Ej2&л7�x.�,B�4�
��w��_<���qٵ�_+��;�d<�M�d�秨���_X�WR!�����X7 f�1G���4����]?T�X,��1z&�I�Ų[ \%&�PX���9�XWzm�q��3�u�vnJ��RzɹfK��3ď�y&q�̎�at���~�>��f��S�ꩺhއ���"��]�K�t�ЧߖC�>���G�L��Ϡ�=�R3Q8!�+�9q�=s� ���x)��F�DZ3�*��e?�9��7��4�u6����OI5ڧwb�:��5k$<&������;�#�6�s�A3tጘ�S>���u���ls�uɧ���� 2'͇��H�O=q�S*w���P��<t4u�V��[�h�c�~�ca�����~�GO/��,3[��Al�S��֌�W�H4Z�ξ����/�|�øU̘�ч'�S��Gt�m��|[#A�k�\p���~s��R�E�ɯ0�1�wmo4�h>��Ƞ��p���z�Fh�۵:�]>���i}�#����|@��,�n�}s@u�C�H���׼��fע���6�?��{_�e'aq�5���6���DF�S��Jkj�ܩ�QZlP����a�M�_��3%�τqh�� ���������l:[���^��nR%>�=�_M��m.�U��^Ҟ/�@�������ΕL���nz�e_�]s]k����"g!+���
��[]�/��A$��4��N<G��Z����47�5�I���T�]�u�i+	71mpc�F��鴕ʤ��nb��"��))�o�XK$�08�l��&-��a���D�斄D_�u�U곓={Jj���3\.�_R~}Рs������ǿL\�H�WK�ħ�%����L�����x�V�n)�*�0�$��8��W�q&ꨢOj\K蔿f��]�z�P��!\�ˤ�P�u _)ꅊ��("�y�Q�.d�4�T@+*�5�U���3���n���EN�/:V�W7���A)���E��u�u&�����/Sj����M#�n�rIg|�:���H�ط��\�y"~�|X{��*f+$�YqA'O�,���k1�Aǈ��nSs��P�<aZ�KK�5��!]$^�\C�Ь@U�ή\�w�ӥ�r�#s�J4Q�- $Q�|��|�i�9�g Oo���H���{F���4���󶇷�O�bR��m�ƺu
��/.P�Bo/����G�����֎zb|:l�0*�g�S ��s��54�ӣob�U���L� ���W�������Ӊ!��3�!�N�.�E��(��ل�X��� 8U�}DW���y�Z[���I'�w�
{��CT�<&@8v3�d+m#�q�Đ��9>��<�Ӹ����lG�Aթ��q�NcF%��2����å	'~;���U^X�k�_ʶ�;��ҎFN����^�=�u���U�,������YC��<� x>��y���Oe[C��%m����Pf���p�}p�C��eb� }؍<ߒ�+K�>M^��D|;r��>�I�	+;`R��Ǔ[7咸����p���j� ߡ���`8`�\�c�h�^�,��^ ��#�'��g���c��J�hm#d�!���f�8&���ws7�v��6�3���<ǫF�E��߀Q�:�S���ԇ�W��:C�y@DnBDS�2��!�/J&х�c��1\��u�rFl6-�ϖ��}n)3�DJ�O����q�699��OF��`kۼ��:%�d����ᇮE�OS��e����ɸ��%M]~�(��� �R�9�a�ɍ�EP�d,�g��{C�쭦�S��-Sw��\�n��D�z�R��m�V�-k2�;q��|t��#<g�x�q�xV��$)4�������A�8A��rC�a#f���X�0�v#��Glb�R��9�Pr'����7Xp�f��U~�5��[�>m|����"Po�\w��/l�)pA�Ԧ�UiM���H$vν���Q[����Q+�f�%�=Q�kſ<�	��<�An�W�#f�C]*{G%���f�ݠ��~�9�h$h>�ԛ<w���������|��qg�t��x4�����*h�q/�i��Ah����l�k��W��٘$e{?�_��^;uY0����	����zT�>a�G�,��u����ƀ��۪��y��l`��C#n��'C����KB"�0<��<Q��1Rˇǅ�c�1�1������-Q�J�iS�ߺ�v� ��~�Y�z�M�����E3L.��3������_�����s�^�%X.�7v(;v�U|
ԑ��{t���X���
ĕ�<�V���K�"���|�FogA1�qrW}Ĥ�"ݥ�ځuŘ�$tΚld�@����M�o���n�w��LۣJq�왧oװN�S�oz�ک��F���1�8���?T�id�B����q�r�Q�����Y��/�'��̋��H�Ot�n�>?���� :���_����y`7*ϡ��=~;~Cd�n�a� 0P��8Y���5�9��f"J�/�Ӛ`O��2'*%����5͚9Z/'&c'*�j�����V���O-dqq���y|#�o$��ܐ:vR���?���Yd^Kr'M�o��[�"n8�
��!�JX�p�}��O��M�﹠�󡥺)`��-5��<N�4���	)��IC���TUuv�4�o��pYU�������%X������}�1}.ׁ06,`x�L�p��T����#��ԏ�3��缅cM"�f��J)�./u�5�5b����kb���ګ��NRZ�^��ea���Sy
�^�N�9�.K/��#N
�v �sv_�I�T�V�:֭��ܯ�W�4p?��u� Bh����kx��7�!&_Xq�ȶ�odGs6����~n_i@?���+Ӽލ!c��E���LXp��<�m�eg�S�X��cn��W� Ue���?|�i �����xF��\eVC��m�O[�r�M�"�kv�D�i���߼�LX0��J���R+�<��O�\k���e1��E&=&���{�`;��0��JE�ޠq�6ȂjF<��k��$_�n�/����?�]YKfO����ZInx�(>�f�e��}l�y'�;SM 0��L�}��oa�w��N�>nQ4}��mDl���&�^C
>�Oؐ5���O�L{*$��qy�]��9"u���PS����M��z���TF
���Z�)��VC؍���~	o+*�=_b�Z�&�u�Y������ȗIaэ���E����W^��ą�80[��vf��K++ת�ũsv�dǙ����!��������ϢM�mf��vV��"�	����=� rm�%���,�e��>'��f���[Oc��:d����� N�;�BWz���Ɛ\]z�$����m��k��FO=��Ut�{�O��}���~;NnNN`�򌞁��WM!ە��)�O��Ά}9ӳ/R��#H�⾺�q�����:���N�[����>����V\���ydY�9�%��JO7OHc�m�ˤ7&g���p�o�l	nIx)��y]���Z�Q���̿}�����(1��l�R��]j���ׇNn�DY[{�g]Ͼ��%]č���)��}@U�NP?H��`��hiw��=un��t6N�ߚ��Bߨ=/���x`bܷ��^�UX��VX#��\U��@�ޏ�zzFy�����̴�D�l_\��ݭ�:rs���b4Zx;�ՠ���k��Q���� Ib���aO�[ݬ��,���p�oK���>^R�(� ɏ�$l�G|�>�]�!�e��j8����}l����|������4gn��9��3�4��3�.�{#t�����L�>K�XX�C�]d;In@����V'�	����D�ga_��==�;�	�`��Zu�ob;�/s���?���ZCu�;�gBW�����u�J҄���zES�LB�\��^#,�� �W���\lQ���"�@�J=�5�:=��̭�f ��� Ŷ���2uԩ��x�j����~�y�9s��yZ����:�z���<'햦��W��/�b�%V��Ĉk ���n�IS����x��Nn�Ӑ�e }�$�K@�4݉�'�q��f��R��%��IU�ƫ�bn���T���S>�O�@�ϼ5Y��E�%�1I���Q�S�偎^��G���-��=�-��zh��i��ë�ɤa��t�D����|a�lu9�FWM�a}:�?8}�E���Ag�=Y�A��W�6V�η���ʳq�8PV/�&���ocTx7�_��}{������ud��8,���'�n�U���?�QW�"OoPA��`*�	{���K�u�t�a�z�?~q���h@�!���/���Wd+��V�bm�K[|���������r�0�ڬ�G�e��]����O��妿6��'�n~�X;��Ya�'e���q�����8u���
t�M�yH�\{�C@��U��C�'���;7�S~"JnEU!�էK�����K�~"nn*2�+�@�;�w�L��j;)��=?z�9�E��@@R�`�`����|Nn2j"n8�K���:9d`��;9��-������a��D�א�a��h��������N���U��l�"��C=��ɔ0����%?����L�{}��5d�G��.�N��|�J��
��տ	[�ni3�iC���?t��%���"���s�����g��SL�l&kf�L�uw�^����X+��w��V,M�F!�0�R�Opt�*��>4l���?~f;��ϛ���9��D�����R�s=�Î4RS�	6��r�m���3ۅ�>=��=���GFs�r� mʍ�)����e��#q<��Q���W��
�a=߇R�^�i�hQ�.�9q�(H�M��1�էGD��#���q�7���4j����
q���_4;���,�M�c^��	�������B�XW��u�c�o��P����@����EՓC���w��	�8ύ��L���~��!�����w�:,�t)�p zo�k1���ԅ�g���=e�8�������G�xC	)�&x��-��5 V�����-��b�[��j��#j����O����1r7[�s-9����k����^t���W���9�P2���|w<k���-�,��r��Ρp�
cb�u^c2m@lFnm�Rtl0O	D�R��"�J���RO�O�:a��B5���n������
����̠�R��K�I�?�
����E���a�<�_'�����l�V�:[4����.N΁W'+����|<�J��VXd!p�$���i?�������?7^��a�h;�yØ	�����KG�=�����*��_��8��P���u]�[l��7&h��j˶,�赯�k�|�@C��� ���s�ڀS��|U^n��h��u5��.��z!��I�ϔJ�n�{���6��Ɋ����p�lY�&O�j㖶i �ɕ f���5�|AH�N�v�+��O�C��Gu0��}��n��A $77TEQ��;���"H�MT�V���V�@�����fT��sby�#�D��}��4�yݰ�g���L�V���5�/?&ό�Km��ߥY�m�Q�\��b��P�'����6��l�^څ�t�9�`2V ~Đ�+�Z`��LL՛G��t<��.t�ĳ�0����'�$Au���#��BҚ~�1%�xt ��膷����z����i��g 	��2V'��|[��t`UU�.�OTfO�s�5��AV�tC�ɣ�Bg�a$��[�ĨK��I�12D��
��Zl��a[[�To�q��u|u�.�~����R���g �^g��"nڝ�L���M�8ν�$p�;`���a�MT��o�-��|u7,���4:�p�-	��<�62��[ի�!}�> z��I_?�:����4��q���Y�>'�qC�y(�v�|'�rUͭ�A^�F�:�{�ulLf�t���W�1J�� $~��X��1\?xp�"v��j����K-�Oݾ:e�Q��.�ڡ�O�+�EzD��0tG��T5�rc��-m#�	BS{������(w�#����+�ڰ����]�9"���Ir�l��S�r߻�ð�Q���݋x�4ma��c�����^�R_��
�����@��'A�MQP�r��W�؛ɛ�N`81Ǥ����)L����L��5V���Y0�Q�*���B�����i�R����7��P�N�bf�>��?$M�> �4{�z��~��a��X�e�����/�m����Y��I�@����X�ƪ�,��q����2��y���L��k>]�����(}U4��	8�����JO[��B-�f �h�e;�"<���E1V�-�)n%Ȩ��$���d���nq��c��/,&�*���6�޴"q���ި՞�-Bx�n�g�\G��m�啕�D��މ@0�������i&����¥�Ԋ�bҶdʔ��?ݝA��ѧi�4I\��B���˒�g����z�$T�p��23���#�|��i���EG0S#�������ՠ��H�J��1;�i��by|a����i�e-��]1eZ)1����ˌ	2gR�	w��⭍S��k��Z��f�R=sh?�:�M��:j��)d�,+%x��qr�d�N�i=�Z�k Vg�ƍ�mM'����a,�Oد{�3�n#g���o����O��*���ƀ\͆�X>W�7s(�Eq���R!��C��	�	�N�F����ʹ��H:9�0C�"�����i���zVE���=�)�{?lh�5��9][{B>���� e~�>� ~��y����,VT�~�F�����X��T�����m�c|k�OG��i�4����RxÁ��;5&|�^��󎟃��Ao!9u4#(�c#=�1�ۏ(�Y_,:sE$�_������7G����f��a����2ls�!�㡪'�nq�A�{v3f��TG\�/F<;�\G��%��-IQ��)d�`N��<��ᗙ�Wϛ�yA9��A�ӥ��Mr���;|<N��B��ט�_���m$/g<f�Wrjq\��$��]�Z���s-�#���`TU�f��m�~�9��}�gv-�Zp>�؎C�F,;p� w��{>x�'�)t}rR���C��c-CY,�]k�lh򿳧[�.�&�D�pE�]
?��:�V�'���pY���Nٜ�8{�e!�+��.6�2��I�|�M�3,���>[��C�����a	>i��ƈʨ�4�#��`S���/l�~|q}k�K8v��vꗎ��w����x���ү���g��б����	C����iFJ�^�GtG9rF��1��_T���J5��o����B�ޙ5��j�V�:I�%`���������ϫ��%�^���Ֆ��f�����Q�P������J��I���%7�5%厪�[&�?K#��Ō��m�*/.bF��T�����YX���}YP������;�`!~���g]��m��ƺx��	��d'�#�)������Z���x3L5�;�VqB�s���.U���Iڬ��� ��-�|�Ì�*R������{����'Ծ��~ؤ�-ƭT�p���HD���x�� ����s�!�+YZ]�ؐ��^���v�i��7��c3�&��W��-��]�Pg�@k�2���#����ϷҬcf%m�����f��1_Q,��<����,y.+����⥧�{�1��Z&���ߝ�y9^�q}I�e�D��~��w������c�f�S����� ��n|F}���v���a��ܗS���l=1�������T��&���kT�O�4S�/;b��y��%�
v��7���wI9N���فK��y��Q}μ�yv�2�e�솾S]z���~N	V�;\b�
m�v��g�gڻs���cK�x�/s��:s�e���MG�0�< ��2;s������W���W���:u/ާ�/?cB�$�[�<2VL�{%{,y�>u��n�ҽ���p��sxz�>�0��L0g�,�0�aԽ��%j\�L�(���T}�+Kg����i���)�Y^���i���yHwW�j�]�����T��^��@�\���Rz��+k�cp�p,OGqj4���a��;�����4��;��ٷ��f��2~2�I
�DK¯���I��T����>>��j;BΚꪁ�?z�2ӆ<<�����E,���&��w��g���T�Q�0��@���CT�^_6�4e(`��u=��/"/Bm��R�)�3մ��J�ov��_����E�>�v�uݩhJz1�r�F���:�H��*�x�	�R"�,��z�9E̒(��shNT�E$R��	 `_�?ͨ)�E�����,F������{�Ҥ������/{<L�oTu_��/Zm�<\bG���1�>̿�^�)wu�Z8Z��)"*���Jz��^�W�K�U�!����Hvo�������Ěx���[���e���8�d��2ƱI_/j_i[�Qp����)R�8uX)(�l�����~oZ7 oF�d/$�B,����[\cP��x�Ō�Q!�hE�WdP���8g��q~�W����4�\���Z"�����3%v��-=O�~�k���lB���퉒�-'n�����蘶���6����J5��1գ����Z�gUuf���M�%m�q���r�<ew*��iAVQc����͠���B��f����cWU�J�Xi#��);<&�y�I�X��tD:��_� ��cW�W���b������#���ˋ�W�{�ٻ�e�B��΂���gv���5�a���I���99�o���t]���	gH��=':gY �G��e����L��c�Z5ʺX�G�Y���������Z�,�[p'.����|ƿL�r;�y� 5��V�r����� �Jn��=]���z �/�e|��^y�0>
)"������Q�ajzt�`�7�d��bNuz7��38?y3F�"a	���������H�d`3����`��b�g���_�Y�?�~���#�Vۻ�ƮuA�%o�x�헩�3e�f�o�ќ��I�9c�e�j�HnϤx7��}Xo�����@�0g�w�OK��[[t��G��B��wTzPI�G���p�����,3���q6���11uÛ5�G�h��^Um��D�O�v&�I����d�������+��M�;����'HU>�8l��sZY���c*�e���eV̗
(����ݿ�� Ě:y��ȚfY���Ƅ8:=�LII	'��������kc�� ����]Z�6�i�����l����l�92rF`��ըEZ.Jw7�� h��H�eM�B��T-��f��=t�-�9"fi��F�~e�qӀ�ƸTB�K"U�y�dH�dA�[B��?N�k�4c �DJ&�b�uQpH7!�n|����K�2���ݙf�RT�,�
C�[����M�K�f�@��X������m(�8�k�Sl;�MxX� K��[�m��N,d��_H�q9���4|�NW��/AJם��P6M ��`�H���)�DoN��d�_: �q	w|΅�����T2�jQނ7f�nf|�7�΢J��}�%PG2wW2gm��L������hL���Hr%�����q��e�S���U�h���Ì'�JH3�+�����0�Ʋ��R.tP�nFvh�!�C��dv�����vTw�xz.TpGY����JV!��c)����k]����ɧg�O�mځ����"p<c�"�qB�.��Z����4�Y��G����G��a����_�%� e���9-6ş�ڛ�
�fU	0��<QW�ꆫJE툠���o�U�\�K�����%�A��+��P$9��:�㪀�{�r螤�yz@k}TuR�AHs�C�T�_�
^b�=�<��xy����+������4�N�2qu�(c�����볕�Z��n��}���h�00�}���u���.M������48�Os8�\8D'�؇�~?1��q�/_�~���l��ۜ�G%��_lE�y}�l�2uv9kn��j�`r�D����k�.>͢�4-K��;��cUCm�w����6�ru�F�hZ���K:<�g?��՝+��N_�n.���(w[v�J����v���<[{<V���ˣZ��w��t��<@��
Z2`�q#z�d@D�t��D�X5��hB�}s]ԊeTM-�a� �O%U�H�����Zbr�o*��,��;3��8v����.�ف��+�o���ͥF��WA��+<��͂�u?Y��pVLa,�[6(M��u��lq�qfy�WV�E�|�Q���;�}R���2��=)�m��D��u�i�JI��P�i5�g���
f�poջY&Ֆ���U�-AK��/�/u�B������L�O�A����6���P�yF���N!,�RS#1S��?���r���зt|�_������8F��;�rַ��ݿ��(�V�[ҭE�����:���2�6�0���u�h,����ٷ��n��l��P3f���ƒO�㬑B�������w�?;.,B��<�#"n��*�.Y��T�t�`��C�Q?�Ը3��+�Q���HF�sO d�����G���Y�����s�Ұ�/������&d��'G���B�M�[�XgG�Z��.q�g�l~���k���@���%���s�!?
�����vZ�y�42�
�	��p-��T d]��R,���/-����~���Ob%�3�K�w�z�jcv����N7m;b<��j����Ko�����-0�Mu9��#r��G?���OM��r\]4�% ~L�w�<*�@�m����Ak�V[��WS�,���������z�թ)(��%��ε� -�����^����b'�O6��C�1��բ?Ƅ(�_1�G-�r�rFV�7�7���$Rʹ�����n]p;)���\[Fj�m�e��f����+)�}Ѳ.��ų�9�������s��:��J�M������_ �����&���Bl�}f|Y��U�s�����m$�����֟�)�:�dQ�t�����Si�kOkn����$��/$L�V��fcq����W���0GbN=]&o0��c')�$��8���M�,v��)����І�%��s�H��}��r)�\ո��0{�V>�YP��@��W"#2��E55ZTɪ+x��
��Fv�$�S�E{!��b��)���Lj�������H�k���Alķ�O:ݫ"K/cJ,����=Żo�;RuZ�=R�O��IM��K��t_�/H�nz�Y;�X{�=My��>�q����A����u|8�<s\><E��R�c�����2�=��;�Ѓ�5�7��8��hZ:��Dr��U@�܃��	�#YE@���9s<�w|9��w��8����K��B�!��{���%���d�`�<*ߞ�]�<y�7v"��瞏��nrq"���.ך�v��8*{��*ha=-�Cg�J�$�^`켼�M�3?M=�z��_��Ϸj�
'ɂ"g���R�\"x�$e|���N�n_��,Q�v�c���6F�t���v������R�_
��V�*�k���夢����e��0��I��W��"{�����He܍�����$g̉���zs1�b{D4	˻!o$��Z�gn����rf'y8�2�2ꮗM+���\6Ag��c�]�s���K��[>n&�E����!+�}���J���.�#׍��֒�k�ks�pO۫=�S��Ӫ��-�}BN�j�\����[E��
���j��&~�b�R?�{s�:��Bp-�n����������z�ҾW��)�W,q#,�O�S�e��-����;��4�r�����6����%!�O��9]��4�*��/�&����@l��q[l#��Cl��ݓ��8�:��?ͳxխD��'�j��;"��&��Vh�l��p�Ń�=��~#I�;�	|E��C�'��}\������S��t�K�ڑ�O+����-v�X
{M��B������/�����N��r����D�2�Y��3Z�$���	�w�� <SQʸ��u���[�$�j�
J��,�o�?3�nAڱ�;�T�Z��<�����	d6��}?��FOD�Q��ȼvw���,�9"`��g+ӧ)}_2��n�A��[_���=P��pq�F��v����Ƣ��PA|�b_�+�vXPY��V��9�Ȫa�զ�����8�W��������ۢ��#����`}�qJ�Y>����C�CD=7��o��B�� ����1o*�]��t���DO��1��k@����@kW{�<��㴕�f�
�:�
"Lc*�@
K��k|h=��n�n8u��{�spe���M`8��#"{Ǻ���=�v0}ܯ���&Z=�č�?kbs�	��ƊC�<��㩙�tM�S�n�h�6���Mk7Bh���{�gͲ��o����ys�T�5�J%@�V�m�����M����M���O�h5��@C���S[H5�CV�Ý������[��nU�Sd����s��������k�GQC턣]Y\*V0��D���:q�;׶Q/]�IS�:������~.�ӟ�L�P����������t�ܽŽ�]�.��2�R5ǭ�y���j��
wQ�r�uvUR畄0�k*F"&)�營�O��5B+��y��v�gz3�{��m�ذ����]wx��Q���2Xȿ� Q�J�'A,���خ/%�u"֒n���^X� �p���ŚT�Sx�4�=>C
Q��g� �ۖ:V�a���W��k G�1qͪ���OX\}gg���<����:�Ƨ�߼��S�]-��;��q,���Z�o���F3�F�� �t��ɰ�W���%s[��ZV�j��vǟ���Sf���q���L�<~�h���FB�+X�gq�c�	���8������du�V�A���Y�z��`�a�U�/�c���*k&�T ޤ�n�v�ƍ�*��G=�:�o����XE����[����[���� | ���vw������\|qa~�_I�,��.j<ꌋX�V!�@�52��_!7��T�F�yg4bF $� ��X��E����:#�4����U�J�Σ�N!�_7L�H\I��Wz�!�U����]aC��K��lS�v
ϺlE~����R�Xw�A��Xڃ�ލ��=P{���8�K퀸C�".C�b8�=V������7�����e�R��N#cc����͡�1܄09��l���>�����a0˽SZ�CmObˁ;�0B0�
8���h#%'���r0�<]�4B���imc��#���p��+w7v���o�$d��Hk\$���4��lzb
�Hf`~0X6������t��sb�ܑb8Hs��.l�������)�����y���r�9P��.�O�Xy���bC =������"�ՠ�R;e ��P��֝c�5��ߚ�K��'NN-\���R�D%��D]�Z��W�0���m�J�7$��Ax2V� ���(Va��{���J���FUUtL�o��[ۜ.�Q�.�ETc�{NKi���G��HEx���t��	�b;�ի0���A�X�Z/�hO��=;σ�T���*�@�	!`��/|���g�gөS'��}����OT�$�={��|�D9g�i/�1�& �35�H�ղ�Onj0}�����jn�[���1���շ�U|7M�d�͔J2bxE��Q�A��o.��2�?ƅ�"�0�үʣZ{�3�'�����Q&��.`>�bd���^�Hd$,4S�e~>9��<rx�.�i��W$���YÚ����A�`��)+�q�c�9��秆+ʷ�\_��Ħ3��4��q,_xuu������0���2L^?��Φ�����t�u��\��|G5LQ_˯#�ߑ�~�),���z� �+œ������J
]YY��R�,ޓ�2_�cl����y��#(��.��H�u���?�p���ƚ�m��,q#�[��n�v�[�k������!�����w?37��U�Y}��^�7����|׶o!^�3��}����@��B�-�$�"D�£{'��J���+W㻛j\�L&C��X�p���=J��'3R �8C@���I2����3�B�� 
Dֱ�)#�~}��,"M��� 2�bw8m�.%h��%``넴e����+����Z�.�'��h��H(�\��ջ�ԇѸ���4�弜����~��Y/,�Q$c#^H�0�@���u��;�� ��f( ��je����X�+y�>8T`ِ>���g�`ƪ�8�Dc�څK���`̢&w�sEe�C���o���u�Q���ҍtki�8�]J�nͤ̃߆�)9�6�������0�a2}ac��*�F��~.��3Xe�BqI�T���LW�魯ٻ%ҷbH����G�<},u��cX���)�ѥuT7��G3��Hncּv��A?�S�a"��#=HG�iӹ��b��N���o���Sx�I�&�� �$�dn���Y����o���Q֋��@��]�lxg���������/Ϟ9S�R��ªX1=}4�<qB����_Kwfn��u�{���c8��m�X�BdT+����g�W��/��~$���K�w��&@7&�M�����ĉ3K��8��W���$D4��a쇄*���'\k���9����;�j��vN��Q���o4�rb��Fg0R��Ȓ�����`jI��L�y��ZeW�z�2��;�X�P����z�!�C�"uk� ��.~�ᇙ���.�U�� �����/��<���
B�%�6}�G���'�z��}O>�����&�_��:�Vy��#��������6������2�A�3C�\�`lr����*��ĉ��]�_�8)�J}\`�[���w�<cNizݵ?�/�:ݰsͬ��x5vY�;\�Y;��9�u�ر�|��x�6��i*������h��?�h3W�b���|q{s�+�n�~1*�Q���*"EuJls� D���x�7H(���HU��� }��@�d���]�DED �i�E~5b��(��2���B@|%��Fp��Ã@�"^�i�aJ}CǞw0J2K~�\r-�RGʉ�42N�Y�d� �Z�E��#�8�Շ�T�h���-%%;�ܫP�^+���*]�k�@j�~�&�/������+�`>����@��7�1͍�@$�����^�i���܃�)���������#̜�	���
uI��"$$N�U]`:�a��wh`��G�N)<]����n������M�A����x9�,���k+�����N���^OwW���`��,IKp�����b��;�����N"��K3���Wnk����Dq��{��Hzc�f�ci)���f����O��5��������6Ώ�Ҩ	�����m�\pQHixsF:��>�(���mb|Bii�<�.�.�À�޲�+��e������\t��,��77ֹ��Dͥ/r/QN�<Q<�䏥�~��4�h_/gÐ4�hɐ��!�L���<���8o@L8À��_���o��J�N'�u�-$�Ї��>�����/��{"�������r"?�Q+�P�Uw�j�w3����c����O��a�rX������ql�d�q-F�u�!�ꬒ0T��%�*���ȅ��Z
�f�G�b:�W�͔X?(��/�i�?��u����G�Y�����;T��>u]2��&^�G��:^No^�?׋��_8����/�u�*_�;Kfzb=9�G�o<��Ve�e����>O�߭k���5��p��Y$�Y.��0/\^p���>�T^Ɨ1�ƌ�������q=:���|r��ϲZ�12�U�Y�;��m� s��Ȯ�����F�x�s�2U<�v�^M#�!��̠y����#�k�lJ6�l{����o�:E�X��m�n�v|PZ��\��=U#�1p��Al�077���ٹnv�:%�@�XY�@f�b����"D�"���>�^d���W�X��Dh52�
r�	U�Y�v�I��H\�!�6�C')�P����Dbi"K��l�0��䍣��i�G"�"B3��,2�}�x�U�f���&��@H#%�
ˇdU��9�U 	醰T��m��32G��h��9̚�|�u%D�8����?6��H��8���Y	���@X�7�!T�8�D�ʼq)m���������mͅ�AP�-�`_ ���Wq�S��B^M�wq����0�1���+��h!����3������D�~c�\�s�^XI���r�jws��� g�Σ�7���y�=����U�Ž�|g��r�z�=s�h`
��4q�l��T�-�x�o_M�'�Q���2�[��Q���xq@c/�l��ޏ��Z��{�����+�P?��h��N[�ǋ�K\ԋ��eL��r^M�F&g��Ĳ����y�0�3^K��������۷7If���遇L��%&���>�$��eOw'��^y������o�+W��o{�Jz�z�*��(�����Buvf�X䎫Pgb�9V�0�?�|���?�����|6]�z5}�k_Kw������G�IS1H5��JbAʸ�K����\��㻞OP�Ϊ�x����
�"#�sZFͲ�/�i�|���c!�U@��{7U��I�L ��̀���\u�VqZ�@�ŵ�h��O�L��:T�E�9_���W����C����"��@�_����E����<���3`0����p�3��8���?-?��bLH���:}���\�>��jp�����]������C���y��#�X�ȃ�*=������*ߺ����Z��a����j3�2��1g�����/C��F���Ĵ���z�V8���5���t�1�}�vT79g���ϟ��훔��f��i��-�n�L�����D:$�EM�߬��<r�֝,�u��DO�3"ݷ��FD���Y�]y��� /|�?��jb(�@"*\�1?�3�cٹ���8�,R�	��En��*#��i�Q�
iT	�q�abt�J�(_Į�Q�0Y���@ə&ୈj��	�)�1�6-�U&����ձc�����{���:������(�Q�De+a A侍*Y��!�뉓'� �W�ʅw���V8���S��#E���e�5�`J�w���P,!E�d�y����w�ԯfF8��}����e��G����xƫ����]$�I�361>���p��s��}�&n'��F���(���h�Zg1?7�Ff�4-o�+�孝��Q�D��wS�N��@	V �P��Y)��1Gށ%>�I�k�kvC�Gӑc�Ru���\<7Sr�X�=ic	K�T�5ʾ��t�ђ�-�9�~�=�����z��������:��f�1��@����T�sL%j�J�P���퐆�^���a`��D� ��@�ב�!������{�q�H���Zz���L�}�ݓ��FO�������t�������\,}'�Rx��8�,��!����N��U7��`�i�=ƾ�~�'���+�S��?��B�������� M��#����O�<bxD�7�Q�f;&H F8%�={�x��u�a4J��j�NpE�Vq*���T��I�c�̭�i�M�׌,%�`���O\��B�o�#���q��_� �C��^r>Q��U��7?^#�����ʳ�[��%(��u����iL����2>q����E���G^�}�ˌQ�\&����MS�-���p��������<ޖ�Z�_H���:�I�a�_Xo��M�S�Ee���7Y.���������:�'�_�y[>.����?ʷ���&��@�ݐ�|����R+�r�3_Ǖur̒Gl�F^q	aq�i��V��d-�X�ީS�~���{��X�3m�n�v|�Z��\� =v���H~桿Ĺ��J� �j�J��w�B�"��HZ�W�@���e<\C"&���y�*#����>�噑�+�d����ʊHSd�[�i�N沽�W��,�(0�H�o4�;|D�:���򸮘C����B&��|���� +����F�t 1܃��CJ�0�^tb�P<lZ1��)T��P;v�L�<{�8�Ȟ����W0ܰ^�a�K)QI]�e�@/��؂H؃	����(<J_��p�Y�jp��n0���o��Ӻ��2V:��EP:�ճ8+C~4b�v��rj|�������J�k�A1Nkcy�u mKǑ�a^����_�M��kX��j�jy;�����i��&F;P���*���Z�ǐ�.� ;��{0�o��e�u�ct��'��ӧ�k��Z���>X��$��w��jO�@C��|6d��ؤ��V�Wky��a�ˆ�e� �j���Ŧ���9$U��������H�x�5�d���/�R����V������sH���<�ƛ&��QAݪ���P)�B��473F*�i���1ǐF��I��/�0ⱀ��Bb�����f��~+=���Ń>�N�<a,�h�1�3C+�ݯ4�n��@P�����ȸ��u�����Z瀿#�ߌ�X_>:砎5!�1�� jN�0y���@�w5e+���h���ZQũ�כ�u�e͸��.�.;���F���4���A��so��8Q��)l��:��F��39/���v��y��#~xDѹ?"nk�3������p���d�s��(����
�ڵZ+Mg^�q��gl$�p��D�։xQ�4_��a��7�����D�Ʃa���o\��O���"@��76<�M8�׿ÌUfM��k��Y��c���pq�cnU�W.\���Z?mˀ�J۵[���x���Y�>�0W����Ϩ���ׯO��-Ȩt(�I|�D2"��@< 0N&�$�*b'3".�H���DV�i��w�A�w�"o��,?�-26H5r���8�(S�o�+ӹC�]~U��״2]2D2W�ӏ45Vݙ#�W�˸�[���%���m#���wI
�Ah^$�S �B"\�ْZ�۵<�'a��}�Yd��0����ŉ����X�v��!Ś$�������(^�v%�A��y;�������5QC; �D�����ˈ����B���:ժ��A�gցvS��4��vQG�C���(�q&H���c8���bq���2"j�ibl,���|+,NNMa�n8a>mqN��znZM({�֊�s�i�������`w�8~$��ю{i}�2g��)�����ǰ�xGw� w\��-S:q�T��c���=�n.�c�b)�pƌ|�6W�TO���4�a�a��v�P�c���?@Z��_���xq\�dߞ��v�Ly�(���p~O�N����LH�<g%Su�G�I��~>}����c�?m������}��_�
F&Jw��"�R�=����C�H�`��W�q�=W�"8�)��臮��rjr�8z�>���io��|��/����ӎ�;_�Fz�o��OgϞc�xNf�]]�t���H���<Ʋ�.��2}*��W �#ƿs�=)*�vu^�c��q��|��&lZu��c=�6GL/3���s�1�z�󏴌9\&~����5�0Ǵ�9V����Exk�G�����~�Z�����;����O�?]+���ߖO��[X�1���}������[��_��bRޛ�8[�/\>�(���;�qm��e������R��0���[?�����7%�:����帞�&���f����%��u��-�
~�݂-�9Oj�0�s��oU	�芉3���[��8�*�ohݓ��	c�\XXػ�����G�]6A��8�6A۵[������@���z�W�WOqH��\�r�aΌ4�L�\0�퍪]7� B�8*ج���3X""�h��3�����R0J"%�f -��$�D\�DNX d���ޅ@MoY{R�̓��^�y�ee,#yi��^�I:��6��G&"�u�q3�xh���Ĩ[�A�	�Ț��D�T2$�@ܡ~��>��i�2�`��3UJt�`��3E|�C�s��%�������
�Ր��8PL=^N�9�؃����k��k׋$]G ̧Ɛ�@Xs0�t�Akt��}ô� T����S���6�=�]�J����6�H�hz�ޖ���a�<x��Jj7�K#2��X.������:Rbp��~�Z���)'FǊ!�(����1��ϧ�^(���փĨ��l��+nl-���ͮ�b��N�X����Ō�v�I�wn��]����g�(7������~:��g�҃�>���T�u�J��N�ads��v�k��$F.�����������i>�|��=�r������P�l`E�{��t#�
�bZ�\��1~��?�~�W�u�9̟=:�E��_�ŷ����|���3���\�9u���j�0��0���Mq��8R�1�)�&&�/4H��F
92��l�r������r�Y��{�?}�;�I����ٳ������s���n���}	�j����?�9�K���]eJ�ɜd>FF�QLF=_��4rH�Y	���|&V�|�)E� \�ܜ)���g�W3(�5 y`3�� ��.���sR��o�����u���"�}G��;�q��"��ǵBOY��s}8����4�yG��s=��2ޓ>36��k8+`(�d���E"�* ��z������:��&�8�E�j���p],��!̎�j_��5D��R��,�&���jk˷�s���w�G����b�7ڏp��w�ϻUo���Ɩo�a�������a�J��4r>��^�Hx�禚�qr/D����&Zɦ[�3V6%W~����ǿ�߷�#�wL��v�h�@�>h-�f��+{�"�:�����;w�Ar�ayT�P���\� \���'�~P 0҅�D^"?��A��M�@|�n�8)@B*�^;�6��6#Y�t�/R܇ᐰ2����<]�������75��C�k?$D�{av�8"Y�b�e�H,��L�����U�U(T��Z���"Ꟊ��/�3��jR�bt�!*@RB�s9�ؑS!���9*a��"p�q����]ލ%-8<1��Q��2ŵ^Nw�~;�W�o��1�0E;������)��.���V��Y+���W�( _�g����d+���%v�5�ak޾)�y�f��j���r�T��N�rem���4
�?��M���;s�͵MX%�8��Z4�Qw<�FNK3+\��i`��r��2f�o�F?L�JG����o������)�r�s�4oFsgs�D��8��=4X�@�p#��n�{S�뫪�������1�1���;Pݴn��H����i;��=�?�Q��!�,�f�i|���u�i���(�?Vp�T܅v��-�*��o�:=��O��~���~ƋF,N�>YjpI��S��>p,)�<u�dq��1,
��˨X޽3f�����dr3�ȍ�
��K��ų�<S"�
���@%u,�3�G�0Y�V��H��r�1��S���1�C$�*��ᵇS���i��<�C���2J��$��U0O���G�Jb%,���w���}n�M���fJ ��t>����@�o� ��ց�qs�� ���o�w�!��c]�/���Z�OXԉ�CQձ�`�ܠ/��V�(C�ud�����(�����.� � 0�{��xW��]ץU��k�\n�g95n��@�\�XSr�r�o������X1?�r�܏�up�p�7/��:Lu>Q'�[�o�V'uw/ڎ,"��y6`��oy�w�bmw�3�y���'w���իl`�w��)ԧ���-��+{���-�n�t���������������ss�#�����t��k�$[���Z��F`����H�L����F������?���B�;�$#��Q�87�Ψ��(����yK��ۼ�)��ęgV$�D� �؝4�y{�����85�P "\�o#1�b`0#�tZ��eh;#`��
3�@���aq/a_�32�Y� ��4eW��q�;��\��%b�w7���vLL���4�����?���\T�Q�s�hx�(��r�I�!$ͽbmi.�A�C�V�����r�Q>[��%u����x�Ȱ�\T�j�ڸ&l��DZ�+��r�����Ǎ�H�8��٥~M�����J��528T�tqO�NYb��DEo��w��k~�3k�C���Zm@`qwVꍽ�b��� ��&F% a>�Qu�G�3Z�"�[������zag--szm�җ�֊N
�����ŝB�����G��[nR�ق���"}���Z�M��X7�@��3*��o`�3m����2����S?���'~�3���;H��y�����/`��U����
�z¸޽{K���k��=Z�S�\�L�i�+�;�E�����/���S\����V�6�"�4���]�y7=�̳��;wӽ0qgΜ��{���F��N[V��s0"ռ��+�G���[{Ώ����}1��7�߸����?�j�`NԪdl �r�ձ��ZRIT�����w&������Zj�v�U�Ee�C�w���;��f�^ǋ0����@�33���|��"���8�k�y	�o�k"��$�0�u��N����F9��t~'�Y���E�zc���p���z�G]���au�`t��Z���P�D��R�$\����0�q�6��NS��v!~�}r��?0E���f���Ի��U�&�s���5��z�}�#����s._���=tw>����&��=만Uؑ ��-�n�v|�[�}1��>?T���~m ��/��/Lsap�	�`A`�ǹ�}1qkw�M}�i��Dj>�@t�����-r�aE���ir�:/�օ���A����ݎ�����yG%E��4-�D$�n��!w�њ1��<D��N��I��9�TKd�)UA���`<T'���M*����{O�T������|{!.%���E�!c� w�\V6aR�e� 8��C=ͳn���!,F�$S�HX�a\f_}=-"����)��/�N�PP���.��}�B�s�&8�¸ XY2�5�����;�~q%�E�#P0�*�HL&�i�n�z)���!��!ΟI>�������J�z7�T�4]$���)f7���Oϱ�i��i΃��\���[Xk�������`J0#�.�i�ͧc���@)�h�٧��F:~d,�;{�,������V�����'c����9�%Cys	0��n��n��&GG��Q��68[L�
wGm����a-���..F�j�	Wz��_��_J?�S_��U_��(�]�Z`F�u�ڿ�J���7�xS��X�k�΍��y��lE�;����J�;��$>���i��qT3�W� ٳ�etQ��.�a�	5|1���T9� c9ƌ��ٿ�"ĉ>�w5����h�ǐ�TR&�TW.�72m�W�� �󼭣~E��'�׹�`�f毄pun�0%Q2W��p5���j_f��Pu�uJ�~�Y��6��[e��.&	��<)%*�H��Ȃoa���	�3\�y�Zv8�H����]īG[��o�9����3܄DUʤ����|a��4�Z�Y�_  @ IDAT'�:��Z�����3B�H�N:�g&Q��Uf"-�N��ߜQ�6~RN����3�Y����:,/�I���i^��D�3sg�4�:E�U�����S��N\�t^�'c%���.l9-�����<���P$~�֭[a��'�x��ٳ�;��Km�*Z������0�@���z�7~�7FAX_A5p�3W�U��>�^��wHwD> E+c E��#�#BE,��5�"J�#+f�h�
�	�a�y��i�ft�a�wC:VK�b�Q���Ȱ��V\�S�%�,��l�JMd��3,�ԕF��k�%UH*�����`��2B�`Z$fU/4����
�o4!&K��!�A�=Lj�7+%[!�@q)�LY7�l�	�D9z'Hyd�'8���&�r߾r�X�A��[C�K�H_:��܁�(PSgk�.��"!���������F�����d�萈g��6�XH�4�M��r�UWL,jw�S�]w��J�
���Ey#��4Y�r�믽�րi��N���!����H�wt���ZI��+���f\�H��BOQ��v����A̭��!��ۈ��bj|(�?�8q�D>2�a��b&Ek�eG?0��W#�,.�ۘPW�srl4EJՃ�IJ�P��D�'���\,� ��XH*��'����O}C��wa�����g��"]:����V1lr���C��{�,m��Lj~q�Ǳ�e�޳�%·/�-MZLc�ddx�yFO2�B�p���Ąf�UY
��!,IV}�5Ҝ�FwnZ�̆;��q�T�Y��j~�Ň�yW�Q0��'n��j叇~��;�niwǚ���
(c�4��b��<T�ג��� ��Ƽ}(/j�׏*m�&���/N9����~�"��8�PU�P��bY�~���A��y�.�����A�o���|���\��>˫�h[�sz7��;�DF���a'쑿0�����q~�&Bf��56��E]꼢�k��o���v���i�Oı���p9~2|��o\���E]��8�3��ZKж�a�cҲ�t��:��x���0�Y!s/wa��}���˦ӳ���k�@��-�i�6s�t�K�0��>��wЃu��-�[#P�dg�B�!Rc9�;���@��g���������D���*�o�ElFx�>"?��@A.�o�ƕ ��L0K�+b�D���2	�oK�&3fƍK$Uϳ<��f��|��8[ �0���0��i�`�2����� j,�!��@<"7�l���z�%�����89;�6UH
�ź�n�5�v3-o`^iV7��$R��Ǡ\;���j�v�
�����`O:vt�e j��-RES^i����>�l��������m���������!D</�U��y�8���v�E��侮�mڍ�V��.���Q�&��ݹ�na~}Ǳ����8(�6v��>T;ON��1��� ���\_���Y<X)waܺ{S���_^[FbV��G�ΟMgOO���uip|$;q��j���ŝ����*��{�\�̅Z��ڝ�*,@�no��##q~	
\�V�
t �fU�퍵rwc�؇���g�x���O|�}���o_N���s���t/��;�ʷ�8��V�K9,7��9�N�>���ē���*1�>���F�v�D�5���t�ϛ׮C�u��jrs�B:�#Ϸ�!���i�6}�
���1��%c�q���t����QLX�o0~n|@����I�D�s�Q!c�P
�������8�;��c�M �Yb^c��0�UH�C�����\#괖���e�`�TsԺ��kMk��t���^��ɽ���������.;�q9��}�0�WZ#�~�����kb��� o���4���]�V��/��-��=Í������g��伍s(�V�y���D=�Q���>��q�<3|�7(�`׿8���_8�K�U�g8|�g�|ۆ���k�n�L���c��mMϒ���f�u��><����،�q�#�.�'v%�]��J�>g�n^�x�a�~��WQ�oY��~�[����@���R�����t��>H�%�U�>�9�	:K�`��DB��s�Z,�)��a"���"&����*�b(��ܫ�:a��K&��Ƀ2T5D��UD(��dH"�k��`�dp�I�G��'�qZ�j!�O����;�[?\z���@����������"�`�d�r�eX�S?�`�����=��t@��3��:Z_�PZ�]!�
�@����LtC��BlJr��!��	Tº�\(���A�x:�N�{!�NN�y�g��]T �S7y�a�}ll
��0T�j��M�Dm+{Tb�߶+.(	�%Ef���C��f�� b�S7q�
vc�� }�KH�v�4<0c��䑶�3K�#0(�����	͑�1���K�H��:�ˮ�ܗc���Գ����Y�+z:�k f�Y���^.mm�����Ň�G�}$��j�M�T憸����Sŉ�鴵�]\����O�ԍ����4��*'ߙ�]�noDߎL��V8V���X���#e�,vָdtc/��Ponm��=�H��c�J��8q�d�(~�ϟ���Ow��*�L���B	�}����.\C�0iǈ�͈��,�� ��l�\W�\����D�q�z*��W��"H�C祛��cKC)n���������BѺ[�oI��T�o+�?����Ȩ��Y�o��L4G�zG�<n�<L��p)4ӏt�yQ���pR(-v�q�J���cY-&�y�Q1���[�c��ru�z��
��J�+K<��'ֈH\3Q�w��V=�'o�2�y� �Bg���sI/���E�n<�VZa���P]�Z����VY��[��'}�m�!����ɡrbA0������i|��U~�w=����' "�Wj�&6�!w�G�_�7֗�\�T8¶�	8���,���49�庮�ƻ�b�s��m�5�0�dV��m�d�v�o4��S`r�����_ˀ���6`a��]��-�j�6s�t�K�D��{==]���ֻ��8�����|t���b���-�b���0��>�l!z	%�R�6~E,U����[Z zӊ e�2�¬t��6�S'2�9��N��-�H������)��_fHd-#Dy�X�\�V�@�+��I�����.+�]�8�/|"w�+��~�1���>p��[r�	���,�����xcN��ĕ���(�!X"`��X��H���rB;��a5�;���Lpv����3{�x������n�=~*�\t�-,^^���P孖�E�Y/a����J�4�l���h뱄x/z��9��[r���>HC0m=���A��ͿpS}0[H�8/�/�!�/ݛƱp7F[-������`��˕ݝ���lq0ԓ��o�����i�.E��T���9�b���8{�B��?��ɋ����1L6|(�=�11��ɷ4�����J��\�su���4�by�n�܃	Ez2��X��B�e�V#��ff�,v!����xya	���l�H�H�ʏ=�x�Ѓ0>�/���t�ƍ��������ӧy�$.M܁���KS�S� N�xҰ�������r舎q��|T�����o���Χ�￘�?	@���2B�9��9'�b ��a���ɰ wi�I���9���'ߞ�Rm�
4�#b|!#v�Dյ,�L�ZD�c(�h���˟U�չ.漒�r.s/��I�W�����"��w�OV���O�#~!�w¬o���C���7`���Ύ�]nNӊ����Gg��>�k�_��O��fZ��6���[��ͣ{W�č5LϪ}���,�2s{�t�����a�qL#�G<~˴����MC�V��&�&s����2xb������p;������:�Zl~��.�Y��}���*�Z�t�|�1T�+�|2q�k:*��s�ν�����.��XEK���[���h3W?@��ΐ.]���LZ�xܯ3a��ݻ�;�w!�:�d� ٖfI��B�$�Ͳ�$"��C���#Z��I���8�A��O��4��.���� d^��=�!!H|�5ְC�~�Ҩ)xT(#�c7��_�FiJ[XP������h�W�p�R&8[7���jj�7:6���?��٠����N��[���b-�v
�9.�k�]U(����2p2r"�R����L��8wݦj ��^�xU(���w���{�CF形	���
�t�vUE���ƎLCG���F����+������$f��&F����Ma��.-٥`��-&`Dd`��׍E�^,v���Ø:��F74�˾Y�P�V�d�$��`�6 ����9U6{PcD�đ2��!V�G�h/f��G��������ĝ]�i�zla�.�q�L:8�`��L��z��b3=�v-���b:}�g�T|�ӟ��޴���}9��<ޘH##���Aqsc%�7�҅����i�̝d��K��Oo�x��4���Sܱ�����\@|sm!��ZN7������wm���vJΖ5�R�pw��Ť��t�ܩ484���:෾�'��"VGFˋ�+Ν;I�#i[�AquD����	�d�t�N���#�ؑ�H${�6ck�g�����ZZ�XN�<p_z�я�	$q�P+:{�.�,�mU]eMb�b�	��S��#��к"�����,\5Șaq.#�ѿ���j�� ~��i������ځ�~�g��V�:���a��A��3v2a�ymPb-��4��O�aX�0R�g�%��	5��H�e!��7L㸋3r<��x���䎩��������Vހ�G~H߾qf򮰚�Л�2�G&��w�1���5 �#��oy�a�۸�u���#�??��eXf.���߷��D�c`�,�ƍ�8iШ�m7N۶m4�m�ܱm��ٱ�w���s����y�<3kf�d�OCǨɤ�NO�o�ū병
�:�����u�:l�������	g�n��&�SU���Eu�ȯ��W'��V��s�բcɷx�<����e��t�x�W��|h�%_~=��<$`��]LH��7 ���u��O|�	
�Qw�s����7Y�Gg{[X��^��3dD�*V#j1c`f&֟I��]Ȉ��D'w"�Am=��Wk)12G�9��K&r�}�=Q
ߠ䛤��(2c�BIbw��?��o�/�)v�ƣw��e����8K�X�5�l$9bE�(\	�����By3׫?Զ�}N���l�2�8�98TbS8e#����m�CsM�P������t��u�����/�����XOm��� �V|��q�c���9)��ٱbq�����Q��)%��c�����mڴ[�8�Aڧ����o��YA+[XqD�?7�)�Ka��SE���;���#���<FQ�ߙ�b}MŇ�SkŔ��)��ɩ0Z���Q[*2D@�M"��u��t����OvsOë�"T�Z7�bI�.$+���a �w�������#���J��ݜJl61�"�G���{wE�22�bHi�찴�T�P<ɉo��өΑ���O>���b+:1�/�ϱ�*���5v�F�8���o��2��lP.!A�땪_� ^�u@� 0ރd�l���<i�lu�pd�T;U�l�j��B+}'�N`�A%���/u6�"F�qo\Y����m�{(�U�<o���~��C����_���`��|�b�Ռ�o��"��q�;c��_��s�6M����?1I���ew�t�&�5aBt�4�EP?�=�٫v�a�?`�?�e3#�t���z��SA$^q 7�Q�Q���T���\&c�?� L�?�S`�7��vB�	�,�P����Pzq�����/��ڳR��ݞ�T��&��ҽօ#������%���5!n�
5�3^:�ȡjcߋ��z���U���k]w4v���6U|���r�������)���?j�9uՈ�>�l]���'���N�cl������H�Gn\'�����TB��F��,Ӳ��5u��I	���� 1,����گ?��Ԗ�����#�"2@�k��[eɢ�f��>�m�8k>k���311qQ�
�&b���!g4E����)��EƱ�*N��2�P��#XҊb�d�*r��ꌷ��35jc���P���2(dc��(�eV�j���{� �;;[����L
��'3-Z��בB�a�%~���b�nM�IE=�J��R?�+���q��E����^�@�������a��$��E`���� ����dD�`�]U���b�#!$U���Zu;\.���� �m12p��?2����_X����/�_/ޔ�E��C���ݶ��E�i�M��IoVڮ�����%V�����8���{���s-O8Z�I�2`k���/e_���pE�6�7�[�KA��������},с��@z����d������,�;��| ��ʪ��<�P>н�F��~Sk�y��z]�F�*f�֞�������l�~gL���O�x�%��`�6ü��c���i2�t�]C�����o�1�U	&2��K�;���4t�!;��%<��x�&�OcFT���esOS?���c]7W8`��/7qVh�.��i������_<���\���e�OEK����.��2��FgZڛ���`�Y�:<��x���pX�MPx����		{!���٧�(M,�vB�
`U_��jLG&w.��Y������2��"�I���WMd��u��(���zE�(�BAҀ�m�]e�cA 	���͆cCR�ˍ�����}=�cSPb]�(��t�������)-���:�����\S|=�9g�Ff����C��צּ��/��V��/[l��[���#�Q_�t�G�.H������+�UW��`�-�/?pĝ;�1�iq�-���s��Z�3�>I�.�W`���಑V|������3���ZqId�m �e�2)�+����a����qn�����p���4fY�̄�8���L���>ƵTy&=������V{�K�f)$�\�������������T�L���,F��a?�_��W0��ԅD��A�8� ���ow3m�[{}�n$�FZ�������1�&9S��|���;ӱ"o,�_��";���ÿ�ĳh�ٗ��y#�:qU����@��x���Ѝ��e�G;�g�i䱠�z��׀	V�M3�z+s旅0��R����8�mi��D2��O��QVU�=�/�����/�=F�/ԣ�����,�#�Uղg�N���tRFx���(t�S:���F.�'����)��|���h�P��P
;ԥMp�66�=��w��}f�B�U�xG\�K�=���"�\k���V��u�qzO_\l)��nk����<�������j�t����ҕ�eO\���.|X���P'�՚����6][em�����d6���K���`�h��
M�G�^ɗ}�6�/nCn�mFuf���w*Y��o�CG�����2W%�y�Hj
L� �����s+��\�q�����Hg�Z9�.oB���.�c�5X��W&�[^��!�t˥vo��}y�����_|����q���q����/m���4Jye�kO�#�Ex��/v)��f�$:1S7��s��yn����%/��:3��.����U�8��d�e��2�cQμf̈�c5V��9�-�Ͳ�	I��<�V�_��A܉�^Z,�wF�pnD��!�����ƃ��e�%t"E�0i���(�Oo�-��3&�N�Ϩs�ϯ�=񈷜mzp��r*K�t߱�9/��ګ*&��H��8� &��l�8{�Ϥ''.P��Yj[�s�mwL��3��<Z�#v �^gU7˓��A̋H���{)�G�n�j�������j��V����2�VK#��o,f/��/'h�}�H?􎧀���'��em>���۳j;<�n4%�!��a�F?^R�S��o��x%���!���H�!U�P��4O4/
����U��Փ�ВI�G΋�[���`-A2&A���],ʺ,!}q�峻#�-&Q"�U��h�;�L��,�����/ �`�dc�{�/��tCG�4���V�/�ZR��R���Q]�6e? X���Y��G�)?�����L�ݝN����u�e�3���S�h���f�c��J%��/Y�$���bѸ�N��� �������ػx��tl����\�я|�mq��P/Ưl��P����-{Qa�����/3�2}�P�5�xu*،�[�$��p��S�(TK�A����u��Φ>�'2A����,.�l���tM�C��]C%�#��ba3�;�|[[�8�՟��ŭ�X�9=E�� y%/�3� �bt��ʺ?w6-V��Y\t��x��M�gGmM�\��H�r�FF�t�]�:�v7F�X���Fiz_ż��W� .����7w�X�^��zP�bYl�П_l4�7?�9��-�}ؑB71��~�V�zX75��X ����}��*����=�1x��1?���ЯO�Fɏ�M�K��8�E���6�3k����nIw�VsV/��p�DP��ʱ y��T��A>�BH�/�O��%���(�ɜ��Q�����ɏ�e�R��8.`���.�:p0i;k�"��W�,>���df��֬b��~QQe���1���sv�uk���NX�Uʌm�V�ײҙ�?�i�%P-�u;�z>����ք)�號oGk�~�Zo�4J)ڥ��t?u���˫�:fwٴj��qb�t+4:NC��?��f����x��*�&9��=ד�ֵ�
��K������oV�`T�����}�?8ʵ�0����Bw'˟�:�S���Lv�SP+���֐fh'�0'�?\�Ԙ���>�nXQ�l쌑���[㚙����������W9�4�-И��F��Q���X�7,9I!j�)8�t�[����O����0��ѝ��#� �L�*NGA��� r�Bqu¥~���d�0��ʈ8���$��7Ӣ�:R*Ԅ����$�V[b�W��ȷj4KH�f��1���]�����?~S(w��be#7�������A�w�I�}Ơ�j�H���`Ӯ�S>)�/�mґY֙�	��]�V�MR� |�ӱui�Ũ%�^C���S�S��I�Z�!�_��|���O�7(e_^�9":q�`�,�'�khη�|�[K�A��/��n谮�z]�+�K�T�����:�E��LI7=���}Ax}l��n�nM�X�̛~�,��k�j���HLef�ȱ�C��@<fTX&�K�c��'��_TXN�.V�]ڶ �� �{R"�_x׀q=��Z���̞�5Sced���?VpXRNVV�g�l�9�|~��L�f�-�>ώڣ>_�|�7\�^�2
/��~̌̌%?���d?:} ��(�
�$���������
@|��OX&���AG�?��[
�ڊ�SX�c������~f��\W��p�m�L��(�mXH�bB9��D����e��5�u�hz�T�r��g����'���G�%;�?gY�L�
�BE�#��� [mb��B瞪"N���e-x#r
�������!��vx^�M���Đ�;Ԛ�;���$� ��=�D���f�>,<���5�Ì�|�O>���2�:�N���"��	M�{]>-�v*��{�|'�~E|&�U�p����� /5�I��2�,��6�$�`�m�Ѡ^O����s/4<:=-���o�{��~E���T4"ևan"l�����J�_]�
�@��
ZD
��Ę��x�L������2n2Y�b�$O֛v���ܚU���Y�L��Y�
��TB�-�����ϟ��B(��V$������`,!Q���eD6�V^�x�Ω�-��,D���D�B*����
�ReQ!���<D�R]7��1H���4��K�>Xq���R��F]a<��Y`�\���1(
z%�hwrK3���l��R&�Z��ً�.��X��_��CR����E�iA1������p#�2�򩽫��ՙ-P+^>3�z��2�����a<B�nH,F�Gy8�)��B6֕`4?���L�a�4�0B�ڙ��B������I�������}X"�GDm��W���U�A��9��m�d5{�fY:d�Q#�ÓOC��݃"�Hg#˾��~d�®���>� ��K��P���©T3�7�)��`���R���=>jim��f! �ҵ��Eq.S�ux&;Y��k:Y��ubE��)c0ա�^`��x��l�q�v�˳o[�M�q¥������@�Y�����tq�h�hx�2�,ҟ3鬒�?cJ[=��>gj.�DiRt'���{��"@��p��fq��J����6~��]�ܜ���E����9���X(�8X#�M��8��A�i�k��M#6���!ڔ��]V����b-�1/I�!��kh�,�c�ܼ[�ʸ��W]A,ǝ䱨=1?q�ʤ��=���t�kBG>�N��㲒_Ф7q]���O��{*"h���KSw�*�q��;�j$���q�D{�:u���j�۵��u�!�^��?�u	�x�h?k��/�Z�lS+���;��� �����r}Mw�ot�`�:����P0q��6W���=kYzkT��9Pn^E�â/UoE��r�;�[���/���M-�������|�j��b����ϟ? �k��@ɫ���5{I���-��<â�7�y�4�Y"DO�5؁qB���e��i8$�I�8�+<mv�g�D'C�>C�����GV Q×@���ij*'ڸD���}���?��0�M.H�6 ��4�;.�E����a#��E��zд���B��$#�%�t��HC ���&��B+���xn7��\���ֆ�F��s��p�����n9��Q�\�A�wGT���c*)�e&�:���ZFǀ�4 ������c�������7ҭ�@s���n��T�󢻩�#���U��Eo�JH>��H=9���O�U�N���
���9�s[���������������6
b��(oQ{��fN p�o�tL\>&W�=͛���\j4
Ūf����Ҙ���/b�����F~����\�|���Y�M�NG��UI��F���1�������+,��Tc'*�N���wrVF��&�=��s�9՛D$2:!�O���
�˙�����J�����h�?-O��}���W�:;�f5k��L���w8�qq���B��kjk�c�6Lz��ݹ�젙)��� ��������=L,��V�-�E4��7r�>��Nw�	����v��$6�-���d�}ُ���aq��J-C3.۹�̘5Yp(�x�t:wڠ��uԎ:�Ԝ�2��}����L��`)�8�(�&��Ai��|��b �5��?ԏ�ٲ��L�&�J�Q���O��os�	����`WI��8���Ц�n�Z�I8��^'<����|=��N��-pO�S%�L}�=��fiD{m:+���-e.��M�vZ����up�Nv��׸�n��7��s�`�����ޑf���̏ ���C�5`	��I�r���U��D�W�}ⵦ���
O�Lm���7��HPc���jg<�Q����u@�ˡ�^Q�`������F�0ů�[,�#"�8'��ed��o(Y�F��$��r��1��\�D"�>4�h)�O^LQY������Ƞ$r�,7gHX$�����fck..�B��X
fQ }�j�'ї����Y!�K�YJ���|���d,�Yғ�y�yZ��a)3�o��Z��1����7���MJ}�d�Q&z7D5��;��U���!�	�	��v�������X��P���pK�>�����d��UD����y�PP�J����ҍ0��-km�������Pl��[��d�Uķ�X��t�mcX'TP�����%�3�W�2��A'X�}�r�mI[v\���/Nm�g����K���'�ɽ(O�����rz���;�
K�&ԅp�����w��s��̞��ztP6���}H��ǒ>b��2��3���!VE��^,���OkG���$���W��6r���o(ꅬ�QU*��5�[��?� z0���Z������%�A.��.�D�dE$�ی��oU6�� ��c�S�����ǅ���]�3X����X��+��a�  ��2�}����n#�#H��Nnam��(�T��^=����l�,�G��lց�e,;W�j8��?�\lH�iR<�S&��J������M��˟�&,� U|��fQt0��j�6��ö�N�寖q@�z��U���\�N-�&��*e�{�h"<�=��,������v �"_��؇�E�Zn�����]l۸S�C/�$��n�o���=���f���.X�Bwwt	��1�(�M�#&y�<`�vk����<i�[�nIuLʿ=�7��R��e绵.m��FR0+��H�9z�I�:r��%�L�ۗ��O:�:�+�ㆨ�cB��<IhV�F=A�y���J/���P���ҤߔjVΰ<�GW�5�[R�'�2 s���@3A��_t��
mw|F�1Ĭ�Ey�0��|¸<ו��.��W�� �nך9�'p;��  �i�A>��Eif+L����|�-����J&:�QG�K���p,��T�HL���:�s?zB?TsaW�"�W��������*-�Ųǅ��*k,�`'G�@vD��
m �˦<K	����ZmC2�H�H�M�͉,#u!��^��D�ow���<1d���ݬ9B�S�����\�����Ћƀ�b|��2�XG�~�6��������tz�J}1���\�.��N����r9�T>����X�������]�5͂|�Q�=(��J�6�<%�?�މtf�(ie�z���+3�Fј1��Q�v���Ϗ�W�\�/���\�o���5��2$��y;�7�;3]ݼ�f�ʎi-b��GW�G��v���^��-*,J�b���=8<�����1`~NO�Zk�6��}�L4_�]����b�Zmֲe�����&m��cz'E�W߇T�u{X,V��&������w�A�� -ppp��wu�`F_<�M<˻4�4�x\�f}ϯ%�\�X2.�@�7����h����JN�&��T����ʹ���X눳�`̃�U���V������pOGS;�l��ϵ�銋C'�)RǾT[o'3�ڎB	f�/�ЛO��5���[�\��u�N�Zd	V@�f��|���.�����y��u?b�������͖~%���/��c�z�(S{���e#�_������N<�-��4UC��F�:�����6Cr���hW�Ϗ-�\��}&��8����y������;�֐�DQ3�(���MUI�TlŪ��f�"�}+�=���	H����AK����X�N���>�2��="b���BtD4����ߣI�D����Q�Y���l�amF^��6m�Z89�h��������S,�����+��	i��r3*�jy���Iix
0�]j�<x�)O�1�!�I��/d5(��W��3��r��<�r���y�'
�R}��),L��)G��ՕA�T���~���KUt�N�H��R�X���T:(P�ѫ)l?���0����Oc=:��������@��6�yU���p�	��!Y��cg�M���;W�1&|2
�{~J��(8��{U{eh�����n~Bl���9H�����Q�
g��S;Q���U?�ã����H��������V�H֐��s	@�w��m�5�����,��+W9��T����k1Av
��e������w����H.Z���24V>u��pa�munw2{�����P�9a#�Ȁ7�\5|����7�׀
s���|��i�s�xS��$(�5�p���	������-$H�Yv�:��33�4BYB���i`q�X��/f��T<f��� �ו=�"�(�Ǧ�v)P�}֘��3���Vi��H���!9#�Za�΀9r�Lȭ�S�T�B�'����'���\j��r%���j�����ČRmX����=}��H��7T��$��$�)�d����������G��:5��V�r��D���??IQ
�,�U�U`6`	�J�d[��J���J���0k��?��*�����?��$m���m����,5�Q�����`�s̠�J��&��U�ˠO}p���j�K��ͤ�k�V<`�[�&�:��F��+\|#�����0i;���1�#�؎�P�D�]��j��I���>(��$k<��F��e�?���R�@GGE9����pt]:����h�Β�F�+|����V�\�r|2u@��lo8�f�ɩ�c���<C���n;H��~��Ȯ�/�8AP����N��9�~�E	3�����?*ZE$c!+o�o�]��_UZV�\���v���yP�K�uG%K&���R&���H��aZ����[H��R���Jwe 
/a�r�xZR&X��9?���0���(�L"�r��^I�?�>L���L{���*�s��W�DE�T�z&��3��Ef#`~N�d�ľ/��^�s�(�`��b�n��juĔ���+��e]��	 Nd����k��K�P;��fO��(�y)�M'�=y��!$*6W�lD�Ni+�͌J�/䇕;7����|��&n!8-���ч��G���S���w1t0��ߛ�~����#K(d�E�\�,3��T�з�i��b�!�2���_�yKw�~\2U��x���~�������|K�Њ]OҠ�Lv+���6t��C�Nyދ4�$�;˥��c4��3�a��Ɣ�5�H�}C�8��r����(I��QE������c`��tn�G �0���_@[9[��R�-U6�,՞_dhrƘ!LM��Z��Qmw;4�[��
�x��9���M���M��W��������j�.o�-���/I�ޖ��hw�	=��J�?F�W"�;˵�o�Ju�is���C��ʕ��f���vۨ��	$�T@*ߗ���H�m�m�.��������#��=��c�4��4������>�����}�n��)�XS�#�VW `�ž�wMx�OB�����M��Xn1������G�����Ex��k-�b1ҫX��7��]��V��[i�/�;n�E�5���V ~q�IW,{c�U�����@��t��\L?��oT�M�t}Ϟ�c�3Ý4��� �i�nx[,�ܪ܎u��w9
����e'��c�`����~�� �>$�&f�u��<��<�ϩ�o}��r��v�!"P�8HCcw�4��0�c�XU����R:�!T�A�1lJT�n�0կ�[�b)���N�6~`�=����[H���	Т�8|�P�s���T��u�E~���}���
O�c�8�h7�2"h���Ќ�:?�Y��K����Y ���NMt�l4�w�Ȏ����?�x1�B��m�,Y��B5$EB��Tx0��г��}��vi��M�4�e�gP�3Ze�n���G�.�|�F#]�L5Y��A�yw���kN�B�{����&������vE:�X6\��~���&N��8m��
Q<��s�ȵm5�%c�m����
�]+\%����6�S�4�������6����!�zͻ��z�o;�S�W"�S߇���=���z����v�ïx������:$�oq�iƫk��w���	�.���Ǥ�2�ƿ4u�4M��W�a��khQ���s6���ķ�th�i��s4�c�O;�ڕxU�+=��f��rҾW�Y�]9��ϫG�
�G�@���*#���۝�f�>�X�}y6��a���Ь�Z�b�8�a����G����S�Oy�ϗW
�h,�=gTkwt�D5[z�E�X9�y�J��a�tؖ%��9|C��_��C#dON���x�6�8�T�������b	��6^�E��Bɟ�$7ۄw�u1{Wbg�cL�|"r�
�̃[v��a��Ls��W}������w��-��1���7+3�����~��o���:�-!
��3�\x�}Վ4w� �������izD���E��B�������ph]�SK����PR �g��6��P��ku�',�����}n:���d���� ӌ���{�I��)�]�>�ْ��{��K�t�oy��{+��=Fm��`�}�p�u7���+��|7�|�L�1�%����y�{��s��0��UZ&/���I������F��W+~������[��{��2��S���������{�ұ�V����?�y��.�{+��Oj��nf���TP#$ҹ�U�D��������}�yz�2K�vea5{g(M�u�7��<�����!��������%1*ؔ�%z��N`ߘk�CJ��g���O����<dD��aܵ�i3�!r��Ŋəj~�c(��pO!��Ya�>�|�i���B#����&ju��!P~VIh���A�܋���
�	OMk�TA�K����!WGlGw�Q�]]g\�ύ��%�4��6~������4Z!=�����d��U�iG�RfΓ?aA�ԛ�+x��Ӂ?�v��)3�F:���/�o��Fu����ܖ/�]"|�Ў���� �)��.��c��C7��T��3Ny���=m�Z��+�;�K�>O pL�ܚ�R�2AGkZYOD�K����+��*�}�$�p#�4J���F��������Vr&El�B���VW�˭�&� �o���Zח��\5������b�xbE6ݶ���L�f����<p����5Tا%(M�=9�z$,���l����2���huQ�����wp;�y_�!�c �|�̹^�DLq��Ҙ��6/��y���n�P<p'aǿ�/9S�LÉcS���y�Ƥ;�[4N�,�A,%�%ܴwqq�$�ү]�� M]B`�v.|�w<��7g��|�@�-Qd�w�C��&�����ڽa_]�v�zUi�����*]!jXS.�[Tl�r� D��9�Q3qq��L����" �1�2�!�{�.?L����dv�ǆ���S�Q��:pݧ	Eo�K����e���||�N}�� c��U��4���Ė�Љ�]\��q�VsL�0�$�ڷ]v����&��>/��F"dS���[F�+t�B�a�z��L��|Z!M�����f���r!���I��f�s���TP�$�ej���9�1��-I�9��
�P���#t4V�)�Me 3\�@�*�2{���|wf���WLt$-�)�j�PW_��)|9E^H(bVH+�c�Io�������F���bh���t���ڦ�t�5�h��#��*������p�jmJ��A+�\����S.���;T���Kd~�ݗzs�az5������)���$=�M��n�5Z�C.��%S�����w���Z�W��S)��8��(���`�bn�
�<zq-Ԯ�I�/iƇkR�����[���'�V%�S����Q�ӞJ�R��R��lS��r\���+:��(�|�1��c���鑣I:ݝgWR�8A��<~��&'�Ѡ�?<����X�����%�ϻ�|���|���pF��X��S��N�
r�D߇����lSOO�fv���2A~���*/�ʾ΍KWi�%D1���v��xKV�=;��^m��\��]�'S�=�!3�t&�:���.O�3�:�,zӇ��/w"���6��?�K8V~:����)��f[6:G���]횷�2W���f%�S2�Q!ݟ��&�}��Q�i��j�
^���Z�����[��2����!�Z���?����(H��l�Ŗ�H����P�1��q���Γ�����bZ{�!��j����f}��R��9[zh��#c����'�0|���kK�ͣ�� �ヺ��pz��R[�{~���uߢFι�8fa���<M��/��B�-�-<:0�x���}��v?�f|d�`e���s�OK���?���A���	����n�λ�$(��t��~��ʗ���k�EW��qz`4�?�W�����[@�CR;&+�!�Tdo6�"���G�Eޫ����TR�Vs�I�_�j���}t��"5�����e^�� ��̰�wfaX����M�c����O��(!�p�.#J���_-��?S+��#��(�5�>D���{(�s�،$p��_������g�D��I��嫴 V teT2K��`v��@�w�q�H!�����d��aF��L7���9��U8E��U���PC��A�3e����D��7�a��QD9_������Fj�D�}q(�����-����y��g�m\W��l��k�D(���]���{pq��3պ���������W�:�t��X,���.Аo=a�a����76�Z"�Z��3��G|e4G��Ja��B̖!��2G�Ǩ��w�e'βl���,�*��L�?�7F�hw��u0os�)=Oۨel�jͦV�)C#��1���ju�m�[��;*��-P���5W��/y����@>�2���-v���_�Q�-\nˋ7��o{unB�%���{=��f�]���2��ϖ����G���Fx���d�6ZL̹!��)!n�$9��}lh�R�p�Z��6� �-��k�M���č���3����W����%�@a֟��1�6� ���I!�|��&;�����r!�Seb���zNV���qt�ZMx :@p245���@���JM���S�u��]EA�c���7��5����os�!eʛB��8�F�~ZZd�� %���N��q�8`6˯.���=�ݔ^��9�l{RůBK�ќ��l$^wClIؔ*?�T_��r�z��9������:���L�^K:}������6q����Y����@/�U�pjZ�[k���һ��~@�߫=�x��j�WX���r5����)p�=*�߭V0�P�fBnw��%2	�(WP�[�9�cz%:�Dz�)��>;���$2D�h�/��\
��~+Y~���V*�ήs�yQ��9�Tjӌ��7��#��ET�<d���0�P?A�8� A��ZZT��=�/�^��]�b�O��2�V	F(��	�W:8�V<I���N�ͫ
-���[%�UF~��L!�Pq��-⚠��1w��q���[g��ٞa�����@��b��t�[�M�^�4��lP����R(�nҐ6�d�x�9)��b�1�z�����Vl�����ŭuEW0!L_/
4Y�cz-�����fc���❈��e��_��-ʵ;f��ZJBѶv�]@����r�&sXt;���+3��Z��7�f�i[�kd�8��-�f��%�E��k���T<#�Ye����0�/]vD�#c��Z�9���Zn,�Yh�������GN����Ka�`�fTt��>C+{�@�դeo�lߊyj8Wg����.}���̟c�9?rT�r~���O�=��[�V��Fyf�G�t�"Z{��ۧ������ ��Ĉ�8��ȡ�U;�|��� B|��������2%��L����ٴܭm�zWǹx*�燧�_oA$���I��}~V�>m�
 $���5����t��Yڨ��6��X�j#�`:wVE���H��ڭ<�]6��?���k��G������=�$.�Ƈo� 8��%t+LBH�X �?nu���/�G�T��81>��q�)����c������EIT�/��p(��n�[��s���v���/�2�xPl;��������ݚv�i^�,Wz���[<���TY����e�Ǚv�9���)( ]���f�[C̝a��u��J 1��ҙd^S����1��'	e_W�1]Q[�˼H߼��G$�I'����^r�>܊��_�p�a���?n(DdC��C��A;=�d�p��3���)n^�m�j�1'�8d(��\e���G�b!�'������N�|�;������`�J��$����?.��v�[� c]����-G�����R?�V4'={W�T��%�ńV.Y:�c���0��0̯��dXgXHs�N[K!E�M=6�EÙ�4�lP�g],���bH�4B�5oj����ΨL�K4��$e���Ɏ<�$�"����;`~��ykoX�k��^��\���� tO��x��?�� �:k{D#�j�)4xnx��󟑡6�a B��\2�ue��P��oF�N¬~5E����~}���o.��+�b����}�G��I���X@�l߇x�PǤ�]�z>�$<�^j��ٖB]~�i6&���<��$�����ngh�OO�*6�F�8L���$�S$��W4:�yp4|�Os�x���Ǩ��Z�4zb�A�P�C��95zM�6ř��8�ss/�ܣ�E�7�8�㥽��Ý���k�O���R��?cJ�k3-���u�@Y�.a������E�fۘ>Փf-�sm�?;�d;s�-��J�o�b��	�Q�!&\����^���SZ�{�Ð��L�xH�[;詖���7�{�����|���ap�ڡ6����s�*�.h��:����)KK�/����r��$�ѯ�s�@�������`mo�hF��],6��s�|��U��R�iU~��7m��-
n��BP�ZVɃ��*!�}����+T�}�UMU�ӕ:D'�e�پy�����;C�ҽ ����Z���!�;س:��%�O0�����P�g�ʴ���):�������c6��UO� v��.�My�	���|�oj��� 5��dS����a�:/3GJV����������G���(:��r��=�ڊ-ǜ�e^�v��~�&��~����M��0$7O\&�D:�6uNqr�T�_�i]R�^c�	^�Sl��N7��篚�L&u���3G�c��28��z�5���>J�=�3MǧɖA����I�,��x����Z��+����o��)�4\�Xm�3C��`��o��.��0�Z�e�#�K��R�<�ԗt7#�(>4��;0Y�cx�f;��e{��=�	��GRbG�|�Tϣ1��D�Pg�T[$�h
 ���3�LL1���;h�~�� p(s��L����-���=6��	6���{�a����x�(���[��N�S�S@���n�N%����.阡�!�^���>��\?\Ǳν�Ϲ�^rn�($�o�F�F��g2(����Y��\�;���X����$s�^.k�i�٘�����J��7_�F�ߢ�
(��% E�ȥ,�J3�Uv���-f7������q�qj*~ф�'Ě��m*b���(Ÿ��ۨd��P��nN��h�~�܄�jF��MӉI�p�vX#� MX܏E>�p{ uW����p�m|It��~�`u�>�����2X��S�
�>l1�:�bk�9B�l�_a���9�`}�KL��J��^p��n �ċ+]:o�+��� ��s��?=@P�h�D!�ާ��(��m{��n���|B�����5Z1�Y����~#D�6���/qE�7B~�@��b��H?gw�s��"����%ф%�F�B!�E�����#>�^��mg*��N����gx(������6�BE���u��F���,A/y�|O��8��K�}����0"�;���/_�G$�'̎�:�T(&��oR�[��I/3z Ċ}r�Kz	�:�J�D����]i,��&��I��)��C��~[j}�W�0ePʻ�Bg{�-O����σ���ِ�x�J8�,�L>�׻�53U�Q��-&R�\ѪW�]u9����{P���%[�����!�pn=�2O6��m�
�����(���p�~�G����b0�]��滉�9zs��f,�r�b����b�!��5�d�B��gh�KJ�jQ��4��פ���V��L�-Q�Q��a!`<�%Y���NO���'���M0�����u�����YsچT}9�8&�q�pF�IQ���#�k>���t�'�,�G`9�S$Q�v��oeH��{��������z�,����n�L��[Ԫ�1�_�S՟�%:���4_�B�*-��zo+�ꁟ�[�4i;C�^f��E���C/�6��m&�YT&ݝ'�?��\���9�#�|�=�M�W�q+[��n1��\�K.��
O��&��߾�f�����о�"C}7ϲ� Wu1�����`���u0_2n{\�����y�&WY��s��$XIkͧ�
W=NT1�0��\ @���!�AsrG��bѥd�jI_��U
��KζOW]�d�I=z�gi��V$ʦ��甛��ݛ?U�^.^�t�A�_aN�X�sʑ~}�9��d
MSgϟo�G��łB����xKG�j	ҕ�Z�D�=X+/���zC.��i�"�qױE���U�H�V�jok7��A�M29�]�+��{��q?w�6���Z�7��*t�������vpԕ�-��=
>�d~l��d<��8M����XmU��Q�{�B@8;��,7�h��2VAV�U3�!<0;���`/R�E'���AR�&�硤(�:�W?�_+�~[���)�&�-�<6J�����uW
QzW���V��u@��zܫ����}��bA�����iʮcJ)���3sv.�|���2,�ߺ���w��ބPF���L�tL��2� ��;�Bq�*X|M�۱8��!����X�s�Dj1�2�&���(��b�
u��xۅ�V���߬��lam����6>u;o~�[e"u�!���$�h���ԩ��"�O�'s���Xɫ��fMH�6�t�IĪ��(���jc#>=���֗�.fNH�����G�����#{'R.��P�=��߈���Q�87�9iN,�OJ!V7�_�����A��I�ω/x䪹��h�i������=[h��|��ܐ�+Й9�)_B��)CI���|J��|�I��ܟ�Z�@\yj	���i!F-[�ꮾ,��v��sM����u3�uy�6���I0����W����Ԣj����.Jk�D��*��s��1����H?�㰗�/��!��U-���<��+K��-Le�ͣ	�ǡzW~:��<��/$A�U$U&;��k�&�?z�˧�L�2[]��gJ:�4]����qe�<#��~os�L��u����<��Aqȁ��C��x͵'*�4AOz��j3�����k���	z�2Ң��S1@L*]�[|��x��H��`s��M&�F��Q���	��ᥜ'cȐ�{MfK��/ɯ3H���j�^s��K��3)�x\B納�Ǽ5 ���ly�-�����(5d1lL�%�I���y�3sw�T2H҂��w\L#��,�B�tkl�y]	+��B�'9��bn+=I���\�equw]�-���M���#������qn��w�I��M��Ԥ�>�'E��bD%g���b�g��2|.�R\�(�R;I��,��A�gs�XQA[�1K��k��G�=N�~�Q%W1��}���p6���l�� ��|��W���ڽ6�/�Aw���Z=@�d� �]U���o�1䧥��7,$����P�yxf�mֿ����Z��]Cw��!k�O��O����f ����;Y�#q����`V�0���;���4�t�:���j��9ism�^�)k3td�}�
_���\�O�����\v!�,�g �8KE�J��^������paN���0ͫ*�q��)�J���l<��E3}GӢJ���Z�I���ř"�NV����r�!�:$':ǣ<�T��-"S�҅>��o�9w1/g��y�i|��qS�[��檇yj����'?�I���Vb���/1���nI���!ka�|��֒�����@+��6�s^�C@4���'��V�k�W)>�s{�j�@��I��*G�E���ᛑ�q�҂��e� ��`E�e%���H�D)^�@�[�荆�ד�%�|,�AM���N����L9ƤL	җ,�>"���	f��LN{��py5)X�M{�i-�����u�C�l�t����a$�,���2�2 e����jw��$Itv�]��(����efE^ڷ�q
�XҍW��P�%�U�Oֲ��;��Wl�������5-~N�zL��|�[wH�p�Ӄs�_'�h'�% +`�K�L�x��:?�-*̸xlW�h�z�pTPZx爢)�u�nE�ZI�\�Y�I_���]+|D��,m����jQH��Ld{y�F	�����ε��g*�I�⅕ɏp��_�e��Ď����%$1;�w϶�9Jq#�XG�f���DYiN��cs����|�%ьg-� l�?cWG��ё�>%J��.��ÿ��M$O\��//�X�Mo���]o,�3hX�E��V�3��G޳�L3D0��. ����؉\�y��T�M�׻>�r�M����4D���Gb�O2������|�6��8�"o���&9�$���J��	��ڥɚ�h����LF��IIS�0����GD�<Y��+sB_t�c�h=�A�:VA�~3zn]P=���emԖ<zA�U����u�C��0�Ú�_��DC̷��Vt���z<� {�PC�~��BCE	��∤6op���g�g�2��h/>�fB�m0?�8���
e^����D����f�r�w=$�_�u4��m�*_��D̝���4�?�-l� G�}Q{	h� ��ZM���(�i���c��c����y#��f��Jm3�S�ɷl
S�D���s��M$�B}+������%��rݾ���MCf�#b�To��_A^�p��r�Oh�Y�x��}R�⭉ἢ�-��,sH�c���>p8�i]�@l	����ͳfs�p�70�
;�)9�9��d"��sqfho�Fӹ�/�)9��&*-�6?!V5��]����a�׹:`�˙��K=^�s�-���^B���{z��1�	�I�.��G}j���]�A��z���[Q�q¯d�f���ASi����=�Բ�D��*�VJ�Q8���ƽHh��+��񓑂�x���g÷W��x7�= i~P��,���=��֡�Qψ`�[[����$�$P��C5� |��.��t���}����8� �X*(O*]��e�hS���d<�q�֣0'�]o��Z�7��U2D�K�kpkϵ�2Vxj��,�m�D��Y��&F����?证�Q��˭Z����L^ҏ2�J���{�t��<�.��Z��Cr��N�h��#��U�$�[����'���A�%�$f�����P-C���:��'3�,G�����J��Zۆ|\��XԄ^a�Zk�C|�s���$�+�p$Ҧ�:U#'s%/��9'򏕡�':Rq������EN'���
fe�k�`�N���5��C�ɘlb�}k���ɕr�q�5�_wjN4Y�9W'>� O����܉n���@�R����#+a$
�Om3s��R��#��{o~��z�;w3��q��z��1AJ��9v�݃]�"O�C����:�OQ�P��J?t}/_z��]��}r�X*�����?����w-�p����M�Y�s9�t)��154�]�!_�jw6�l
qz�i��G������f���A6̶j]�J'K�<�j��4B�~�j�l�ʍb��G����쪴.Ø��	0[����TsF������Yv�5P�v��y��l(.u����%�@�Tv���Oh[�8�%�=�H�ާy�u�y:��Ҕ�t���V[\k�!:fO�z�4�(�acוNh���y����Y�ݖ=�SClh�e��5�Ø\U�Gx��'���G}Z�Yz3��v�8����)xt�D�0ҧp�C�u�tJ7p�q�����y�2�t�9�^�0I���9����Ivů�?M���c�<��I���d����XLm1Nj�$W0�<陊�hO��	SX4s��L���_Mr���w6;��|�����^��Eʍx��j�ؙ?S���SԽ����Ҩ����I�V,ط�{�d��Ojו��h|�n��F�c����7�N��oy�����,$�G�kY�o�B�����[��ب]�|��+I��mo�÷�����;z���OE��˵�#� $�G9?@N��]E���'6#�R!�V����Ŋ��ra#�RiӋ�d;)��&(Q�]�����u"��������T~'d�:�*S?)� 8뒔W?���>��-2]���&�'(f8��Bmy�Ya�JS8`a��1����ds��Z�J���+���^����7Ьq�La��f�W�n!�w'��SV��qu�fCtmD���uY�K#���cl��4x�"���<pO��h#��il�)�Oa�{�b����Ֆ��N�IJ���I�����c펕te[���6pdxdD��-Rrj�uxذI�z����$ͯS�ޒ(��xk�1���K9��ߋ�׀.w7\�̢�	�VS���4~]�9vlNx�lّ�p�#�X"8h	󥞎�c����3[��ڄ5��M�����0j�5�B����!Ј��s���S�=��z��A�}ť�0�a��^$�t��i?P{��ռ p�����C��}9��[�.�UXf�'��mRG����iI��4/%P0�]ͺ�&�=�婫�R|���8L��������*�f�}��w��x%+���`A�ؒ;��^1�K���X�f^�;|G�y��=����xb����薁��b>fķ)��%�d}+{��|o:���������>ۤ����,����9�I�޶�ԩQq�{�&�T0:���,�닗��W�LR�޵m���"CC]�������zⰓ[��͠O�y�lƗ]��.��i���]� h�0�><qVQ��S�$}�N7~����FO`�.Z�����E !�kS`�S���)��A������__H88T�D��/x������Z`��D�}{�.+�ԱhP`{P�S0�Y*��1<���U���Ӗ��&.-=��YǍc�RəE+w��j�����ջ/:��$�1���9H�.V�S"���C~���Ɋ���g4�"l���kA�>�,��6��w�EϢO����GN�U,���F:�z<�/�R�op�X��(��3\�w���d�E��z6�7X�d�%�5v��Hv��aR/l�=N�)�&톛���t���[\����i���sͮ�C�8�P��CM�$������������"F�MT�-@:�s�"�9�Ql�[	(�y�I\9�_���v��\���8	ZH� go��WbU�cN�I�ݦy���4�7=���6J�~�=�(xmk�0Njч��{j�����p��=�(�?#�n�p�}j�)ٔT�ҙ-�m������f�*�b��� �m�����PR|p�t*��"�Mۂ�~��� �gw򂲑Bi��*�
]Ond�Tq�^N�"�oo�4Ze՛hW�N��.3`�)���x��hP�!p�`�E�Z���N��2��c1�̖�Pw�iy%@X# v�ư�Y�7�!Nj��}�(��ޣ9Ӛ��2b|�Sܙ��}�Nz��Y��Q���Y����]�Bɂ w�8#Q呤p�^�eW?��zx	�����Ivj���pw]�u^�K�]>_���xQ��H$��g���\�ݿч�	=3n�<?vղ�p��4���$��>FwU�{���Q�M��)��ۏ�*���_��H�פ��H?��!R�Ɛ8���Ҋx�+����yб��?|+�����S=(T"K�`�@lL�����U��E!V;������|S���E���jw0%��:$V�3���c.���8�o�i:W��Y,������;32ǳ����B:��0'@��j�O����.�4SH��
� �8�g�[S����]�k~�p��,.�/b�u^�a���)�C
�Q��N����i��o8JK���њD�N-���)��}V�=�ʙ?����K����[lz�Do���`�����z�n؜yQ�t�b6$A\���8�ScO��Q��&Z�(�v^4D%KB��36��d@V�8�Y���j<H�fB����|�$�GWx>�̋#�+gwR�/Z�R���X�~Y��f��9�ݚ����Q��CA�H�58�6Σ�F-���&���ޱ�1�\�v��uC�P��d�n�ȵd�y<,J�C6%��ddpJ��!�T�Y�T��ן������M�r�nKC�lm����B.@�X�B� Dkn���/J����kf����g������H�΅ݦf���fO�^��"б�f�����v+�.�)8*d�ф�pĦ�j����g�c}.�pŸ����Xs��Æ�ÏR���b\�9���S<��#�2.�3�-�l�*��y!�m����O�u��^������I�������"Y�=)0�v?���6�Gr�/q�	�����z��/~�[��]��⇻f�b�7��%��0��1�ép�r�qQ�ƾ+�
�싎�)�Yo�o%�S��,B�W��,�0M��ox��>�Z���8B�'�,��l���=�_'�9/������6G���Ymn��>�%N��bF
�".F����	�8�\N*�(ߣ;7?����oگ��}�z�M�l������!,Κ>���8�8�,�u(�21�T�<=���l`+����#^Ab	ݿ����a�v�����0�%j��A���?v5�~��V%��N0�l���I�$f�I�����r��O�gJ�ؕ@>�^G���*�����)�^!�/"�G�5 [��P_��П���ן���m���7GSQנ�	�%#���mˠ؁��9��/��d(�K�:٧�,Wvni�Q�K�Eˋ�jf}�7w�l�,���ܪ⟊P���A9��Qf :�<�R��@�f{�m �����5yYoo�x�_@0צ�%�I�pJ�7m1b�e�^��1}���|�tn_�1|�k��EB>����m���q9�Qi�g��Z����M�lX"B?cV&�Q��a���RՃ�V��~ .�,J�ʡ{^����9�+�|?�+��W�-p�9��$����B���M�Lq&�06�e���G�E�RI�mR�����osh�wg�͗μ�({h�dH�@Ѻ\��D>@?��b���;�و�����?�M1�4��Jax_�GO��5�Q��� �}j�r�^"�6����E���l�E�(�-iLgC��&j��� g��y
�[� zj�.��e[/�Ef{���`���7�R���Uj�g�&�r?�{��fq>���z��u�e~VL�H�q;l��V�??B�|:w��aQd�%ͨ�fVz���Z��O�V��ߩC�t���`e{�F�.|��1oZE5�$c�	�T2�a,��;N'V�	�!R�k�������)�f���M"�/�W����
�%���n�;��\�<�\&V����}G�9��}���tW_�ط�+|��V`��'!MO�S�-�nB����T�/:�6ȟD���nl�=ꓐ�� ?�cSb���@�Ag�����<r,�2s~Q�T��Ļ��5�2\���PûuD��(�֦�C�b���I�+�9�-�@
&�6�鍁�g�6�rF%.j��o����o�(]ˮ��}n�Y�58��hX���ۊ�OJݰ���y+ͭk�����(tG�S�z��O&��hh(J��	�V�uD��r>2j�4��%�1�e�஻)�����n��Y�����2=T�G���5m�A5E`^ɬϏ���F��6 ���O�^���DS������M૗ꍹ��z��@�J�i����vY�Ģ�TV��z]Y��e��v?� a���*���#��îV������O5�?�g��+m\rq7�V�Y�'q�Rx�O�}�O�-�jd"DD�����&�*g�}�<]!~@n��1i�	�~c�W����y��[���H���J��Y{�h:t���Ө��n0��)]��^S���$��r?�j�]���*�!�L�2�s�(ZP�Kb�4�T���X��6a��>q�h��PujQwt� �0�_��2J��kʦ˦hXy����vx\��i����
[�``�[]�X#�L0K^��P��]����o*����N��@��m}�"#�F���ݽ�._�t_��о�.fT�����'�+��]�,� Jr�:�b�e��&��MXd�&n��9,m\ e+�3^ϊf'��Ú&�� �j5�h��'"�J0��1��(������:��+yi�B�X*����J/5P��mD�⵺���A��:�D�xl?N��Ei�&#� ��Z/��|{��LR�7��ju������&(~�`�t������v�l6C�a˦��5h�l��(�����μ�N(���T�^y~�+7(����kzn4۟ok�	4J>���nRk�����Q�:�9�tv��/6�&��.]�ָf}*�3lr;�Z�P��ȝ��1{���X87	�Ӆ�T�
�-(���;C]춴!Ink�/АC}CE�Xf󔋲�L�߁{';����xc�&��&��A���u`�)_�Z��t˦Ka�R��� �Z�%Vh>J�X@��]�Rg�>�)2͹�ׇ��>',Ƽ͠NC�m��ۅ�>�������J�<M
�/�+��0m.�h�{�l����UM/��������h3�vۅ�F$��9�t����x���-Al�cK�k��X���h�a���_���\�fL��1N8���e �_� �����K�:ӗ��33����he�����^�{�彻#Z���Lw@�kU���.��^�+z5~(�5���|��������I+�{ ���c�F
n3fA�]��G�}���7�&t���b�����gˍV�IG�����ol �s��Wِ9���-��f��r�$�����^,$ �qlAm��C�;�F�|��=I�G2�e@����J=�ip�a-����;�S��K��3.B��<@��@\6LMf��紲-	!�OF��I	fy+�0�<8���@J�N5(W�|WO�W�R�&�G�\��=B:־�/<�$�0�sk��đ$�O��3�LF��\)�G���߄Ű�P��o�~P�c=�]4�z��e+�͵$�F�C@����'�T�����@�V�솎I������U�e�����Sk�+�cO�4q��g�߈T��|нm�;v�t�{�ɶ�^�N4�o*ܧ���)�D�L�D��{r�}�F�~2et�]����_n��y�0ٲ��Q^�8��y�o���Q����<m_]0Ss�7��}��B9m^��N���V��>�t��}���=��u� �H�V���@�2Ꮲ���9�ￖ����6�5~Og���%�R��ƫ��̈́g�/������۴Y.p%o��:��S6�������H��88&w���^ǖr�v�t�G�2�=����ؒ�~�������R:
B9�f�u��=���9�>��g����l|�}����5Ta�Y�zD���0c^�n;ַ��^�R�e��
SI3O_�a�b�B��J4y�g"��zy\rn�S����k-�"��T�C��r�Q��Q�V+����z@06�F�u���$�Yn�x��Ͳ��Fe�X�L������n�6��F�����wb�����?p�|�M
��0����K�*�;�z�H����������A��g�;
׫6�1
��^��O��6�X����y�t�y ������i6
�'G2�&t�ǛcyW�����(@�]\�T��'L�\���[)��c�a����.6@�1����\ȸ����`�#=v��X}o�$U~9�Kb��G���2vٝ���!J���ąM/��gm+�5#����押�C����7�2x����>xӲ����^���1^���|�:�o7�]�5�-����\���e#" �w�@���Ǐ�>�b�?��F�[��'x��ÓS{t������v��������
%�r э�VD:�	�YIW���nǯ�[)2i�S���Ǘ����1�EƣF�-aa�S��d��jO�D�s���ƗmN��#���nNGsYlA�5\�n|п��Ϡ+��P��/</]���$�_ئ$6$�Qg�����(�XT��D#�d�;�����I֥X��A[�ME�*���d1t����M���f�"	x�=�'Ț�ٌ��{�������pB��Įb^#�b�)x��� }�S�'���a0չ'F'	��;"�Vzu����H���y�g�_P��N��aF4v�t�e��$2�mQ�h5��֙�#���8=����]��Aؽ��w���
9YA]�s,�A��{��~Ј�����#�5�է#�CvgM��nv=��}$��k��]�������n\�Yy�~���R�Sǟ�%+��3;���J
އ�jț7�ρ7l<����HzlCH���^>o75��o��6��@O����pKeh��i����ڦ��&a|n�y��5�a$O�.-`���L�o��Eh��Ol��\z�������M��RH_��:���)�|���������iWQ�鷌��o�_K8�ix&L�K�,S#�����pقNt�dL��{�H����2tмQ>E\ 8S��;�8<Y�y�ّ�G:S1��KY0Y�ۉPd+�Gܸ%��I݉�7��SQ����}��핺�W/2�*��uZ����V1vE�������Xv����\޲8l���U�Y��	�Z~��^��T���׽:,�c��&����������j������^)��p����A�^I�s����7��e��4�2P����V��duk��$��.��,�\�~�'�A��7Y��Eu�x]�-�й	��f񺦯�_�;���7qx��h��d�l�����!Q�#�RD�Ư�~|gf��W�k��7C�b�V�,��B���f���G �v��l{W�=T]�\JB�L��}��вJR#F��z�1C����ׯ�6O1�p��i"�z�� ��HK��&�a��,r\g�C(�4�_Q�>c&�f�9��]�dL1�ށ�yHu�۱H�<;���1IL|�m]l��D m�Fpո��q�˭����H71���Oa F��!���O�I�����9��2�{�F4�PK���S�֕a�^ӈ�O�G�~PTT��/FBX�_��O�3��JoLWWY�/�^D4Rv�A�(.4��صڲ���X�� (y��a�8e_��6O�]oA���%����=��F�i�(��� T�n��8�.�� JX��o<����Q_�Z�̟2�mΝ�k��,Ӌ��M]}I��ΨDTn�7Z>��ԦF�ͧ�c)\!7ƫ�x�!�gx4W�z�(~esn��Z;V`��X\���~��|E�D�ww�w�?��l�M�*�����	�[��i<��_"���+��=_�Ǩ�|��w��7�7����7�Ў�cOEʲ@��F�\Ȼ��I�ƭ��X>mU/�x^�M�%>dW#&AAA�����3��5�Hb���Jf���o�wS��`哺�8%<�.n��G@8-(@��`K�����5��M�e^s�W���0���mO�LB���z"�z�C�V����zY�S@b��ސl��'�,<ٛ���X��<��:Y��� \ ���*��'�K�\����uT�����.��V�g�������퓚�q�j�n��=
8L�O� ��������Ka��� �	�����U�9��κ���,��PS��.q<�����Oo@4[���
�!��9�������Q������� ��Ls�F���6���E��а��l5LH�)r�Ņ�(�ڏyZ�H�����z�h��@P.�؋���}�55�@��Q�=�E�׀<�Z���>}����j�Z��x.o�ec֘��i�}p��!�]nf�KCٯ]�t�է�6�n��$�([��w��x�zc�F:d[�\c�;?Ʌ! ���Ͼ����E�,e��Ik�����v9�(f�A�&d�]���2��ΠZ[���d)�z�
d�y�� �[�y����S��^n�t��EY�g8Q�!w��G.�c���i��̏Z��싎�DA��J�����rȾ+yO�~E�
`@rm�=wg��u�С��s*��v�I:���3���z��d�<��[�����o�?����&�Tv��t��q��1�J�tA�7ςC�O!%�Ґi���-3�T3�n���^B���px�3�2ABsC�v.b�4�"�|��?|T��C�+���6P�H�U,��3f����`D�B�6����v$�M��8X�]Y,�NM�\�((5���Q�|{d���j'�G��C����i^D���K��`�)�������!a�
��R;�hI�|�F4(�$�ys�=�r`A.���9�P�n��� �b����~=���
��j��=�����\�o��=nٗz�iCn�~x��.��$�F�#�䒼���h�����<��c!؄�y����;͇"�I^��&s����E�8ĆB��&���(T��'��hO�rl��Z�1s�e6�%x��N[kqU�g��B7�_�QhZ+qˈo)];5��и�m-Q��]o�j��2|�����+��*�d���=V�m�&-�贆��CȜ�׏���� &��k)/=?���#&���Z7����e�5E�5��Y�=И,a}����ك-�Ou����g���!3�GA��;QT/At�����K� <���@�P��a7�(�q=%�c����]�~�eT{�w���o�"�_h�@A!���W$��#��MD�S؆��#(X��D-�by����yF:R�	��[���2?X_)R�7��_(+L�Ҿ�zDB�pK�za۾�Tz����oA�#�|��=��v㏞�
$ �t��B]@n#e*&��r���?��VDf�C|h6����n0����MzÚ��q!��T�Z���uwA�>�8�8�C,�煮�t~;%t�f�9l|���8'|����{s��5��h�v�0N'�A��&��H������#��O ~�Y�ש}
��l0��!��ΰr� ʧ�|��1��:�pMWF&M'����Z�fkު{�Qg��fN�Cy�"�����[��e��|N�t�6�ި\�$X̰|w��X?=�k�q�ώ�S��y�}����ʷ��ln*�CT�hd~�t>j	|2�7�t?`Kj�m5K ��M�i�7�U���=_�Nt.
�I�Y�����3d�7铠f�$��0V\;��P<:���xDp����5�9Y��{��@�f��(M-�Bt����#�}�*8Ox	�`��dH�{�U���3+3�f�[Ȣ�]Ӱt�$~�&�	<J�r�6;�d�KP*c�DkR����WW�Ӫ������v�y���ZĒ�i�0��M����Un/}��R�i��#u&��4��q���I���g-<�O��x7$�e����Ȋ��ϸ��_`��;��LM��ӴE�;-�`Pg���d���Zy����+bO0�7�yCx.��sF�g/Ȧ�}>�s�戱���������r��܀Iɯg�+d��4[Z�[��{gUS��͝��φ�g+	�=��Q�m�Lx��Q�Y�YJ=����#h5z����Լ(+�'!��g3���28'!����у"�R���A��^C�M�����F9�y����7�����A�=cK����A��Mw��᝕5�E킛O]c���������F�qmt��E��6��k��u-��F�J���-o�>/�A�?��I�ux����ı�VQ��H��OH�������Q��3��� �%���Ƣ���lђB�x��{����3�q���<���2��(���%�њ�1�@oTku�|�_~�X�ȿ4�65�ż���}�ؔ�<0dʔ.�$a�z��}��?�$�8�����|��mr��}*y�VR�x.�����vfЭ� -2/�]�;z���������Wמv�.*ؔ¢�������y�������"�?Q�c�]���g.�UI+!���߫�9���Rz��Q����5+��w��K�V$�]��Ufx�m!̲��"�r_a�w=��g���j�-0�~�F�2��z=oi.����� �ry��8�V��8^E�5,;�@A	/�zv@��$�|���#%Az"
~��}#p6��/�f�F�N���ϑǝ{�4xЉ�NZ��W%�5���fD1��2ӕn.���3���CJ���B4�̆���eT�ץ�dn�G��<,l�b�s�&�Dc����ѭIz���5����dvE*Z��O	����E�Ƽ����ϖ���Ar��YK_s�q��s�hj{��-� :��\��v�������Hf �q��nj�D�?�{�K�SU���J���c��Ɲ3Y�N�.\���������3����&f:0��ǁ�1�{�~ط*����}8���_�i�rq4G/��0��8j~�(�?_��D���:�t�b���4�]"Q�c��Q�����0����<z���ehA����Wx?[��)c���JǮ��_�t�^����VV�����B�s4�����ȝ��mL��Q|�xk3PD��'��Ұ%{I�Q��I��?�17�O��M��gt+�bƗ؅�E�^4��Y�����u4z��^�
�."R�x�B'��_u �i����2��Z��@7�M�;/����Ӧ�ŧ8XZ�ذ�-��k�\��ԑc:��w�K�<��i@�l:�CNf��mDF2���z��s?ۧ�p*-N�n7>9��ap�Y�YUI���1����pl4=�R�9ٖ5G�E-AG4�t�w��Ce��=F{���?��˟�8���Q�,x~&���fW�d^��jwT����ɹa2ҹk��;1����5�V$��ex����Y��{���H���;g��{Zgr��C���?��t_e0�� S�bCL������S�.ږ[.�@�1�����i�y�>�,w�A��; u��s�M�?w�ei��q��$c�n��k�.��ss�1��j�uZ'�IIF��n&d��%�lg���P����KI�c����6)���)%��Ep��Η�Q��Cv�!n�!f�}!~�{;�TE$*�l�j ��qBP49��\���Yx0������@
`Ύ���l��Emɓ�iʶ�jj)d��#V�F[DL��v�iO���x�# Q�]��9*��b�c�w�|�I ~�'�V��Iw�9�G�����u;���7LA�`)C�<->�?>����2��rOeGC��R�9�Zl��5!��hAKù���w�!yY�R���d?��
�Z�W�ٸ� d&B���SU�%`g�ΰN��;�Bb�az���!u�v�I���z��qLf�>EM9�ۅJ.��pK�[M�A6t���x=�_�V����4�|q޹*q��������� �)+Q/Z[p���O=W��?(˔���2��������ආ�~��t�od��BD���%���׍��p�j]W'y��1�nQ���7�%�!� ݈�� %闖z�.�������n`�������y����u�ϺW< ��N�#yj�&&��������r =���WRj�ct�ڔf�?[�r"��8�-}�M;ZV9��u�;ڮ�p����&�=�r����d����V�����S9s
����c䪃��kyLT_�iv_���N�)�:J���6�Y�s
Z]�ګ끍zf�Qs3���_�n���2�Ly�VvL��y��u<8�[�"��M�_ _�H�i�EE�� 	V�&)�'�\��,������x�]��4�Xj?D8*��I�2�����U2-h�!�[�[�[\ڛ7.��wr�?He�'��=���R��`T��@
������֯���c�M���(�]�6���.�����m�Tr��N?�bri��j�xg���GD�҆��)8Ѯ�U��-zy�{�d���.��3mf{�|��3���c��л�3��B�gclvWV�0�J��.N)���$�f����)u����c��NT� q@w���́e�������BGIY���&Q=�?�L/+��w%�Tn,+���!o62��6������蕆�gX<tPZ�w��&��qG6��N��Ǣq�������;8<��`4�.E��G]<���m���k�D�
�Z�T��C{3�!�����ب�VkKɆ��T�]�!�H;yFc;��r�e	B�EÅ��)85%�g��7�#�ݎd���>5(13��{��prT#��"��l�Kp�J�c���Ԥ��!ғj�3�����Q�!�\.f�%�H.��oT�ϋU[yBΟM"m��Bn��KRe���1W������)��\i�L��;��e$��^��ve�VK�VN5�l��/7�jL|�C4���F	�-Q3l8�����"6(��*�����v��O��7'�|�5�:ST��82[Q���R��� ]#�^��F1��v�|�_����hוyVR����F~�E��oԹm��f��á�j~4BY�:H�?����Pn����_�t��0�[!&ټ�;'Y��'�AC������y�l�P�.Ec�(�Cw�d���UP���͵��J
f��{%����+��)J���y��u��\�,	X���d����G�{���tAQt������ԨۋIc��;_xm���_ǈ��9/�ܜm�Aq��A�.�X�����	1��&���cam�z�.���:��UK���r\��0��l�BǍ�q��"OJ*��L�Ƙ���r�M��j!ps
����/��ҌFPb�o~�t�^����iǋ��w���`�z�/u��m�~�YI��%��͚�"%��41�x��k�\�L�Al]�J���Ȯ��(�r.�t�.Y�h6�Y}X>W�@�]�Q:+׈���!���	��c��O�Wߺe�`)P屜A`bD8� �_�`@�;�e։�OSL�H{\h[���kh��=S�.�|������Z*��H��WӅ���d5DF�(�:恉C��zw"�:����M�o���ag�����klΟjS{�؋:O���m�7��fY8_�ea��Ж�K�Y�Eƫu�t�]L��T�Oa�}D����**�����b�o����[޲U���!i�����[��s��)ы�_�LƇh�K=��54�X:ns�/���@�Lg��|�nm`"q�74�v�ӨpJ�1��W��ωIJ#�x>�X���4D��8���g�9��|��\3����\�'%��K G���ܫ9{�86V#�0\��#M$Ѿ�D5o�-o�vY����s���_�ն�3���3�C�87�^ޛ�;(���m������J2�t_�!���5+b  9J��_쓅C�c��20?��?<���*������)>�7���j�����Ich,hM�������ǿt�R�X�a��/Ð��o($��P���A�A r��*M�⟔t�1���!+�'�W���1'|��lc�
S�������׶e/l��o�����T��!ex�~����w�lS{|77Y��$�y�@�tf;D���N�d�������l�W�5��������zw�'٭�����G�׭i�͊!��3�U�)�;����>��]م��/͘W^2�.���*uU?���~m"?�1�.ޘ��c�LdoUA�X6R�:��(���W�_�}�2�x��
��FV�_���ȉ�E\��u��a4���q{-i	��m52��P��!i�rq��`K�s�/���|+��tu���T{7�_���qz�-�4�C�C]$EQ���\Hulc��{c)&&6�Tj�����wo��oR��^�Zfq�J)��u*��+��t k�����8'��o��2�߬�T�p×U#LwKƄ��yX}��b'���KZhӥRRp����;���I�TH���=a �;ڰ|n$�-~��담73��O�z�� n��m�8� n�{�m��=������P���ۿ]n�N)����tQ�-�=v�dVnXe�ޑ�h�ĝ��*�T�t�N�[?�wb>� _ʸ�}�ff㿑ڬ3z�x	���5��{ƒ����i���"� Ռ���أ�	�T�%�|'�˦�/��kkk-��.�� l9���f�`꿫S����h2T����ﾟr_���\�^^�0��<�Ey�P�0��;{饲��W� }��=�r�)�|V6q=?W<�/����z�\{�7e�K��o1��V���s��P�Z��G���ԫ=��[)ۯ���(sY�PgO=2�i��<8��*�hG6K�q�W���_>.9������J�R�k�>T]��d[K
+��g`�?�$�^Ja�`	��`۶�
��4�-�/�v�{(^]���[1�u�'r�~<�H���<V�����X������}*;}TJ�',e4��H��O��s5��I��'þ��>���̓S�T~��9$.ۜ�R�^&��Ɛ��k�۸��,����J��ْ�Rϥ\�S����G�l̧U.�/�>�2��!>�k�^�L�1�JLZ��7�������-�.k��kR�@v���,��_�b�]�u�o���d?:��sHm��n��=�ܰ2��Y���hx��r�^!�3�c�Q�d=�J_��5�s������@�A��<���y�c7M�9_nv�y�0�AO:��b���n��$A�{?���><���'���ۆ��	���_�.�e�6j��
�P0=I�D�J�֜�)B3��s%��&Dw {�보[ùÎ�a�D�O
��W�~���Y���{�q꾯)`�s|��(�ΐ����څ�e�Ӣ��k�ϛ���������g�� ;N���S(hwdA�(*�����CުvwALNI��2�~˳1;��hB��8@�$�:.���GK�Q�fT�8�_�Vo�ɱ��~ԓ�&�����{��5�:QҐ��3y��!/x�u�(��wr����&�B����`P�}��;Q�j	*����~�2�׈i�àT���ZZZ��OHb�^���Xκ�jM^:F�"��Qɽ����ׇ�F1oٜSoEX�0��e*�R����|��:߽i�����h�D�=á(���6��&�@�~a���q�k���D�O�����A�[�ѧ%�e�Y��_e �Ɍ!h�X��n	:���%Fh0���?n��űi��0<�5�L7����:����&�JrьN���Fi���G��x�7l~ҕnZz}�v;a��7���h��kHj(,��I�(V�`�D���h��}��`�ٖ�/�;������}�^[�>d�Ћ��|�Mظ���ozގ�7x ��`#k՝#>���w�qZ"�����
O������Vˎ�9����凸�g��²Q�j�{�U'���r.���EA4���� \_�^Z�=�D��D����q~,��^ndNNnN�%����fu2OD/���\}+�Wr�.d�S,p#�ui��>�^�'�!�a7#�1�=kRqT5]��}��6�D�]��'�*�=��W�'�=���ط	�w�9< ����k�����Az6���$D��";ڇOV��>o4ߞi�m���.��MVl0�����78�0��Y����@W����vMxML<]F��^�� [�r��?2��2�u�Py~�X	3���NTT�������7r���b͙NdK=S!Z�������#�T&u�����Ec��)[AX�
�S��^�dJ)$��I���n	�pp�
pX�
�(����0n��?�)��R�G:O7"��@t�âN�����_�"T��.�O1�˶T�O�-�E��6���C`�żk�LV5[�,	-f��2�[5����Ǚ�fT��,`�r���4b�+T@8�GR�{�
k�F�����4�|�0s������P�W��'U����-�Gg�&��{#�I�*���3�=����UY������W�W�kUYN�w���"����萶`�����^�/� ~O�)Z"%��1G�X���Z�x���H����c8�����|����)H�A�|����������h��ꋈ:I�8�f�v��\	��!tw���~�B�	���r�������#F#�/ut�!Ai�s-\�*/�K# j�1�J�} �,*��?7���1q6~+Y�&�����v1'��qa�y̸l���[l3���4�I>a؋܏�,7:���/�ֿ�F�C�a]>�N�3�vo"�R����7�{���p�~�;Y�e�M{r�׷ ��S��o�3$&�:��
>?2pwIG��4z�Q>�� �:�`��:s� �[y�)��E������^�\������n����4����0�j�b9=�5���#���o�G��x�����,��Iة:�ʣ�u�������NlQ�W�i���B�������F�P�"[ m0)�7�ǣ· ,�P���;25#C'�M|��gV�`��9{~@��L'���R`NW�j�r��@�`�K�,���4�����dE��?O��~����S�-Q�kg�j���QKv(�i1��O�8���3���:���5���i%���^pB"���s���%U�[�E<����Jc\�|b~W��케k��]�dn���^,ϗ,g��/7���K�w-�c^��R�3�ӭ�@S�m
 e�A���Q �yV��S���:�ޙ�v�� ���Y+bs��9�
9(�"�<�1��-�W��B7����|p���H*���Ct��O
;���'"�-2<�y����Bp\ԼeS���d"{&�d���ӿ��I���A�M�y}ῶ�?���"R����T;'ϲ�����Zэ��.W�>��U�ǪJ��+M��Mcv�"ݻ���U������1w�|a�����]���:���9���c*oX�ȴ��@@��D�}[ �t!E+��22��N�I�CY ���E ����h��
g��ڋ�L$ϋ^N���c9+%BJu�)��z1���=u>����?�h|�挍��VT��r�h�I�4��Y��Z*c·54I*��ș,�+����l'f
ڻy��֡�;��H+��Xj�P����(�|�F���ݠO�{{It��N/�IH�ew,�SO�=ջ]3ŗd��12��o�|-u��ɪB���x�=�=�GaO!V��&i�73�)n Ma�r�oǆ�1�۹�7�[o�"*�?�;6�*��y$ɉ
V�[��B�Ҹ�� ��7�<��}G��꫰t�����Y��&I}/�H����4x���#v�����n3�՜<�r I�C���Mn.Mj,���q��c�PW��Cŕ�eYJ x�clig��C�/��l}K�@]$�U��`��4�G�do�H�d,��ұ�����~{����õ$b�mP����֬��c�΢ٕm0�jDCʩ��O���D��2�⠻���U]%�5c�'�U�ٖo�&��tw�������~��v�-Q�n�����`��>�?����e����\�����l���4�K�rh�:w�[��ޫ��N�^je�rG���V�j3Q��k|"}8�0�H}㹰��i��L�ju�U���m��F��"9w,;8�MZ����6�I��U�9t58�'���Xt ���YkOLG5�2,9mp��0�]��0� �ɛ��SDA�IB�0n�a'��d,|a�$�z����A7�;��aHT��*�ϒ!TM2	V�ko��-�J,!�co����w�H����������b6��شB�����ΨH	�/&>r(�7�'?��ρ���b�:�!^=�������K<�%��nz8�ֺ�7�K�&,StW�i]��\���M8h�����Cߏ�׺�:�ٙ>L:��p�d��;����[}�i�G�}!�]�϶XW��>+�/�<ёz�e+���~�o��qc5�d-T����vʏ��Մ����i�N��vC.v� @� gϜ'5 �un}���1x��t2!�l���4~�7�+�7F*�fC��)�|j���o^9mC�4�~
]@! .�1F�Y�U^�Uz�q�M::�xHL)����@]r��.�0���	-f:������o��ؔ���?��	D�3�F1�b��C�+/�nNg�`�F�>��9I�s���aL�d����/��j-�G�w�V_�ݥ�,h��/a�h0���"iL��O�1&�})()��2�*IQE톫>�jB>w�8Yd�pY쪱�9�y5��">Qk�֓$��~�i[U%���9*���dt���n%43����{[��材��=9�1��vH|����$�ٕ���VɹSY�B�_��+T
�*��1�l��uf~��h�|z'WK�f��Ȧa��fg�F���ģ�lK��L�_L�'z;��ic�`������uB���Cq,~��]-�����a�+��57^�4��8�M�Ď�r�n��5�)[�8j�Ɉ����mg#6z��4����#8yf�
	d��'<_lZZi�`B�p;��
�������:-��d�*�Y��1Ź|k�Ȥ{���-�P_�M�f�ѐ��Ire|48Ak�q�l�����~}L�\��o'�9-��c�9�&�o��X���	M]�lOn96�Oz��=p\H�eZsWul�T�ރϹIa�+�b�H��h����pa=k��}���<)�+~ �J;�\K��iQa{����+�%��������X;�#�)�E�p<<@נ�ݓUb	�Ü�]�Qf�v	8���3/DD=��C2of�	fVᴲ�h�h���j7�j->�~P*�+����uG��3��Gԥ]�_�2s���p|/C/���b�+2-��GbA��=�ʢulo����	�(F��[0��۷r	��;&�Ϩ=T~魐�3ք�P9
�9�k����z��L�M@��\3-��1q��6�3G֥��'^ 8����8+SEe_�ެpX�o�������mP&hv4��d��?~.��KΚN�r���ۧ E�I=���&렗�S1�#���S�ҡ�Zp��k�<ς�jǤc�b\�Lљ��O�ҫΆo<�����.���ש}���"�v�$	�۠7�;�7}!�ŹO2([��Yn�c�Tj��}���]�w<j?�(�����?���2�9Z.y�0�O;$��-��Mw0D�5��6y�M��|���y��9�<�g?��LV��P��ꐏ��U����]�i��/�+44����f
�m�m �[�8K%�y"b�p�}c#V�*:���WV�;�� 4Wߴ�ïw)����%�����Lb���[M�K�¶��_l��:?�HW$��Ritu+��`�_�s�``٠�7?�u�u���aw-�)��N!^kg\��g�F�TO�(����#$Y=Ev�#L�?�X���_xNkO[�g}y���ȍZ��<7m~���|B���|k�N�r��G��৷���H4������s�$�WD���C�o����H�Nk��i۾�K�{��NH�~68�Դ4���(|�Mu�]����w�z������K���uX���#��U �6����0	�������{0Vr�b6kϿ&�!`�{TJ	�ʦ��cʝf���wu8�;J5W���R��������U?�WlyKS��\�����0���{���{��j&�,\��X��-�r�W�-����4<'�8�~Z�bd�0εr�b�+��%���S���>��ٺ�3��5�}TS�I���c�E���\^Y����{9i?�}4ۃ=j�k_&	�\Vwd�+ܰ+��M��������p�n�������< �+]A�U��j�#i��9ٓ��@����&P�s��;pѳ~�L�X��q��j�"&��?S-���@�v!� ������ߒzZ�_��A4y�9�����2m�A��.��h�¿C� ;{���,h�l����4Ht�/FV�������[5��\ݰ��bq�"i�l'� u�b���~z��k�m"����D�T��ؗ[jcR�ȳƠ�k9ˠ&k�I���2ޜ�$ԣ�د�ݮ���6����:n_�a��I�i����wt��b8�{!t�)h[k�����߯�J:���2�G����V� �g������M14���+�d�S����e�]˝�EPת����z�z��9�`Q�{����8�aϲ�q4���HB����o�W����J!�&�͎vܾ�V &���7_��"z)�e�_�fvƶ
i��<����6TZu�O[w]�3�|r�F��J{�9�ڈ)��s����|oM7!�1��N�y��b�W|��V758"���Y�=�����h.��g�1zo��|f�����V�.���;7�"M�I�b���hU;��8#�Wr�7:^�������o�a��M���z�T���&A�rAG��l��Ewܳ�g�O�Şq�FM����z>�OMA����n<>�C[+L�b�ϧ
Q��R"]�S'5��!ݤ��a`�c�������!�*�fV��qf��l=A��U��Q����y�x�����YGX{����].���%�%���U�ɸTv�^���mf0�w����--�~$..�&~�k��8�fmD��`�=��"%�����U[D�E��
F4A��@t�}7����Sӊ�ʛX]|�o��F��!�LM�QI�ɱ��kI��.���Ձmd��9C�C��Y���֔��!�n���T=V�o���wQ�Ce�d�b��j��!���:[�nx�Q�٬BH߃�~F_�F��-'(� �k"Nͼ���[3?���j���S1�Ik�``Xw:�.�ƁMq[j�\O�?r�u`'¬�<<���]ϫ��57(�{>�lS��IA��,�%���V��DU�_�f,�R��?��L�K���ʌ����v�����8pwh�����2t;n�i�����v>x
����)x
(��`D���n;&i�~�Og�L�}�x��>��UKI�M�?�
�dX�0U�u�ױ-�I���v�(<r�+?��]�{Pf^��V��ewm��;�V�eM̝y�S�0�"��/�E>�n�� �s�|�46{t��||�g�8۞�p���<=3_�g	���8vW��7�W������5G��Ȏj@\�����c^�: ��:���G��|/�� ��$8f#o�?Ƚ������@o��m�?��@h��$����	���ݛ-��=���������~�E������/h�-����?u��9HV ]	]�x�og�ޜ �
���Ζtc���s�9�]���B3���/��`��JY�Q������(U<\�js�7{��L��V&�gS(�+E} ��͍�ѮN��J%���g/�6O:�RU��?k���h�!�����r����~R�=8�RѝEoj��E��9օH�&ED�&^U|�J�X��O\��B�_#H1'�gK�f�r��;��=8=Ӟ�$޴I"3`G�]f��l��\�NТ���A�Qq���U(�p�eWxL�Q�)���6�;y/���Z��>�ˊ٧̝��Կ�	R|t��:`U?�+������T?�l�z.~��jK��5�Im��$��S��L�N�W������R7��l��x���q�z}��z[�py-��e���b��I��і#�f@��opq5����q��y�����mS�'���kv�}������3�$?��Y�v�]+�H��Z-v�3�}��EH�� �h:@EX�&�����:W�g���r��]'T�+�i�#���с�{mc��返1M�UR�+��b�늪�dd��gȬ����@
,Y�,�L�훤�����+����;�6��8�!I�p� �ᴅ�o,�Z{�����+��s�����B��7��wS+��g""���`�������e�;q��!�����f�vp�&���|u0��p����$�Q
�~bE}�
�μHĺMKK�]��~.F�#5�Zj��
A�{��%x���Z��Xo@�J1�ri�΃�g ,a���a�2O��V��.�I5Nd�-���:M���b�b9���,Z��@��}(�E�Y�@����?|U��sa��ٷ��U�;H�	0�s�������x�EB�q�6���G���������Ay��M���tD���-������^�3���VRKn�Fi���)��ʁ���ܠþ����6�}���mXe��IkB���>2Զ�����'��������KV�Dj�W�>+C�+ۦ�N.d��ʙ����b�:@�*|f0�������վFW@�t�]=���*���[�7��W��y��=�ȼx�FD��k�&RLK{�\��!�t�~tA�V{�n6�5,v
+�"�b���N_Q�'IR��i��sgT~TP	c�;Ƭ�K
�:�t+ߴ\@S�{Ծu�W�{�nU��k�p�Y��������+������̸����1��7��Ǳ�Y�\�ox�~���z��֌�E��KH�j<^�Չƒ?<+g]�^���>f�즦y�7ɭn�K�M*7�3�S�;��I_���>0�d���w���V	�c����RQ�8h�}J�ɞ���ߴJ�0SR`Y��H���+yf�h[N�����З� ����:b��7���ݍB����}!�'tf�M퓰��c���C ��t±��ZS0D8�fD�xz����rgh�R���;�KM��TD�`��{qB<t��MR2�JV2> d�n؝��Sq����	ӏ�v��/%6�b�j�b�޾݁ݯɂ���-���u�JI�$xj{;�V�܎�7��>�"g:���^�����������C�/�x��:�tY��$��+�ּr�<L�^�h31(�1��O��W�3Q�U�w�\U�� ���c���k�ac������!���E0���.Np�
w*�f@�}���I=�$�&�V!�SBc�0K���AZ�\�x�R+.�HR�}*4:��G�����N�"����fT�b��[����ෟ����y]��oV��Ǌ��{���#�ֲ׿�_OV��O���>x=&=Y�j��Ǭ�~q�o�2��_4NL�ib-#�D��@�|�Y#u �J���nqbv��0jvVW[���P��_��������h@TXIZg�fI�����ԥ��Ư, �ه��.���FW��� ub�X���F���A^����F��d}f�mJ��} �S��~"rC}]�Ipy���%�糺���ɇgg=z[F��2�x�6���<��m��������h����[=֖��	���Y����A�Dʤ	<�(��%^9�"Z�B��v˵�+� ��gg��X��%��/&`K������=��1�*_9-:'���)^�`�O:W�+VH3���|�|�ȁY�0��W�%���gU�)��<����}�*���@��9Y�0��y�z���W;��E?��yZ)�a"1��jOU���`�o���5���ԍ���j��Y�e��j��b?����o0¬�b��Nj`O�.��m�@俲$��q���=٫�``| ���x����2���0�ckGL��[ş�V�H���^/���ds �+����8�-O��v��0f��K�a�'D�B��%�A�N��c��[&*��������o9T�a��8�Be����v����qn�Wˌ�7���5^�����Or��kɸ=N
�Y!��� �!o��oU�(�`w_,��do��3a ��o�X�:A�'LQB�0����n)��>#��S�Е{K"�͡&>YA�;��WUQ5_+����]HiF+�[�3M;��oZ`�������g0?X��m��mȳa [�K�|�Ñ�|#ch���^�	���/���\K@E�L�l������9!��~�>����(A�!�$�f������ l��C����=���4(^�Y?.��{�	M\����4�o7�E,����y���z�����,	Uzei���?�������!t��1�Rg@��k��xaE��{���c��u�v�`���ܮ?Pu_k\��x5��0h�����J�ϬV���#m�Rd�quSaw�j�g|W��������e|0�~r��\��t��T8w��\�(�R�W[Z{���	w��oƘ��Ȕr^�I�E+餗,��8/�U�|͞?��MY�v��..���~S딙j\��m��#<���v��z����^;��C0��:��en�N_��az%��y��X*O���l��9f�>�|����Xa)f�}}�$�ߢo5$���rQKik}��`"��f�+r~]ZC�p�!�)���bF�w�~8[�� ����.B�7����	���3=�Wć����S-�,��3~���V;�{�`��uΪ���O�s��>˝i��f�g=��)�� ��"�
��э��C@鋏1T����H�d�|�U��S<��Vs��x��D�C�f�fj
2�)D�wv�F�KH=�s^%/۞��F�W8߷�����\�`���'�3*ȖI�7��G���l���Pϰ�����;��ȡ;�έÆ|>Kq�w��G�,�c�v^v�S�Z��nٸ���V��Bd�RuR�j��M,yW��<�8�mi�T�%���S������(<�X�̬+���9j��>��å�#L�?��M�bNX.wp�9;�}�qO��&i����;��"�0^�ed���2i��+Z*N#�/���x�M��#��hX���M��;.�hlV�<�\��9����0H�M]�cᩣ߿�R�$7NL������خ�N1D�-�!�Y!�p��z�ޤ�`�����V!������[�[U5hMYI��桵�7.�ڃ^vqmMqg�ø|�f�,u#�{�^�3sЮh@5����� ��Rg���yS/`�wZ�WJj���?�Mm�n��9����x�$���m'4JK�R��ýR�"^�	�B�������ng(�|+!}<a�}�S{�Z��63��_���^K�jIbC�?��
��W[-0#Rd���8�˾�Gk�,ĮN����U�W+և	�Ŷ�'�����CN2�T� Y�/��m�EP���j�i��U`�@]>���oKZ���B̧�Dc�����lBR(�!��b��G�@��M�L��ܙ��<��l��~� ��c�].�±��ˤ�������ۧ���)���+�Z�я����S�LD+/8��)b��z~ң�x:S���p�n��+1/�X2��'�#�r}�����mW���c�o�;l>�ĥ�����a���uݘty,=��+[�Y�7�r5ZI��nX���^T��*�C��~�a�OrXa����_vV���
}q�ѯ$��0����ޞx�x����$�S�Xe�-�ܘv�,+�k�����k�yc�:c�7S)��/��PJ�V��c�eq�,��_�g��>RN&Y|��R1�-'ygn R*���U��
�)�GMu��z-d���Va6��@��Q�k}>�%�y�<Aܸ v��s�R���)v�	�J���I
��[�R�hH󾰵��G�������9��`�@�D����E켟<^���1�����/P�k��N2�ы�ݚ�*����{��xoc�X���.-Q^,p�*]�X���2��m�V�X ��)�G��X�,C���A�z�. Mį�y�&����
%q>`ATf�7�3��=��ݔ�>ޤp�<��c���/� |�j�!�-	��+�1�	 .F�Kve��#b��;1d����t�t�U0A�{ʦ��M�
�dr�_��p8;F��_�t�O՞~�|�����G
(������A7L�gx���ɸl֡�MXD�Q���i����;h�盭�=kX����?_,vR�o���	�u��k�z���U�Ǹ�w�FI�h�ri�)�,�Z�4���)\e�u��(x��c0��W��J�'��3��Xe|��cp�Tڄ�"H%�М!��3�骧'�Q���`�@��q>Ҏ!����kCXH[fa���m�p�߰�<�'P����&�¬��e�Rw="���kʍKD���^r�����^������>M��( �ۓ�M�1}��Zg��e�!�lU�q�({�,�Ϧ���(Q7��6�\��X ��͹���p$�!ު,�3����rL_Q��`�2�')�n
g���O�d�M�3
��	=�:��l���̰0�>��{
�:N�Ab�p����5��tSƥXη(�|����⹻����$���kT�R�Ps��0�ȉ����7�����t�������A��_��op�%�Yl�����2���WlX
���}%��ٚ׿�Q�.�J�¯`��d'��-�x-l���)�)_�Ddq���O�/�hα#Sx�[��l��r��iOЄ*+�@���q�d�	}L�V�r �AƺZæ'�v��.��G�N2�;;�4�π;�i�U�*�����qw�^γG����R�,���BA�:f'����D��(����f��='��/���-�Q��P��V��aG�%��G�o�J�3�ͫ��o�y���x|����|DT쥙��С�����\O�΄&��
ݪ�b.�����R�R�HG�ɝ���ZĦ��}MIf�m#��_�ˈ>�%
@��` Z'�[6�[�.s����Z��癗�~j�]�>���ϟ�ؚ��_�2�Ս� }^g��$�/�^��Z׏���v�pk��)wk�e���:��~��2d��F:��q|�]�����m�q��N��*�:@z�Q�Z)�N}���[g6_|i��Z�o�L;7er�X���X_9�#r�ׅ�v�f8���a���a�B&_`�%�:���_��5�������Gh>�N�t�y�e:ĽP')�>�R$ �I..�sC����83�WV��N���]�c��mC������-"3¸����u�{'�Sjj�-G��P/:�5M��H���� �o&И`�QLYLɎ�BGB�wr׾�K����,PiQLٮ�������� ܣ`���6�Oct�Ə�~��)3���S�N}��1d�7v�/m3�,��4�f�x�������&�e{`D�[.(�[�OQN�s��M����umL�����#�u�y4��z�����xH�X��XG6�Qoux��k�]�\�!��7�Ѡ��K�`ש�cM|�)���	��P�!HL�"�_�\T\V��`Ē�'+`��woF� 7#7p��P���}���B�k���o�k-�Q��x�$�~ �M|�'������f�豑V+򽩖ʖ��lr��u�7}Yh�D�6�C�V�C|�|˹�3%^�T��&r��� a1b���صb̸^
�k%��3�%v��`\�>��݁C],�f��Ӡ_E|ʯ<e!�H�X��?����3��xf�  z�q�	r=1�5���?�B�6޸�&���y�M4��;�߼�]�>�O�fy�D�W<��f�-%�*����H�$��U����.�.����2���\R�bS�w��C�aӌ��t��L0+�z�H�hZ�Ln�1(���cbk��cb�xw�s�_��N�I� 4�����UHS�c�'����9]+�a�.Z�i<�a�1I=;�Ira�riS��x��9õ���(�b��~�_l��I�l�Ro4w 5S��3r*�A9����2.�8����,�Dz1[?����򳷁�zÊJ��)�+�Y��|��$�Ɋ�=QN���0����ګ��thQ�����&2�˓ҹVy����K�Y�2�㍱��4��80W����*�R����L|L&���#�Ӭ{��c�-�`�.�iPT���%��C@:����.�B����:������{ι�a?k��Z���Ѻ��E��O�ܩ�ut]�6|3=���6���T���F��v?c*��u�$`��������|^:h���,>G����~�þ�y)/��s5d���;�5�ym+ Yv�IT�h͕h�����1�2'��G��<�u�eN~����4�b2P:��Ĺy��C� ��_W�sl�z�ߖ�K�U�	G;��9�9�R�r���{E����.�!K�y���mG��-g��d��J��!�π�>�'$ L	L>��*Ŗy�v�=J�yP:�d�9F����Z�T\)�ع�Y`��Ǽ��	vh���۳�R��l)�[/+?���4+�e+�p���H'�3R:��L}=�n.�2N��e����1�x��z �?��-#�#z��*�����>��z):��M��c�;�m��LV�����r3��Q��i�Z%7��)�Q�r?�|v�2��4�ۥ�,2R��_vLۼ��ڊ���՚[�g>�Zl�3�]T�M����2�K�G{\���PU����;�$�����D3ߤMvV��տH��hS�5Ӻ���r�+zz�7z���k��������mb�]�ϡ�i��?�	&�sK=�璣�ʔ�_�E��Ɣޜ�9�ߚ���T�#��
��9�e��a��>�,�9$���U�.�ӹ�R5QS'�|�9�gf��B&܏U���y7�:�>&G�$���0M�C��^az<��锸����f>��>F��3��F���Z���`�����X�}�_)1��$^����WU�)���f�����
 �/ϓn�q��Q#8|߱DF`��zHُ6��i��?p���=��'�����<g�0 �r��j��Z!���HT.��I������{������5�0Ō��Yr\�=$9�ŪX���tb����9��~����y�H��녻��������\uW�r�b��ͺ�`N��zr��������8�W�B�uq�ʞlNt��x%���K���v�)�'+NxD7�=\{m8+]���J�H�؛�L��K^��rX ���Ĩ���$噖��k�K�͟Ǵ���P��|�%;fUQ��� `E�<#�؉��D5�?�\��k�I%���q�t�???#!͉F�G��,�%7��Ȫ�M�b��[l\��?1����M�vUm�En\����=[�-βxu.*3=$�S��M�$��.�:��XO�9E���m�J�}!�����zގYX�����1�
.�@�o�2J����X��F��&]��IM޾һm���Q��<*����pS�ۇ�!�w���Vif[�$$�~GT�x��5��n���1x��Y4IKa��H��״��:��2"��5�IK���/-O���U�Cx�K�_	�~�͊��?�W#��x�#�V��9R-�0�M�� ��P])�2}6��0/�\YQN�yўUjQtک�Q�=�4��-X�ܪ@Nna�Ś��b�(	)A­5���ɸm&HӉ�#q�C6@�+1�G~~���:T���Vg�	�<��"��D\�-v�{��v�'}L���+��J8�P��*���5MR���`q��P�$F��m��B�`�P��ѷI�ۡb������yA��zF�������M�ǃ�ɜK+G4�n�\�����棑�ę����U����!5��m|�ϛ�.���(]S�D�X��P��D�K� �'j�}��%��V�u6S�1��x�XC.��7/s�34?�Q8�G��ł�x�e����#32�b��wX}/�����V���oJL�R�4�4��%hj�
�	>��V��77�;v��.�$�N:S�㳦z��Z�td�#��E=��m}��������/�{�iX������#-��&�y�k�"�O*��B��-N��!��HLB}}tma^�ق����,:(��E;fG��~���s��9���|���I2���RʾX^Z4i_�f
�XE_�Q@7�5%������<�Ąr�����	M����ԧ�' � ��\�|t�V�^��rΔ��oQz�7��M��MU�*�K#�K�����%Ca8�<D[.$�a�Jj��`L�r��s�7��.$	�W�����so�$���v�7u)���70N��B)���oѓ�x�>a�����اzh+� �v�t�`J
����#����$U�&��i��,)x�&����ږ"f���V}-n��uf 7�ڨ@S	{����Ƚ�SI5�ј���0�;�y�2�����3-���m+:U��%U@�䷣��Ċh�$,l�^@��I�	H7���ے�A]�\N�9�n
��h�����M�
��ʮ�I��J�gs�'׃�����Y���FC���ULy��UŒ�mM3j�I�#1g_?�7����3�{��+)�� �?�*K���L m�l���O�$ -�_<��Og�ԅS��:�d��CE͊D��S����ɪqkl|���9G@�����������n�b=�I��g��E�^����A�(�|�0���jQ�������ϞĒ&��V��)�+)DX��;������Zp�ܪ����A]Q�0��(b�ג��Ό��*�a��H��,�N��qn.�S�7��xz�����w(x�����'��b\c��!��_u���d�y&�v90l���lu]^�V���I��1�)�z�c��U���`�HR5�U'��D�'
@/�/�ʋZ*A��c'@^���d�����������r��μ)�Ӵ�4�	�.ܺ������CH=м��C�֓��k��M�;����A,B�!a�6e�_Uk�{k|�L�\���ߊ� 4�>[J�
���&c�Y6d y�34���aQ��Rl��(�wz�y�ɞpy���/Q�0�E��s�S��'633�LX@�'�G0��.��:$���{�^{��O����P�{-\$����ɍ����8:�8��>{�S�@��������D2l��ȳ�iW~�
Uͯ����
ɬQ�yn�Y(�"���U�_*�1i����:[H�/ ���HZ�9�3~�X}�h�y,�؛�����Qv�?j(��BQ|�<󔲸(���p^-�U�1����_�V��{&��~͊0N���q�f�B���o.���/��-��_c�d���#b���**փY�(J���s���;�9��#��КN-L#�]�2�x�""�q������֨��WG1֢������}��~�}�����Γ������g�K�V�t;�V��o���~������w��I�A{e��0W�o�񨿿2v+6^|�5��Qw^yW	Sb��������f�%�s"�:Ր>!��V�l܋D���x�/R6�7�i�W_�ǙY3����%ϙ�a��|�rS�(]"^������d�JH�B�kG�s��;`�P��j����"ad��&b�K_��-��|f����2�7<X�-â�"��'��xj��|׌C��MB	2z�����mw�z�ǥ6җBV0~��p݇1�ms��]��$:8��Bd[Tn��!�9�ߏ�RET�����߃|Ge�L��hV��w�Z���	����*�x(�t��x�}��Mٱ��>:Ƒ{�a|A0�δI��q���ex|Տ^���۔Hd֗�'�w�2���	�{����#����K#���p����T����Hq�~3\>iA(����Z���xo����vG\�[��ʅC/�Mf��Y`��2����8��V7��_ȘV���`�����$�'Z��}�^��T��V�S��RO._&
��LB�KǨ�r��B�Ag������,��&�t��b���q�H/�U�����K'��Y�d%X�H_��GJ�cp��l�v���(��R[�S޾#!�-�2W:�O�k��NC�^Je����	�#w�JP���8��������kO`%��;���&f�3;��p9W�����x��0I�qp6��i9�U��!��<f���-�����=�j��ҘT���~� ����s��g`|Y��?��<�}����o��L���P���b�9�� �������֔�8��1d����4�p�3�!/B�˶^���5
�4ٹ�ʹ�Z8H���]f*�*��0���dc�q=�������k_�i?����3���ʅ��*�����&XQ��gpAO�+��`���Si�>����OL
Z�;�,n�r:�)�9��-�����2Ӛ�q�h�]�4[�
Q����]���!��cZ�ޛIćDS&��笁h�Vv���"�n�t��iԲ�V����'���=l���ř��MV�PD˜iPf8�UN"��d�����z��F_�&�����pX��RO��d�|���R��t�k���3����a�9��oc�����{@`s7��\��m}�/��D��#���P�X�_F"�����z�A��η��'G^�㳍Z���n����cH�GN�1�K)�O�F%"B�T '���-�|P/J� �=ܺ��8kjs/ͭ��$,Z�꺌�d�4��j� �^*S���}m��~ �n�D�ߴ>�u���Vj>g���������*��%_t�6����=�E,�,T�h{M�^6�D����Tϋ��0zaxx|>%=�A�ѳ�+��G���1����Sye��Hz*[���~Fo��dp���0�촘�,�Z(SH�ڷ]x-�J����9�i$!Y"
T$QH��x����j�aT��fo8��&$2���*l,�T����zÊ��h	'�I��<s9��V�|�}g_������|�7 8�
�h�S�:^��1��V��-��<aA�B�bZ�l���Ȩ`�M�(��Wd��
G�L{����X��뀒����g�$�1JxS�؊�#�܇AK\k�����r�J�Ȑ,S4��bJ8��yt�;Y�b=�����9� a=��o�B�m�=�n$���wES�����ہI��B�䮴��ŋ����d����}p�Pj_�Vq;�a�����Mډ�k�h$n���}_� �g��Ȱ#�y�@'�:�<�䌚�ԧj�&o��Lj��g��Y�
��Z�^fJ���nQjј}��ǫ`ʑg��'EB
����>�'�M"3P���&r�0u68��!u�)��d�̈́)��=f	�T����������^�i�
���/�B����GD�D�Rtn����uN<w���I�7�m#�����9v�W��)�&��̪����>�wS�	�F�w�Y������,�1�!���c��w�?�<�z�X݅�n	a��ʾ�}���_�Ϸ$?8���)u�ؠ�\dOU�� �{�0��Z�r͖�RN+E�{�k��Xr����	��g�k����g�ރ-fC$1&��GgU���[$t�6��2��F�K�5Sa���?�1�|Q����
�k��>��Ƙ�{�
���h�+
�+<^�9��V�ڃ���%�9Y�'1<A�V��e+�s�T���z/_3$������m����FF�}�������]���Z� ��1�C',I�j��q�g<]�`��l��M��#��y���r�y5T��#�'v���N�,>^%z!.�X��v\H�S>�� �E��]��,���)��}��������)���2U�2����{D�����Y�t���F[Ѳ�]V �4����8��cq 2����}���[�i�d���?_A�*r���@?��f������JJ��/{��TL*��(kI�L@��I�+�,��]��Ԟ�����(���f!(ǒa@��+�tK��h��oִ�������SsL�:f�ݡxj�
����?����Lrr��������"EK#W����2s���	�)�DZ��㰤a��Ti�M*���6�A��u����
�&��/�2�lv?�Ox~���@�!+�-�Ļ��e�������_m�5K��+�qi�����b'��דor�xk�j���ҽ5�Ҕ�PU�I����a��e~:������Ƀ0pWv*�T����7|��6�yM��<܎����|B�_��@�U���I�%��.H�~>���yJT����u?��$p���=%k��j��R6������¯�|��-[ο�{	�����2?sђY���@`�p)����es��-��p~z:���O�"�\tAq/��ya
�h�u}"�l���ʚ��C^N�URb���Cg���*Ё~����/�Nצͦ��T�$#LY��:���=�6wMT�#mA�\��$�lQ�W���b�(���c�����c���a����w�#�K���5L.�+���\D�}�U�o�D�2@ʧ�jɍ��sh�Ͱ�Z�����ظ��R�g�7g��}���o�d�@*9�	]�C�g����g?���@:�VO���R:��r�����0�4�����?������� Q�?� abj^:[�	Ὗ'����@ꬉǲ��J�R�px�O���잜�� �l|�.?i�|;�c�9���i�tjQð��.��"z1i����yOE4�#ȋ��$khҪqߟ^����25Ӈ����8�f�w��%���1���P uH�XKx�}B��w�*,{�M֕�w���G�@��@��Qj�O�Ǡ�c�XR���F_�A[���u��}�p6Ӹ~%U�?�wx�Ck�,�_[%fNM�bB��(�����p�r}�&�"�ow�=���~j��=W�eu�ya�h����vm�5o����v�����٬�$�2�=��q�^�9R�⸌�Z>{_�fO��ꌭI�g���#�;
DOv{�@�+��U[1o;֥�<�׽��? r���ճ�!}��e~2�9T(�m��ǭ�8Fg.#8.�p�D ���j;����x���n�s=�s�㔹Z0'�/���\
a_��"�#=��W��HGОAp�,bY=[x��	�����=~7�g���~��6�M�޼�Z%�A���ͻ��"w���%}�W,j���pR��><ҤCD}�D�� ]�H���IT�2&,@7ҷ�Ƃ�����xƲ1 Οs��(���A�!���������;N��N�36�-i�������VW��Z(C#�]�`^�TTV~^;�lu�]���?��Uy*2��]�+A�����z|�����uYe
��,U�4���
&e��_Y]%w�5�p`��__�m%b��[[��-������`��{��g����`/��b�'� H���a��2lw-��'�h	����A�/�\�����+���Hp|?�KO[d]vU~�ǆi�(�,3���"E%���ϡeѳ��@p��1�������)�%�(-���XI�j�:����';eV�[���Np�/Td�1w�޸�� ��˔'ӡ}J�?���T7n�ւFB�(�b<A4��!��O��S�JF�\�?��<�\��� #��(ٔ���b��5*�q'j՟�[�S�hZ�&��l!�/�[>k�Qv3��!,�i,N�Y����B���~L�(��jS��kÅ�劺��N������弹)�n���c`�ws���w�=VZB&��S�b^5�%��vɎ�)u	���� ��D�A�(��_jn���u~���#���3GU�L�����Lyq�Cq&R�!@�wBp�W�?	,��,��8zdag��I�A/�9��x�<�����<�	�E�h���2۪������؊�����SJ�t����M~�_�@֣��e�%��Ma�QB�B���KO�P�ݠ�dӪ؞g?����#V���M�r��D�gL���T��b5���_P�_wditV�����T��6XArjLȥ���<�VE���sK��)�O5Jφrx~������q*����Z���(,�c���qf��+�b6��٢���_\�yItw���~�:/�#�x��-��>\�Y(�z�N��!0����Y�G���k/�{�ʠ�u��]��^����W+�J��
���>���9㠯<���6gW+$�Z����v1��kVb/��X�t+*�2�fa?��VRD��$ݾ}<�u��2P�To���5I�� �H�S��6B(��J���?w��W����|��;�������N�>g\t�n
p���)����$��)�)�'b�>S*Z%D��>�M�}z�������YF�%�CV�����1���s)c��"'{��#�T87�>Ԛ"ܞp��0]C��3�}� Җ�+	2��5N���o�x�z"�n'�^gD�q2����8�4���0E�9sn�8�'sf��(��<����^�[ZK��e�om��ʲ���q?�=�'	ح��Nww�������ACNZ�����5�Ckk�϶)ROVZ�U��0�W\��Y��w�,�b�Ri�h�	Kp��	�l(��r;=�4��Ek-�����qr�tFb�A���\�\�Pp��\g�j[lH��%xc#l ��fI��B�����MO�Ћ؉�yxMA�6"��Wu�0�e\۫� 웿t�� =�)ӯm���V�me�_kc��.|UfS�����Ym���!z�xOUU����I^�_��A[$�5�6n�N�	�Z�&kk�w�d_��9^���۹~ܧ��m�$�6N'ӰZ�%ջ���7W�Z�[u�Ii96��-t�"���&��{|�45Po���9�R�6O{?_I�Z�w��`t�a�4On���F}��>���!H��l���í����z3��j�b<'1�$-�Â���z��b,Hy�����̎"�%�dQzLS$8��h;��,.�G�W�A2�
�(0-%�&E;��4��+M�1>��O�4L2]=.F���N�+!��'R�rJ���yym˻��ړ���������V�:��p�س�x��O]��������ճ��`��S�>QD��(ˍbP���p��$=����mz.*"};���8�Q�����=i�����aN��J�1�u�����Ŕ�3�f��:�%�[x�a���+L��ޢ��0K��Z��x6����<ǳ���6��sWNB��ƛ`z��>Z�7�mm��TO�
�./_���7���s������.y�r�)�ǃ=��CE9��r�/��9�~�k�W�I��2���)�vl-כ|98!��,S��)�Ȍk�����R� �Zu��2������p=>�ת�a_��2����5*Y���ܸ�F2��p�ǙW�(S��
WH�o�5����Y5�y[e���:�ۗ���ccw�nۭ[��4>a��r���+�H������:P��K�G{Ǜ�5�U
O���"BG���V[�>����q2J+�o>($s>,��u���ͱ������Q�C�9��ju���7��%_bXк��A��Y����i�f+�n�瓋����x~m����t��F��b�?��I2$f�"/�/�OBP%����}U3�+W�UVR�)s6���Ó��k��\Zj�tk��V^<�S�� f}s}�D)_�p�6��Ŷt��L�TZ6��LCw��������b�䳄���d��o:5g�݄�-[l���'��h7�k������]����ݙ��9j������z���NLw��$ -/`~�y�5��\��/�; 3A���WѸ�-fU��Z^�@s �[��F���a�����\8��� 1���� �Ub�l�.���Π��
j���Լ�q�ς��s�CQ�N�'vo�����>𩡩���.����̑�ʤ�hGF|+���`I�t��1ﮂ��/t ���f8KuDd�_PU���侇n�����5MRn?��I�%�4^���E��g��[�� !B����O�cUO�Li�d��6�*t�ca�?쨬HB��!N�}�/�{�,X�b����QoY��tw��5bZ�������aP�����������\͟��IȪ�V��� �M`�R�/���qʳ�_��=�#��Ć��;uUjۏ|�"H�a��v��n}c����a��;�/|��U��pS>^4��@�:W�Q�4�ي�& r��Ӂ���~�}J?[�5�q�dy?+cg=&�z��4��9l���;�>�U,$E��!�gB��V6�i-%j��=h�l�N�B���1���l�K�H��K�E���l�6A�Q��=��
\��kG[���$��G����~{����N�J�%��JPC�h�;�65}���)�{Er��da�L��1U��G c�|,ǹ���[c�H�'`l9�і��� ��g`�J�Z#�2\=�Nf��8PPx/��Cn�yxW�(;��a%ڲu�ք5���m���� ��ՕYq�Q�+(`IN��S�3��/�x	�2��J���[�}X
܋F���R�9R1W���T� ���<�	��}�Z�x�F������H�4˭#�C4ձ��U~����C�DE�z�rw\7V�p�loϵ�I.��u7O�m[�`X4�?ē�x�<��ĴZ+_2_ȝx5���[c�W�XW1��Ik��bA�%�waJkFD�˜��w.�������S_[E��i��yJ�X®/�ǫ�3�6Z-��n���_��X�"C�D�6Y`�Zc�"���������k��L0w��_��fX��6*�!s�go[{�N�_�Yu��&�w�x�Z ��ea�� >�>v)��󨩱�3lк�6��Ƕ�Yk�#J2e�
������h�?=��}w����-s>湶�'~����3�q�
ؠ��&��A�?{t`�Nx~sѥ�� ����n�kX�?���IlS.�+�a�.�����Q��wi�N �҂�qM�?Hvŏ�ɷi}������v|h���i������T�z��~�p�*�7��S��:Ԇ��+��h�7nq�.��0}�NyV�G�Ny�t�<+��%^o���C�/���)d+@��B�� �7_O�o��t�.��!8lQ��L+���a+�����j�i�o�=��I� `u��#�S瘵)�)����ߔ�z��bb9��Qr�e!��j���I���\2�׈e�֒q޹��Ƈ[���&�>u�:�ko]�����#���u<s0���M̙֣�w5V��]���P���L:�yr;fdgR���]V*�����0�yS��dt�+Ny�R\z�d��ٿF�U�"f��4�4w&�H� !�/��)�!���/#����Lx�S�C��b�����f8��_��M�Y%LX�~	�WsZ�h�JYP?
��v�44�!3K�cy�P|,����]���M�8���a��/
�s�B�6��k5���[�)$։mn�tr��P?1K,t��m�׏�i ���Mb�\��C�Hea%��u��||�D���B�p7�x��3�z.9�]�m�����ê��[z��)�DbWB�5�5뚀�~��}a���UT~d|�c�+���l��(�
{������y� *�>��`Ro�S��\x��	�j�]>9)~W|�`#=��B,���@z,��L㞗�&	�ٹL��4)��Gd�������4�h������1�U�c�ul�+~%��(�,��ض7Qu�皦��r4�����M�n�ĳ��W]��<o�)�VLWUw���	��kq�?ְZ�cpI�/�$i,4�c��/�^:ˇ��o-4}�E��K��a$�xl���N�/�Hţ�p>?�\J��P�8A+������ZQ�k'���5���z�"��S&�B;ted��p���3s3�xt#�˹V��ɍ��C�?ek�0���V�ػ�U/�u�FKs��9l~]s�lڞ��.Kc��\[hGU�[�b�Q�RkS;��+���W���l�g�NuRĞ�z�n<�E�[.�z^'ǳ[��B��2.��ypf���[�s�XT���"�����b��
��	'����(�B�<��{G��A�!2a
q+�~@R���p�wi�n�d1(pc�3�����{��7:�H�m�Wl#�|����lQ���M��q3�[�VpS�~S�$R���"Ll�U�@����T�a��I��j��f��O��e��]��AH֗ĸ�hʠ3�Gd3"O�䆸�������x̰ϗ�y�µ��x����d�'s�G��w9�T�tUZ�g��~{����%�����w�Tŭ�bm��'4s0I�㞸|�HM���!M�56�~S笟��������\��i�J�͋y��j������#"�ĶWy c�9�$��K�a�[���RLP@%��(��a
)�{'��/Z�I�lH�(��89g|�lVD?~&�0��_+�ښF����ߎ	����>Y����fy ����@�dn��n���/#�/�(�{��`E��6��\�v���٦C�����_P[ B]��yx�`��g��[>�p9���Ӌ�(Y�P��> ���l�X����jo�p�f����E9^[��N�ou�����p©�ZZ<?uF�(�[ba{���N�2
���(<�v��@-�[�p;\����� z9���6 � m!�������ǧo�-����ow$��)���E�C���#e�*�E�1,�r�ú�k��3��tgiݜ��z�nɌ�ث
ʓ|gw�ک���ӶBq�[���M�s�N�����t�1tܸOˤ�N��������Dw��{��q�����py����ne
i�������wOn��%�B<n2;P�K���R�E |�D�`�]n�!i�k�9f_gj.-p��MC�N /X���g�����C�y�M�QY�.�3u�r#�_V�&���,!w��%3e_"��gi*�U�L.)�(�IF?�H�~U�Y��عS]u�<F���(N�����EǪnf�+��IIyTx�y��(��ER0�T�j���� �23^�����������3����~�'d5R�m� �$��}:L���o�\m}�=�A��֦J����9%o����;k
�Ei4���W'��Q�~p�BEr��y�ˀ�ׅ�Ɯ��|W�){b�ﲥ�A.�j-��^�7��]�#�<����s#t�jn��Xl��\O���z��-��1g�p���
"2/�SQ�޽7^�$2P�,�>q[����:2���rօz� Œ�.��*�^�[\����a�c�,��\�ṝ���O�cYrj���wF9�q�5�]o�]�3(M�G���%��>�s9N�}n�d:��1(����˾�ˣ�A�v2/쑯��uT��Aq&�?�!0����T���|A���>�x���^s�ph�swK�{��d���N�2[3��2���əs����G��< V9A���F�#�ׅA���� ���j��{M��r�t �*��	�)O!���3��\o�q�]^_��v'���0l�O!T�a
3[��:�-�η�'�Jf+0;RvS� �n-�݁������5�:@M���v�G,��-T�S�h�5ܱ�nײ-�Ң�e�mM^��5����W���	��V�?.� W��M���Kӑ�����4R�����:I�P=g���~�'#V�%Q��c�f���2u���(�s%MO~��6��|��.y��KǸ� �?B加��&�K1&��~�7��	�k��0�ԝZ�_s5�����]����FS�y��m?�XQLi����U�[q�V���4ĝHhiay9����<�	��Y&���fx����P���t7㔩�V���O��"'s��Unr*q��%��S�i�o��3	Sm�Z�p���Mh���tGiU!mش~.oM��?p�YڌU�_K���+�Tc�-^	��9J��Ǵ���#�����:6�o����x8y���
�\K�K5A���<��_悚�fU6�e�+��+�_���7�ѵ?�+#\^�_��11ǟ��赖*�	4_�
�a}��*D�:+H����B���/췽��y�@��C�ob*���̬�Y�ȑ'����V�nr���U�_K���͒t�R��II����ri�Uнk��;5�w�c�9K +��`~��:�Mf,���$�����*z��A�y[��~�����8��x�;�zF9NM�m�l�����q	�#��$����8iCq�ޑb�+P`�;/���BKyL��er�|L)����X���>G͈O!�ID��\�>��Q5�|H�󉿃�9�T�
�DLe����9��\w�V���h�Cw2?
'�q����)��Qv���a]eKz��*#��d�Z��_���-5�$���p���A޼z�� 	�&�y��F���ǥT�A��>����Ak�R�q�mg����dH@Z�3���AB���&�,����.��\3z�[���������m���Ū��6P ���e)�x�F�MFNg�.ɞ���>f=���Ǉ(M%��^x~�"ɾ?�j5��4HTm��G��q�v���>��;���?��w���Zl�$�ZQ�7��:�g.W�q�:�J�f�b��^f���E�G��5����j��M븆0�ީԇ��e:���k%2�{U���!�s;������ٲ]�
�U6j<!�b��䘽f0�&�E�Uo�i���%�4r7��Ia�߃D�#�p#5����/I]�~ ��~=��T'�������W������
��O�.C
���t�l�Ӹx�ߤ+�<`���{��x�ޛ!�baf8Y-1�qF]�U$(}�0�����s���@_�>���M��"����5Z2"�a}A$�'51_s;�C9�٢H���>9YK}z��G����/���>�����Y/�b�!�d��f���K��(��j�J�i5���H������R�ө��j��I�5��+Bt��q�)~�AJ�SڶDn�f����[BrZ��bq���8�_4��!9Fx8�ϻ�i2C�M<���,����z$�Ě�v��:��*�hſ��I�N���՟�'H��x�qtm#�^j�c+�Nw���`z�P���;Ј\V��r�<f���7���O��L�T��0p8@���
H*��/!<o�ԙ����L5���t�,�SN�y�h�V5��:	*�����69�7��H��¿�� \����%��[Km����3�*�_Ab��Q"�ouJ��^/���&,.Jy�i�:A��oatw�C�t]v3<�r�에��y��^~7l(�oٹP�pC��0w4���u�ЛY|�)���!9�_JƲ�ךãg��S�I�w�y�d>��sa5\��ǏS}mۜ��ˎ�,oB�@�π�n���s�z�_ጎ��?^�0��Wt `L�<��)�ke6�&���ۇ��8�P�!���������	�d��rҺܽ� � ����ǹ�sZ�f좡~��On�=w87�2���W�S|O���ߚ�+���G� �k�g����
s��]��8��U���T9_�V��"��#u����h�01nNN�b�3gԧ���*�czS�:�͘�P5�����y���<�тG���y���9\^��otf�d.f��P�|�/8�$�7���~�IW�|�`��!���
�JOO�'٥/@b����J�;#�ɬ�:��OI��W2�ޛ�Q�s&;���h6�~ST��K�B�r�р�3=�>���Ž��U#����"��7�*��f�M�gB�+��O܄�T����.��''=�k�(�,�L>?ʽn��AP�A�1_2��Y���Z�l�v�sL�:�G��W�?Ȳ�	t�	F6��E�]���䚱�ĜMr]i���˛�Q���)Q���l8P#Y0�/�G5�'U�����P��7\�����R]Ջ�P��1�h�u���|	��%��84,vIj����AoT�*#��G��x�ͤ�\�͜��&Z�7m<���HB�W`��	�yBB�q��3$F0ro��/�E���Z˷%��f�K�K;"1�-��܎R1螗1�#ʆ�x:O���_�ޒ=�V���"s��}ܥ23�Vm�t�0.�����<%{9�t����桒�@H�C��P܌��[2����[�ٮP����ً��gBJ
]�W�{����y~��[-���/-�����,��G	�Q���r��T�vQ���~�I��w�G<��_�Þ{�Aם�g����.z@#�!5��aO�1��6K��)��˯�K3�+�*_S<2�/��_�(�<t�������<��6�������K���w"w,{k)΅=tەƨ�_��Џ
v������K�ޝş�9��IgE"w��tp�w�\߈Q�޿y�Y���������u����"���Z^����.4�x�)zdAW7����d�uH��e2�~i��ǁ{I���I�]�5Eg�?�*j��xǷ���m��3Yf��[g��Yl���VJX�N������by��BC��B`��?����Eߓ�I�X�0��Hxa�����������M�rx�t>�]�q�[���8(����V.cW�KkE%5j⤽~5�3X��:˨8�e[����w��N��ww���-�;��ݵ�ƭqҸ���x������s��f�Z����=�/��L̷B�g�ța�.��G�i0�e�kM�%y�* �knP+�4T�P=D0���8ǥ��}�!�$}�����$<r�E�"��Y^}1-�\�Fq�ÈN�w鍢�R��ѡ:1�r��;jK�DŹ	9�.G�uO���h��W�T�d#7��r��?K{-��}&Q�ڔ��Vri��v���Ζ&PTR�s�p���3E)�6�-2�Ce�bcN�D�Ƭ�*����/h��k �u婀�=��l:}m���v��x$�������~�L1��X�Z�^���Uh���`����7�gE�ϭ�Tm..��{$�ݯj��m)���0VH�{ͱ���?]�̾�x�e�Ǐ\�k���ۃ���?�t��.J8����,%Vlq_���h��M��Hט�eg�/��2|S��0���W�1��o��oI+M6�[��"I�L1��p��6-DP������̷�i(��أ43ˣQ�3�j�!Q#�M���\���k���������ͶT����_ü&�_����G��<��:I�Y��{`��ֆ�&�s06�J]@��`zz�=j/ӱ?�RɄ��vX�]�2��Y�v"l��{�%64s-�H3�����.[St3���-B]�*���ր&��R���)%��'��]aj=
5�����d�5aͱٖwx!?a�[�Ti{~��]=G\c(�� ��e�xB�2X����<Pd�z��G�JH5�roQ��������=�F�q��o�P
��$���Pw⺁�"��!te����Ӆ���c��26-6C�A4!T�_;(�g���>�7�Ƙ㷞��i-���j���FWx��EcՁ���,xE*�*�r�,��_���DWd�3�_>WYJ},BT�$�y��6�Նo��U��xX����F)��=_r���I������T�M���H eSJ�lz��gǰ@d�.�t�6�Z{��(�J��kEs�*���d�G!��[�ڇ��o�{/m" m�%>�ekM��}���\�7��"ړ*��  ���A�L퓈E�*h�>H��y��B�T��F,��3������@.��v��~�� x�1>B�UҴ�Ô�[�A��JV����LC��@� �1��dg7X8t����I�k��pr�!����$�����1D���KW��=o�b~�l͔���i�;6p��V	�7����s���0@�8����&�s��c)�W{ڌ)W��;�K_n�� ʀ_����8/���C�81|�^���گ'� ˙�ŧ3cM��u�]�����B(�C���A�l�;R�M�P����!�s����khY^mmA�؄S�V>�S�\Bm{��d���޼�#�Hv��m$k��5��<��3�VT���D�j��)b)/���:�&ҧ}>Y����svR	u�ɠO�DG<Mw�^�_�>���p�i������s� ��XZj��Cϕ�9�����3�oW>S `��|"eW�5���kѷ��d��Iتq��l��z����c3�L�.��
{�w��o�}vň�7{s�:z�XK�b�(ӰʨV����zx|�{����}oi{0n�r�"%�-�}��Hl]��#'�Tw|x�̩
߄'C���D���V2᥆F�C%��j�z�<�u3�^|]��;0�$�UX@4��s2cx�榨�j�q���/������l�b!n�M�3S�6Y�H�7�<�Y�/�%&�;�����RH`g�UlP�*B�i������3���������~��Z�v=K��E'[)H�8F����m�`���v �B�I}��[��B{F�s�t��$6{h>�'�S�C,1�/�5�ڋi�,���c�~� Bי��k���H-P�gD�	�Q���w��pZ��p����}WDّ*��a���i��2�Q�2s6�"���鶫�t�r�"$�nK I���8�$d�X��	b?�ͧA�h��;�`7�1+���X����kWC��_֢|�g'᠀�g8iHY^�1�Ϧb�u1�pu A��Į�<��AλԨ��k��l=�GZ����o�]q�:Z�Z��`U���MF� ��U����Z��\�e.�#��L��G�L�ޘ�P�������'S�//������Q/��X�j������� �d����)��r��/n�,�zH�8�Y��,���g<��.��`y�[���ƿel6��@p;�����e�N@n��F��@�1]������̚��*4���JP�S�%��	�2�B��bF�Z���#����es�у��0AEV�NP�q���O�X ����)�Wj��A)<�/k���6��Sw  �R����ːh��17;l�CZ7q(��#�>�{(��CD_qctw�5/��+���@(�;�2b,!�=j�?��l��K�L�꽉-��8�? �n/aVܮ�~�Q�,��7n���z4����w�6;�PN��z.��^�h$�#��m&7=�=b����E^ͺ�>�ʤ�+����!��i��d�b Q�
�|�j� a}��O�ʷAm��_��c�hk��c�M.�y�lY����	�>�4N�����J���$�ܯ���ų�|�R�U�߮8��(���g�����e��q.S��C��?r(/�1������k����w:�����)_����i���@Y��	�s�5R`)s���y~����S���?�w� ю��ߝ����7U���ʂc<;sc�c�	�oN�F���oD�z�oJ5i^mWØ�T�ؘ�=���:P���c0��|��	}py䗩`�m�/�GH��N��K���%�}��b_|ń��l�P����a��)�eË��Q{�E|K�U;s��geB�I�$-��E
�\�Vi�Y?�Eַ��1����O��w��g�e���;Zlb�D���C���,��Vm&յ�2-���d��0̿�\���A ����;aĴ�4k��ԧ4��� KJ[���U��5��;(��=��0�+c��a7�����]�Y~�j�|��|�A+�*i�a��t�>�U��d��U��t��i����.&�-��m�~�W�D�ǽ���AP ��Υǽ��,����V{����	LR|�NR�ԉ��M�uR|�,ͪU�,�6�YA����Q�L�yI�
�*_S�6jM�i��e�%_�ӴD�m�]5Q�z�Gd4M��r�~5[�f�hjwPv�Cʡ�*�N@�=#�/��"9��?w"P���6�&�)zY�e�e������
��'k��H�ko��A�:�M�l�QOub Y�j�vrɼ���ϥ�<M�,�9	�1�:��\�o9�b	���N��`Pс�kUBMj���m�Elt0�h����U�\û��Ğ7?��Ţ�QS8[��%���ڍ�7�<kW�{��ow�H�'��*�~�#2�7\��+#���i��A�8��`�����˴������v���ϭ�@���U�|P���i�,(}a�k�:=s&܅�g�K}����i��%b�uD)��r'f�	 ��7`%v�9�<�&2z���ۙ��/۶����'�@r�Y�$��>#�qX��"6���Ԙ���Ҩzt����_�2���d�+5AX��
�Pyԡ��ڍ��	��
XR�	�~�h���R����ܮ��	�¨���߁��'�Z�zR�����iwH�C�gP�������n�ox���X�ɮ�j��z������2�W��#u7iE1��<S���j��J(�
��h�/ch��܃��5;K���JC$58yC���#���e���0_Q�Q)��!�+@���S!^:���������/�i�*��n9/��R���u��l���m}�)�8��Uo��٨3 �{qO�R��@����r�b9�(�P!�� w�:,C�}�^��|���`�Y�� |���b�a�����O��3������w��N�r����iw7�ͭ�T]�5+��ʠ�+��vFF\��԰����Q *A��FC`�a~����z��$!�g��O:�F�7�� �;����
gld�;������'X~2��B�b�U�gK�s1/H/�����|���JA;�(ֻL�֋؄�6D,�k��B-�� �y��DߜҌ�0���f�1%^�yndc�v6���R�`t�6+�,QitY9���f�j���?������7�a��������e	��0�U��`�^H�{�ĵ���I?�z��]�ք����p��o�U
�}��0.Iw�3��2�����֭�<?7��({Ά�nW�&�"�"�rXA/?�T E͸ޙzS��y�އ$�?O��`�(�u��X2'X�XB��b��&)AĜ(N��:%3�2�B�R=Σ��B`k2�R�*u���B�ZJN�E�7{���8���Q�?�ޥM
0D�����f���b�%��X���Z,t�����A�u�_0"��\�|��S����`i��y�T��)��DU�`���9����[He��R����8��VB#�<�&y��� �������4�98X��3���]����N[|����1��:~Y	g��k<���d҃� Ȅ)�*?bé�Ġ4�����h�nn���he}:)M��ff<�`�����O>Z�̹ʤdc�Gd�.��l��a���tfʉ~�QT����I�^��� ��G<."�������Rq���*�]��� ��A�Z����#����1j�)����ݣ$�+�ZK�B�h`b�����'vP=�
�!BRT<��)x!@ÿ�D��_8��X\	x�neO��7�~q��~��ǇJ���m�����%^�����`��ۥ ���L�:�{�����R3SmѾG!8��� 9`1��˗O_I�N���ft���8��4��& ��������P����z���*�<�j�p�e�Щ��3�����?>>~D�I-�P�G���D�9��x�[u�(ח����8��Ժ=�F�e�g
�󤏄Vq��h���>�"�I�I���u3�S? �m�gc͕��X�d؁�kq���@a�#����O���GX%�Wt���e����0��2�?�N�EeFG�*IQ�~��s�$IbD\�<������<��:ք���ڨ���y��G�
jZH:<����!W�ޏ X4��ĠW�B�zR*��z*>�Nx�&b�J��:X�,8C��$��pJ����ǚ�)s�J����zJ��Z�.r�&xwqqo�v_���RZ�_0�/T���9�s�-C�HC��~���$�/�v�x{��Q�<�
����d4:ɓG�e���e\Uk o�O#T<������ҎO���e~�'�{�C�f�� \���\�b��rV�[��M;�_���{��,��Z{y���6�^&4�L��s}Y_V���͒W�J�5c���1Z�X��?C���1YV6l�U�7g7Дh�c�&v�jf"��-���&�;v��`c:�w�	8�T������2��6�W�)�d#�s��W+#���G�PJ}N}��iU&��7"��ag�H��ҝG�9�\�a�ʹ(9i�+���W(�՚*e|.���O�/ˉ�dp��8C��4]�;i����%,{�9����9KL;��[܉�#�X������z�'h+�+��ܶ���6A��I��"�:�Ȗ�z&�Ȃg�ƆM2�_�{?�R�wżق&ł��5�;�����S�T��x*���`L.|�N9]Ё��_G��S�{�P0�	�jģᔱ[$�P�a�-�M9*�%?��I��e�|�vcG��,ј൬ym�d�}�;X&`$�U�LQ��W�
��	
��l�M��J�]��}%��j�5����̑�Z�vO�,�2�V(U�rs��O�|��G�`��c$��nz�h�a�!L��q�A��v�OEͿU(���VX���ߜ���%U����?EVx��N:�Z}1!����b���k��Ob�۩����^�ʓ�d�44�I+���j83���y�	J�a-Qb����H"ˑ�-RF�����bL�<+w����$Ӝ��^%mx�'�b,�?���Z��%��;�`�(�ɮ_:������q	j��r��+���8[:�}Z��23SM6��2.ޤ�(+�@�.z����B���d{9j�����7ާo�/l+k��wM,W��%�we�G�|����9V�F�������6v��e�ꁱ����)j{{#�Pm�����.��Ox�R@� �㚧Q�����o���_�GgHޕ����v�cr��AT�a 9�t/ga����Q!�\�{,�-�A,I�4�۰��0L�f�%&j��,�_�Τ��{��Z<Y�8������iS��ԩg{�bv�|M���9�:����d.�J�bq���6w,�=�)*9I:6��S�A�°.׈'?��Zc�$i]������Z=��~��'!o�w9~��]s]�'�[��Z�oClW=I̠Pn�3'�ۄ�U�ty����K)寿�~��=�]q�Z����[X�zlZ� 0։���r���f��ύ\W�������e�0�������5;�2}t�9n���h���f�/�:f�?y��}+����i�_}�F�����:
[������Hl�iD�ݤ��K0fdd�
j���	�0��}@�nD$�o1������ hL�϶��4�x�4@��&'�]��|kC�2G��Gѽ��$�ze��
�ҤE4KP�7��6������!�CS��0�W�?v���b����&����0*��V0�ҿC��ЭwTb˅��l��eL7����៟��[��|_QM l�E]OG9l�Woۊ@㠷�q_�8�ׇ�*b������"�#��dT}�p�o���[#�9���1��Z�-ܒ�>'K�d9/a ��͗����g��G+��}�ܻ�zWn&���awԱ��2��B����4<�Ҏ�o��2H:Oal�|�<�x��򡖬��_�!�4� w5�������C�]G�FIa+t"<!ԙ`IIr�֟kd��[_	a!M�n#�.��{uN�]�RDN��BS'�db��J�N��_�ٛ�&�
�\���V
�gvڀZ@�� M�����Q����?�8������w�:�eCl7���c�X��s��J<���r�����%�E��y�U	������ɖ���yV^y{fR}�yM��7-uuz1ԓ/T:%�p�W�[3B ڍ�QF�
Uy �0ޜYh�%M$ �O��<w�/�Gm �,�M<�����4����?�?�bH�w��͝^���[�U���(_20�FGl}��fkz�]�%���2ym	�M�����s'/�T��s�Q�>\��ըK�ًT̵A+��C��#���i
%�顶j��!C2�E�^�L��B��ڡ��8�&�w�}rI��h[�s_oi�3�hP������r_,"�f���L�@�;A�>�Op�
Sp�nQ�j~o����dp�u{4tp�J�<y r8� y�V��N�G��J���dO�Y��ʂ9�M���0t�p��<_�Q���E?K[Q�a�)�VF�p<�������U%���	��#�,�]��,Z��Ť�d��`��
��]��O��{b�50���¢7q�9�i��(����$io�=�S6F�0�]�^���ݣ�tU}�,�X�?'���u��͏qDfa�@Z#.�*�2ػfw)�!�����y� +,x��H�{�M�kh��3-���-�ڭi����!=	�bK�c����J�κ2\	��f���d��"Ɇ�q3O�X��@?��5��CL�K�M��e��őÌ5B4��MA����9`e��3�:.�1�Q�j���PHqШu�4�#��	�s�9��C�l�J���L����b��\M0~�+k8-���V�,JN�y��kٴ�|_��[�$����|@C���וv���h��h;�h����k7��Mdi��������I;D����Ј�Z�� �j���8���a�0$�P�	�M��m�B�����gH�<�Z5'EH;P���:H�I��1MY�Ӓ���
+{�i�L�[�X�o$�����*�&ZaONl��y[wۥg3Io���"Q!uai�t��^!W3�P�����m]R���1�s!���"���a̞�� ���}��έ�,Ռ�94cT#�c�La���W!9S,�����v������8�öTY��S�����uU�"�ʎ9,Z�I�d���:�:վvq�X�!�3!'��4��,?=�N����bW#�m������y�ӳ
� ��qF$
os�%�iK�>��%Û�+�r]6E"���5A�Jz,ԁ�D��wy"�3E�b-���Kۊ���Y�lI�ya��'r��� �!1e���9*���5�ې�����%�woOd�N�ަ�!��gn���s'�:�8����7KE��i7�3i�����pN��b���x[E��Â�ZV����+�ϋZ�/z_^G��o>u�/�c��w����j1���|||�s�ok��(��H����{�rU�}\	�[��
z_a�a�mc�P\i����}�p�/��KBG��՟~83/E|	.	ƞ��luR�����e�|
i#Q����1�pv�p!�i0F�k��.�
>wp#0Y�N�V���.�6��_�����J�PZ������F���㺷�ww=������]�ͤ�&cC���e
�A`^�{6�|�uФ��[ʰB�*�ZgcGW��v��{��{��b語C�MI��vyI_�������Lq��j%z��H��j\f�Ź��R��yZY2DJ��:&T�Q�}S9|0r���ى�R5&�|L����]/�.�̌C�>��OdfH�����u2���m-y�j��h��x[O|����� �9Ǣr��y:����/N�>�����OyA��[5��Q�b3����pA����Aa���|�6��Ӿ�Q�+��Z���}�ር�5�l��q��K�\��'���yv��p��k>j����B���J��ܕ�g"&�Ö��U{�K{".ٵ�����3�90
e��ؚ�T�a���P]�{a[�h���A��/�' �t	[���c�dT�V����C9Y\��VNK��r�	���9��5���P�-#Z3
Ժ�'���"j��c�k����I��R��Zo�xf2��^ZM����6�@������ҍ>�@�BO��P��(4���:6�jqL�KR���tR y�w��i/��o����?Y��+벆w�@U/q�^i�'[��Cf�%��ɜlP��'�t���H�b�,��r���1��ݖ+�I6��+��I�\�$�̦�)_�:�����zƆ���zri�_���'�/RRO=c5ǥqI[���2E�$Y���c'�Z�̪�3�k�,6�[6qs��t		�&y����#1�i��Fu��zXO	�1��Lĩ�����!lI�hQ����H�Mmj G�m������fL���2��鍖����e��S�7���ׅjA ������°���_ŀ^����t"����V&���ߨ({�e��̫{�� �*_���3�:gY>�)��	�g�O_��m?�v�8����ڐ�t=WH�w������
��U��Y�/Ė�������e�!�� ZMv�����><q;/� SD4�8�����9q�9��?��?aix!$�g ����������K��cX��>��a�\��J7p3+O_���\'��i
�K���(����{��6� C����-<����TLgD�ĕe�[[�|�ę�z4�W��L'w\ql�*2׋����Y�%1����?�L�r6��o[
����h#�U�%�H����IGGbdue̸��Y7Q�Ԏ��u����%2T"� �Ȑ�e�vn�`�c�S|��[r��޺�������j���
�4$��:1�3%2�%T�o���y��H�b�֣�:4	��S(#���'-r����$
ݹ��� h{sp��7�\����"���3��+��|sу���Q>���:���'�ޜ�+D�}��M�-g��+q�f2��X�X��^�t��f�E���㪷p&����w�pG6�ܾ�]���c�����p�S/ˡQ��w��z3���4�y���IR� �De��5HP���l�q�kIܼ����ڢ�~J#�\���x�D��F���O̹/x$�������a�'|�ݠT�(HÉ+7��,֥,u��f��񃻶G%��ś,�n�����
[���?��2�B���'����F��A�!Ik�0���f���nXշlȝ�J|�'ۿc�
�Fr�i"�]Zjk-�$z(����:�'��/�,M{N${�oG�/����7F��`Z�G -f#��o �C����)^�9��S�WXD__�I@n<WǸ<�*��7�k�.�wNS��/�722�PwD5U�-qy���!������.,+L�G1�/Y��2�hvd�Ucsw6us� q:���|��)q֯������ (W�.L]�mI|�~i���
s+�4�[�Y���R�P����4]�ȴwE
:��I��󰑄�9_��t�HG��>�6xHP�q|v��{���q]ޝ�̆��l��7�%�k�+?���.VV6ͤ���u��ӽ�177fVd���Ol[n�@2f�7���Ԃ�?"À������?�B�����+��oAQ.��?�o�Z�g8m�v��?�Ŕ���y�5�'��'-~-M�m�D36�aUЖe��K�s U�W؂��� ��*�o1�M�!�a�nx�H�p ��u��T���Z�:u%��$aE������Ac���Ӏ"?yJ�o[��-�X<�����䐖A���Jr� ] c2O�X~j=�xb1wdG>6(�̀泄�^���&�e2�� ��b���leV��`����qB�؍�.�A�4�@�?��g���w��V'uqy�<Q4^��47yzH�Q�x>X�j��6�x��8U]����A_dE+S��ը��2�/a��%�(�f�Y���᡿{%�E����(���D�o����y��<`��$F��	�ƜEgFli]��f��a�0c��I��o�f'v"�L��[��7i��M��ME�(�2�|����țp�t��XQ2|�����f�1�= M�_'��G�29�k�Zu��#�"�g=�pmE�^ڪ��b�'E�[�6���C�bF��U�Ts�����z,��ÿ�A׈�	B��lhwAwA��ǂ{�G)�N�u��gv��'I����<2��$�̭$�	y�)��������"3�����㙋^�3.!��R�pF��A%��I��Y��	-��@��hإ�7L�a15���T���� ��3���z�Ͷ��4��� 8�#&��C���֥�$�RW ~އ�rѬk̾��E�{��꘏>�=WpKZ*����4�T ����C�&,
f��8n�
4��z�I�����z��Ւp�;X��IYG�a\�.E��6�]`n'>��ߕ+V�e���Y�[�+��z�pKG�*��γ���m��=�2@ʽ	�>�].p2�DxŘV�{���N�8U���Ҷb��#߾��!i�����V�*���~��`����f6�Nש[����.�w��"�t��Զ-���f� �s ;P=a31`ͩ�w�c�|@R=����8�=��Ut���n��T�b��y3�N�-1~�����'e?����(J-�[���K��b�г���n�"/�w�V�3BW�Y<���������.Z�Z�o�к�`���7tp��Ƀ��w+��]̇�(�Q���fp"9���你Ij������\l��ܗB<�c�.��<��h����P�M�ha�.�X������ˡ4�IH;ar�06}Ŕ�D8�жʿm9�R�]��N�Ù �s�+����t��:�͗8̣��I�G��g�|��6|��`�F�D��Fo"�r�����O���.M��bR�ឤ�����1D�k�����k'��":�|�_ogZN�wo��N���F} ����0%�}���F�,�-0v�ڠ�h��Ky�\a�c����- �z[�7����"��<3�ڐ ����8���;����d���OK�ۏz����^X��\�Д�Υ%5����tS;"1��n��̷����3D����Uo�Q�9� �{��o<������1iO Q?<��md�._�z�0�^M�>�'C�~�,��u�׉O�ܦ�R^z�ŤP1~��\\����$6���n1(2�P��±��D�o߮�>\��^�ݳ*����A�;LV�PG�,ioK�'Z"`��.1Au��;��r�P�~���Q�Ƞ�;���N�$������?�:�sod�$+�U-��hV�^�(݋A�������І�p�2�iYU/e���B����U��u������\�>^!+ƥ�
�Y�e��&�h��E^��xmy)M5#f~�_g���Ұ��d��7����c���6aSo.��s���������o@�����Q����2E�lF���Un���L�M���z��t����0��V`Υ�4'W���[�i�qq����YO�/�u����dZ �g4F�F�Vw0���'���]��օ�Of:l1Y��#�^'$�9�9�h��b|��J��Y�K^�	�cT7���0��@����#�K'��:A]�đ���,�1x��������'�i�S}1�p���׆3��_�����4�5}@4X�� n���;�d��#�c.�z�났��k�2��a}��u��y�dy��ſ~`�)���������G�#x^}C�:�N6�y��x�^�5���r����So#��}E�7�?���	�G6	UM�ó���.��Ե�Ǚ~!�g�~�"왚ONޒ�
�$�iJ���Ř1�,�X�*#�vQH���	S1aE93���=M_�L�e/��%\�?���b���ķî�yQ�AJ˔Ȇ~1��b�Cw�8#Z�R�uA-U���� ~�)_�rKs��Os<�A՜�p����XB+^}55������p�*yç�D���yul;�tD՟�P�@51޳�$��[�H�j)���I����a#j;��C%�T8���z_�P[�=�z�ڟ[>�o�F�>�+�gů,^ӷ|%�|/c�=
�����/�Rd�����>���)����,�b̆��Bgl}��hb�i��ޗ�N!�ԬZU�ϖ�R<�Vg���
���&|���Y�r�=*���J�����!&d/Z��cߺ2�|@�,�u���#�j֑�q��	��?�OS��۷�_M�E��K���۴�ŷ˳F�I�|K��T��]d�bc��:�����f�k_x3�f��yI�� UGN~��j���8_�ӓb��
�y��Z�'�m�(�?^�⺏��u
�:�p�����D9]z!�pg�ϛO�/�ޣ&��>�J����>L��%������wҼ���"X"�3ؐurӥ_"��kbT�t�J������otCK�a�ېM� ���j��:�$�8��7 k�
����2��b�ҥ���y=LϾ�e�c�0��9`	E��h�J�Ȭ���ā�B"��y��r�^#Ҏǆkw��[�{����|���l���L'�0�(�Ӡ��!"���boD�ЪfŘ�!"�cf��t�v���	�J.���,��dc�:FE^�{�T� �'�ל&x�+agP�8#��}ϭS,Xj�q'KP;fl<~^������vp�ܼFW�{0�~g�l���ZT1��o7}7�1�ܓT\TVc����y��w!|���l�n�D�
,��f��RGj;�#��FA�{�>�����p��<��zeU%�Y�7���m�z�AO�V�W��0Z��,{���u�8;���Ym OR�풓]#)�)�3c��?y��ûF��m��g�P��a�dj�Y:B*�j�׵Q� �ۿ��I��/���'�O������!
������P��[�j�'J�oP5�����K�@V����(���IE�04l4�$�Vd���ޖ�L���-�����l�����F�����VU��uo+���(�%���}���ckҸɆ��KT\�7'i.�[�	�w���q��f�^�C��	_�k먈���G�Y�_}|�)cN1��+�6muM�[f�NxS�hT��=���O�UA��&`d1��Z�ih �D�3̰ߡ�8�zz��Rb"�8�`�2I�R��HnJ�glh��Q�[L�#۱3��m�ee�����G��3��0�\�EE�g�)遑)������FI��d ��+� �P;<��X���ջ	��_�I(��?��I������k,��Y�X�{�eݕ�Ft{��������}������mk=�Z�r��n�\�p��Z��>܆3i;�d�1?vA�Bb��G=$���4��b��Q�/�k�M�mݎ��HFw�rCb�_�?Z��}����WL�U��Cu�E��C�bz^n>q�qg@e��F�vu��j/o��7r%~Z�沪��f9��*�v�:���9@�bf5�磓8c������y���˱dhΗ����Iٓ�v��������$�9)�	�.筭ӥ����o��R��b�����
�0\NW�W�[R&�6�;ml~��.�޼7-J�������=���m��aE�1ղvԩ��x���T�v���`���H�D�9"��.�������S��mJ���x��	_o���ng���"m����/�\9\�SW3�&vA�wSZ��v9)�R�_��ڪ:�L��(#����.I\q%�iK�Kb�b�ǻ8T�)j#��������j���. �g��v1���ؐ�8f�t����$�i~��OL/ym��Z��K�4���:
��%s�XV
*G;���$�v��Fa����ol�|�+ %��s�X�'�{��G��N�XT��c�*�����Xm�k����YYfB����|sXB�ξ��N�����'�S�N�v��>9���AV�7@��P-��4��8�V��/k�F�=V�~Wog,�o�`����v�����j8A�j�T�u�4�� N!�8*�X5p�\��C�Kha�yM��R����)%k^pg�1a�5����ô�4r{u4{樳0�A�,�5$��28�d99S�L����݋������|���z�5s�#��'�S4�x���{��VO�V�t���k�4tj���y�k皉��/����R���������f�;x�}���f�	|_�:ml<�6����B&W{��L��T��l>&�}'��F����������B"ǔϡA�sdi�_�å��(����U߄�c|��0�9���* �w�ĸ��<j�"5�i��D���F2��tl���^�;fR�**�Ke��K�c������+ ������Q[)��c¢ �f<�k�n�F�H���QM�G�R��#5@l�|6�!=^���O����p��K5��r���O��R��j�l2����K�;s��>���5�i$���%��p�����m�E�˪��Vk�(��H]��o_�׮��J[���ou��W�Y��3#ɥ p��p3�������g�L\�9JqUФNh�XF9~�	���k���HF��R��U��R�S���8a!��Ŏ6�$��<��/�i;�\q��d�e�U���`�J#��8��*y(8���������N��Ș)���
�q��ۡ)Is�԰�8�F���kS�y�8D�}@	�}l�0|�C?S{%�LN��*ˑ�d��/4����?��bt������-��#ɨz���!�cbuP{To�i��v&�1���۸EE~F�U���l����	�
�SX��,0�*Zt Ώ�
Y���8��V�|=�8}]��Xf�@��։�].���C�����NU��<�{��l��-6	lª�F;L�ۥ^�Wk�>��;>x8�:��g�x��t�J�&s۽z�
��%��g�r�b��.�c����*2
�O����#��N�(܍ ��,`�JT�/���G��Ǎ��Fyk�Z<FW�O���V�yd�?l�K'�������T���$,q@\�����R�4=�p�jܱ�d�4����sq!c�����e3>h�������kY�?c�G˰V�	�O���z�E�����Q�aKM�ߪ�`q f�o�P��{���S�ҫ�Hk��mDI;a&7�(sS#O	ց�r��̌QZ�����I�\(��	�c{nTg���xO-���1�ή�v�vc۶٦�۶�c;m4N�ƶ�����N��y���=������9׸�kb�~�m�t\����C[ih�[+�[��'�>A�,�g/�l_Ni1�(%c5~�JI���%K�^ai�W�7�p�❠T��q�|tɾ�!�wu8��p�řq]�V���6��o�[��m�F��� �w��'e�[�i��Wzo1<ȯu�7�j�"�ߏˍ�:�嫠0��Wwu�m ��IY�-\�c�i:�)E�)�Sv�M��IY��C/��}lL!W��$�OU���a�HHGΫ�`	�\�9��q���b���v_ܝ��{Um�N+�b@i��p�f#_O+В�c��@�Z�����8����Q�&����]�7�܋��fK\w;�8 &O[��H�<*\�C���nn�!��VN��R�?g�����Y���eL�<*��ob��\T��LB�7�Z��!����pk������n>^����yP���O�'0
1a��:|CD�'��]���y���@�h7�d%c��$��dp��y� �|�ze���G{7u�f�֮��lu���5ql37ңoE;^���I�=���jݯ�67(2C������r'����x3�4s�5��4[�ӎt����`�M):��]_ҦVK����<����QSi;~����J�Đ\���}��8��Q��������:��m�"l����� [�)U}�T�	Vr�#�i�$�s�я�b{�v΃p��5�l�L��\9�2�J�{�D!���6��<W<�̿4(&�1��ݷ}�-�Z��C��Pw$�4�)d-51ϳ�噗�>]q�ڲ{����_��y�;��9������.�.ݵ8�a��f �\���bf����03�J+r�{�ȠCS'��ȫήK����ε�����[��6�rW�"�������`{��2�{��\6{�gfF#.�R��JJs����F�V�u�%���Y\x+���N���T��8C	{�>�a;��PM@�B��`���B&��~����y��L|�Wϕ�(����.}Ն�t1ϩ�~i8�g�,z��Q��u���41��O�!��\*����C�_e(��\��z�)u��N�.��L�vB���R�)4��}�X�&"l�ΰ#m��3ڵ����1��h���ŝh&�ZO(�n���y�g��	���x�6��8KרL9V�#��N���lϵ��ש[���Գ�nsÍ��N}��fb R ��o��ن�F�yz�F��ߏFS�����ʱ�[��"@d����Z]'�w��G���������n#PQ�a�4�ב���+)k�Xz�-m<�c�m�A�����K��Kcޫ��!2�RM�9`�Q�Q����𵽷u>����7W�:X_A�b�{Ao�OS0����f)�.�;��z�콋�{�#�8�O�����~��8���/w��[��>��)�5����v���MWKA���-SJ�����7�Ĕ:��f#��Uz��!�ڮ�$DD�]G�u�����(P�k����5c3lTkU�YG��Ն}��z���.b3Bi(��p���� e�;�O&���Ca�\�Q+ϼ*�/��NI5
)	9�J+���!+b3O����L�J��B�&�g��|�t1�V��)�(��wO;ʲ�g4YFӃWcx<�|G��9��b.���Ck�I�Ї�͓qe�mu�zީzΆ��m6���]j3���׻+~�f��M˥���	��9Y2�yD�"Uj���5&n�e\WQ�-�/�U��2jibF��)fN�T�a�q�}�J�'����Ԣݓ�8J18"���������u��/�����z�g1l!Q�'�����ƌ�����RqC�lZI���Jl{]F��n]k2��w#��z%oh�[����y��� ���ϙ���ݔ�i~��.�{��+i<e���a�����G���{J�\�Yb�1*�mm�7'��E5�ӊ!1B5O�5.a���)�yǖ.kO;;.V6�-�6�VO�����R�7�����h�P���^�/�[v�ZX�z���BԺ������']ov�8iX��#�ݜ9<���3'�Pl�	��S��X��C�\��B�i��CI"�M��t�����DP�][[f6���C�M� Ph!�2puv+~�ۿxu`�z���`Lf���%h	I
���R[�ڠ'�͓�Dg�E�Ԝ����o���E~Rb�+H�Y����S����;ث"
t��z���y��$�_�F=b*��x�|M�^��k�n�Z��qV����St����pp��XW��"����>/M`�p��ٴVt�pʁV�F�W�\6�����f�B��k��J��p�s
~R�	����.X(���ƕ�U�����!�zq��ݮ�B����Q����o;v��W�c/�M)��d�ˮHZ�c�ۭ̰�j��ҹ��c��iWCL�@�b�=jH�8�Ϟ.����%�{�\Sr�qjNI�����S�1����Tn3����S��'�)�v�"�)�c4�/�;�|S*�pb�]L*܌���u�R�	9D�\=�8t8=�ܟ���B����='.�w��8ZoU�H(�z�{_��������
z�߁��f�.����Y������&Iry(�y�b��;�����	�6�"Jڶ��l�Я��bP؉����fQJ��u�*mw:=���|-��H�jO����5���+�P�&b5�H-�oG���ٙ3�?�c��Yd�@��O�%C� �����p��zV�J���Gf�ԊB�8�T��Q<߇���**pA�n00�f�׵V^
��C��������.u.o�z�ݡ��?c5����E�<�>�c1��{ӽK�R24D��%犜��]4�<�����`�s�>�&��:N�v���J��1����Gs8@��ھ�(���B1����O��*��U���,�}W�(��s�����+C����N���R�.$#�~��U��O�&�!���3�7����������j��1ܔ^U�O��FCE���o��d��28�w[A�e�Y�����G'3�.���m��_߉�������{�xz�V��~�u-@"��2<���@��M��0��MS@�G'���؅9��� \���
|�Ez�� Kz�bR���n�ۮO����}bc/��M�Ȭx��$'GBt/~�q���W�BG���(�t]����89�G�T����3���Ɂ���-�'�^����P��_�A�dX�	���q�9PL��}�Q�Y_�W~)>�/N�R�.s��
��TS��N�q���F0�sv�l��s��Eֳ�b���b��#�É�۶�=3d���k�����t��(pi��s	���P�$H�*36ȸW\���;`7�VB�j�wo������[b��%[�!*G,�>�*�?e����]�6���e�4e�).� ���E�hj�0ݏ|�=�&�����_�G��8oj�\�Ai��֓M.$���}L�P����4)����&���bR���#���n���sZ�Q�������٤@�rv���H��Kl�ڸ�jT/�����U!n�{G�sa���_�����{�]�z������������W��� �;)�T�a�gS�fX35N���P���LـTX��ZP��C��x!�sUm�ik�l�4�l�xG�$-��mikT婽����T�qfҀI���>�&l�'�4�����-��"(��WիN��?.�Uqy]����[s"��5�E�L����J�N�b�g�Q�w[���=�
H����8K�fT��.��w|���69�Eι/'��t��21�v�����䏪B�W�o��Q�4�7C��a�ǉw;�����7R@t-E(
'��k�&�$��Z\1QW5E���c��R�8��� z�Ը�"A�RW��HI;�wJ�w8��=�H�Q��Ԓۦ۹�У��g��Xg�na����s����A��z{�o`�7�Lg���`�9���޺qt0S#=^���f'9u�;��u�p�i�}Zt7��;��>Q�D��/��T4+�g� ��}URf��㬽�:��H�&���j�5�A|�s����u&b�)�)*=u����	����v-��h���**݈�Q�k>[a?�;E
xM��FRpЛPYuQ������j�i/: ��0�M	�g#!�#q]�G�cIj�F�s�� 9.�v�^��7���
x�(Y�_K�8�2F���tQ��E�Ë2�v����L?�ᘤ��%���Y�����)K�����˽}.H��0�Dm�:�6�C��p�kUJ9*���m֐��C2��O�P�|����5�ti\�T��iQ��1K�h��C����2���펉�;��Z��פ-f�P{�<;�`�R���k~FMo2F%g\���~�@���}�������q��Z��'�c<Nç)�x�����h������V�̇�W"�8��I�J�����@�֫�c3#�]�l��h��az��1.u<-��__�\��o�y*�������Sgf��:Kʮ�+��/���'��6�ߌ��)�(v���Ǥ�n��''�����D,����EÇΐ�:/�Ff���(0����Kp���4��Vp�mޞ�Y�(���C�}����fp��A�gGD�W^c��6m:I{��~DJ�y�-�T]�MVL<L�����Yh�&�6�,�H���
е�k�}�n�j�mzҟ.PVuf�&3��ļ��`i�^�q{'��A�J��b��t��4�0�m��p���J�~4�Wl����p'*��WB��z��/���1�B�r��q4�"���Y������#i��A�x^K��[[OC�G=N�� �A�6����n����zY{���x�<�}��{#Γ�Gk�.�䫖��l'_�t��9��~Q�t��˄��ʞݣA��ɳ0��z��r	gޘ����c�0r^t��kR�
�?>G�� P{E�k���I����b�1O�g��N�@vw5����x��� !÷ι�A-�g8ԟ?�4Ugdg(>ߝ�؃��K�W	�:=�d"`����#V���q����-Gw�sB�����H��Ǧ��7b�w����пBA�Mx�X&�1�R}����}br��H���g!���{��e{�'�Cܲ��^b�F�� |�^>n&"\ގ}'��\?�1�����[�N5= )�����Ǧ��J��F�X�:�zܪ�W�1O�m�o�H�,�b��LP�k5��Z�=F��ݓ�IJ^��<X�R�����!�rC��t�-l�B2W��+�Ivd�p��a�lTM��$�}<>�X�<�G"R
�/���D�$���B��u��S\�]\-������遷?0{�:"�P/E8�\	L:���a��8�o�
c�3��T^L1"}�"믖��\r�V�GJ>v&>Ǥ��A��	��t���0
Dh�`�ƚ�<;���5��]�~�lLqu��F���@?��Ȁ�E�g.pi�8����l|�M	f?KG�����^M�/?9~{�� ��3�C?��w����m����	�ݝm�y�3C�{�8���m�-��͗�+��r���[�����N:��n�֗�;�C�u���Ք���@�^|���hB�Y�UV3�1��<=���S����3C����ދ�Z���5�J��4^�^�=G�	��f��0_�/xT�Ib���Q���h�}$$8'�0�A��T$0���I�0�n�f�!�ΐ�����#�ڳh#o;7s�)&�*&ı�!�;�>}�n��s���Nr(�Ts{�ȴi��>�e�'����(��|�Ɠ�!ǑD#�Q�'ڑ��Js>�i��AN�Z�h���V|�urVr��C(��O��o���F��}�e�����3�ö���3nq�}mݑ�F�#"}�UY���5="z�w�z|�ϴ���=��_Y��z���w�u���j�Ğ���M��}?�z���d���%"$��r��`�o�"�����o��Y�r�G�v��TF��lT�a��*c�,A��^����~�_���.�8��qj�����șh�zZ2���t��L�%g�4��mqZ��"QI{�y�J�1y{�>du�տ]�~���tO�a�
ZY�-�-o���S]�IXc���t�p	]�=��nK��_��^�C*��Q���qSK�|4���9�)by��a
��\߸ǖ�i�����~�P�4�O����$'%��	Ī�;��놊1�� ������\75� �#�����t�i��b/|��i_Ux��PʮDŦT�$�Hz����Ԥ;,_4������?��2_v���������v4��Q;��=mΫzV�b
W��!�����c��#�}���E��6al���>z��q�l�������S��7[4������\z�3�������^=���{�L|������&�b���C����ʩ%��Qh����\ᰆa�35���:̶��A�q��pk��F���1�Q$�,�j:�K���+n��X�.-�lu�D�=�j��FM�����[@��	�������Y1�_;�яR8E�8FVZ;_�4��F"�(��J�t�Wk,y��O�����*'qss��:6���Nn�fJ8l,�IdJ��O]�e���΁��s�bW)W }�K$a�՘�o�X �/9n>]�<�� ZP���l���z��=�,��6-��՘�����W6|�zC5�$د�ߑw��9:�q�@�]Ɖn�����R��g��G�F�"��o�����F�$q҂�P��*��w]a��؍_�~����Aq�J���o,f�	̒��_��*��~��k�+��ܖ��m�{2��ĩ�C2C^p�*"Xj~��XK��i_��(��|��C�VQH�;��
�W$�(�z'�?ǵ_�,>�lR�����q.$���Le(c���34T��>�%��@#�'+�;<����9fj�9�=�յ��Y�B�>ʡ�a�+��(���u-��'4-Q�:-k�K�ufWحw�Ǜ�!o���[��H���*�K�''f�:YNA'�j��&�d��+9;����(TY����~nD���M�l^<�~���gS�0�����-'쀪�X�a\�ˢ�j�/a�Z0��P�p4��uV;�T���U���8y#��)�e�����(*�j0��ˁ��d�9��p���@h���6�/��>�/��'�[��=$'����zMd�_z��VF[�w_�Eܿ3�8��O����?yO_N��8����8�_8ȶ�;]#.�6{J���^�z����9����mQ-���m�)������Z	��@,�i`�5K��������|�u��9%�hy-`jk��{]����3m�D��Aj��f���==�/4-�I�`��
�ͱ?��v�����>��q������f�'_��8���u����|����Qs�6a�\����'lq��8&�y��B�n0w�ay;Lb,�%ej��jy���}���|r�y�>O��e��HWw5Mbb}I�-��7���d�\�.����l�q~�"/~t�\Ѯ.Y����j��1٢�$�5�^M+�M5�,�ţ�$G��ܤ�=�9fH�sHc�?�����%8�7�y�&A5����`�C#�n�@�..�����$V�M���_��@͡�#��gw���Q)
��k�l��٘�S`�ʊ��-.xԂ��j���VeU���f��YyW\�S_ƹ��
�4�:�6n~E��w�����3�c�1h�?��VZ�-���y��}xc�_�4�>���l5�XPbY�{�w��^+�ùƻ{o�?x�o����؛���f���Y^�p}�{��&��H"nj�����Tċ?l��be`�I������D}����[��ET��uǐ�1� �)[6A���cT�Fa {�3�gs�:w�>.ex�d�]烒�4~�0��o8p�+�����8���c�/�7x?5m�X ~�˜2�10i�2t9�epi}r_9�x���c�������&���Y��Ӈ�T T���Aش��L���.4� LHF��w����蠢�����Xދ\�ϕ����+����㬱/���m-���hI@#r𢞞>��]�w<|�r����%�;��)~
�vM��at�r�ƀ};�^*�ls��YX���'(˓<̕��u$�����P�E8ٕ~gD�|�\�-���% ��m%���-�����gk�50H�K�Z�ρ��, ���z������#aȣ�������y�,9���m_;`�z�l�N� ϒ4�{���ڳz�ڟ,�!�M_q�w\�Y�?�e_�&4x���b��c�7x���=�)s��ёQ@�R-B?�K�DЏ�r� �\�*�PT:fLo��s��A�Vh�	�G]�{�ɱ`�0'�E�O�:�+˨�W"��X́��5%��簶bP�|y�����۷�a��Y� v ��#�'��+ݪ�ޔ��c��띹�q*F0��<��Tg����	gX�-ߊ3�>| Ӑ��N�tB�$[:ׅ!��8]�x���$�m$�[9�����q?x������� *�a-�k��kR���孕�GT�T�[A:�<M����P����{� �N�=��O�u7��W%�rT#L��x�$?G��LqX
-�%8Ih����G�`���&�9�&��y	�P	ft�2���б{\�C�Yo�pjh-�p|��߾i��s�N�5$�$'���w��=X�T���DҒ�<б,A�ո�k�*��U�T�}9�`�KI�]�q��3N�b��5���}��F����aD�v�����z@y#�:(�G�H,|���N�#9G�9}�d-�f֐�K�dP��!��>��O��� /1Cw"���iI�_��>Hv��SpEsà��I�l9��N�h�H����pR�t�S5pJ�	�S�nc�W0?I9[��� 6Dg�y�N���p��.�T��g��q@7�>������yj P +�̨y6�����?Sx3t�y��P�@W��,�F4��%0{��z�#��y���<A?��]{~(���Əű�Q��ѱD�ȱ(�ׁa�k������H�#�~l�>����T<�A.G��"]��e\A�i*:5�ɴ+�0��o�3�EI1#ao�ڞ��L"w�>Pxp�����p"�j�(�[O�	��6	#�e?
{?$�ۡd3"��cb�	����ǨN�%�}8�d�	�EsG����\��������\�E�� 	�E��¹�e.�b=��C8�aF����aL�b�w�n�x%���7C��
���'�s�4/�/�����'A�����g/JbՔ��v��h6D��A�:.y,��%����Bud�X'!�Ya��b%����A�*˞�ġ���A���;KO���?��`}�lS\�Y�{�Z���]�e!��i^U ���̬]��@� ��i�~xb��u�9�s���<�w�b�h�Vf�`h�-������a�}�I�0OD6���a��+�dG�r�E��NVr"[X{�᧴{.vyd�@/I����ԯ���蟵s��&��;��bu�O:)=���ݪw�ѿ�j�)�c:���f������?�f��r�����5w���O�B��o�TQ����g=����G9��C� ¶Q^�����~vb4�z`�4��H������2��-�0-��τ�D*d�����I�����p�$��!êL&�	���m�z|���a�T`��_���Qpk�d���ӗ�m���)0ޞ�4�6ͦ��#��J���!�<f�B ��:Wz��:b$�� f��I�"� ���aa��p�%�9�d{���g�4�F�
�C�s\r���D|T�&U1 �G��B�hu���׊���ĵEa����C��F�u��Y�EǗ�-ø�+A� _�k�7u�!�0�K���'{�f{ݧx� '��>c�}K��ӈ�1�xs^B��]����J�?&m&��i���M���I�X��X�Tn6~]�B�����m�dҀǘ�����Z�ղ�]�� N�￻ ܶO;����*mH8���EP!�YS�.t�ٴV���W��-7��L4E=*5S���;�;�tkM�&��
�ǷH@���C=Y_�a�V�]�*���s�ـ���g��3�S0��#(ܓ+��Tć����ﮝ_��v��2֣���2 ��X�2��F��@���>���>������M��>�_Z�,���{W��4YyO�R,O8�G	
�W�W���t��;�K���&���b`k����=i�ӎ(��.D�	��6����w��E�T���v˰V3m�6w7��J���E(pϱ���K8��_86˪3�o;����a���b
�n�����6�!�T����D2zy�r�f_=9FTD�2ڟ3�`~kUXZ;�����yG�M^ץ�;_��5�^�6C	8�l���v0X�����v/m=@]�=�[��o:�	��<Y��nV~����~Wm�@��&Kk&6�p�)�+,2A�Yljgi��QI�*�+>Z�yك�$%�e'�;�*au�M��5B�eľH%�����x�G����E�ȏ&��u��f �]���c���xb#��J�Q緓"[]�����O���~,J��p��d���K��T�
} ^�5��PO+br;��&����tFCa��p(s$��!*O4�x��=�~6����M��OF��ۑ�	=3��^Y�m �HB-q��IQ�ڦ ���/�|Xf��$�I�ط��0�(
7�G�;s�&1���s�,��57��+�D��~%�q�R���¯�Yפ����WGr-y�h8�Iw� YR �]���y4�φ�Ո��_�୔�,�&��L&|�d��\l�2s��������Q���c��{�ڹ��5-����﨟R������c��h{mھ���^J�>Ai��P��3�;է�>\Ѐ�{0tyF�t����D�Pk���JT��X�W:��'��L���,�&�KG����mF?�T��o�Y3�KF���G5ovO'��Y������h�Z��]d�3�q=qЂ�h|�����M�W[�������57�MB&����.�Z oW��P����B�o'��O�}��yC�-�TW&.�]�Q�=:��`��>�& FB��;�A9�W�/�A����G�Q�h��-Ǧ߬#�0^���W�f.����V����_�~��ܾ6��#Ӆ��!T�_�oπ��7�ʞ!����f��r��r�v��r�?ML����.���;㦴H�ȁZ�f��,�|#�ZJ~W&5��I]pX�]�8[��ɷv�W\[��0=��0@�M����K��j$��j��`�۽ǆ6�P���z�@ET~�PO�����j��L��lv�_�L���4����m�h��i2�Ca
���ڻC�+�;�`J�Ș�J��VP\�c����M���ٍ��͢�Sk�_H�~��$)�e��hX����*	�k��O*R�)}^@���L�1��p{�RPe�󝖫�_t�DaI�[�0I���f�l��>�GĚq
�5 
�|@x ��$<ՋJ���N0EǦn.o�W�?���;ܼ�� N��a��G��a9�2$c`�{�����k�nTv
c�?�Q��'x��Vr��㏘ݏœ�$�;Sb����qz�w�u��|����l�}�Y'��n"��۔h�	��
��1�)� �p"�d���*4�Qh8����W+uW��	�����ʸ<�?�R��v��d|��W�������\�ɯ�e�V��/�^o�zľ܆$�r�0'j�?�?����B���"����4n눔��Y�
S�~ۇ���4��1#��prj����Q��
�+�#8��E�!@�}�0�9~A,�ZCe�qf9u�폤C�����.G6�
���$9�!1���cFk��0�A�tq9B.��%n�
�`�h��.�wȲXT�e�K���P���zYs}��P�|�m�X���G��� _Y�z9@B��C���ж ��P�x�,&m���D!�R:R#�.��8�mʜ֍���()|+�Ge��='_�TD��W���%�n(V��\��ɫS�󬁷�DU�g���Q}n�\Y⩼���s�J��k`��6A�y�y&�j#�=��U�o�-%�$L�%u�t�M6����\�y�k�ao��C�����"o.���?��ߝhK�V�i�_>��V�0�4<9��=��d��@فi-L.� ~0^Q��T��+��PĐ�ܲ'�o��e,'�+���q�]mL��k����/o2k��hXna�ap(���v�L���Y+���Сz�RKkr�tť\&Vh������ӽC�4��S蹳�3� ��;�)��!J��W���z�[��9]�8� *�]�Z�r����QK=P����脆ٻn�C��ѯy�O90�o�,M$���[��)ѱP]H{�Z��U�����a�x3�_`(Bp�'�0����dx�oI�,E;�������? �X$��Y���c!��Wa��./2�-�Vz����js�sw7\�{F&
U�W��{C��۬aO��9�04��*�����o����.�W���4�/���������ý��` Kx�q�d�B9!eD9L{w'*���k���s @���'�V���O����u��������ؠ�h���X*�ϱ,�[���_d��Q e���'�O�/Z��+j���ω�?�B�3H8�T�m"aŎ>ϳA�H~Ԋ�gr��N�/ǡWnU�W�J�8���|;y#G�U	���������*k[�8��~=��
���]N^o�������u����i�GO(�z�0�N�BJ�|�����DV�qĩ����2�x�i���H����(Ht�h����6����y���Pơ�W xl�`��/�l9.�PI���Bs�����X*��?�4�\�!�ǩf��t��aȥ�D�+_�t�O�WY�h���ӕ��"�@�< �Ǌt���"ӳǎ{f�gX
��1�C� 㳛{�k��c�cҡ{��
��% &4�.G'Fl��hS�Qo�z�Mڡe����tYg�5�ߟ,�yr~_Ҟ�oa�����������.ӭ�T�h��R��9?	D_{}�#��f�O0�y4��Z��Yy�U~u6Ӏ�<�5{Oz���A+��]��4�CY�`u6`*Cъ$�4ASM�cS��r�~i&%D�#�������z.]��O��	����/6��n�9�δ�¹X�FȎ�����'�]kO��tH���{��S�dddD����$�j���k6o0�Na5xɔ������[�02L���!d�
+���  �刯[B�h�4���>5U�i}J-	�M���g��h��ԍ�p�!3��6��M!*Π�^h�5�:�g��O(n�{�&�PZ����2��,僩[h�^~@�!�ʪ��T��i�F޾ջ��0_Pּ7�x�.GoJ��&B�'0��S�'�Y=u��+������@��o�^�G������o������
{�a�d����w	���G�_ll�M߿4��u�-6�n�<�zmc�sA���Va��$���D�h)J��m���O�J6����IyY��q�"ڗw-!�)��#��>P/�ϙ*�R�tP��:�C���#���Lƅ�T:���U?<�?��)"��6לZ����p�0���π������Ǧ�}��d�[�?k��_!B3~�Z���A�����������ۡl���#!�<\j���3!��깄'�:|C�2�H�>I�p+d��n�7hz�E6J�a��>�n'�C��"h�T/Cy��RV���_���aښ]��
��Z�W���!ҔM���93
W��Q�#�D�v�iz���ZmC���s��7������{�~+b�Ĕ�,O��9!h���ݜ�]Ѭ��k��J� �Vw��'6��,Jo֓3��] ��oK�6�v�la��q�<6�NUVVv����M�gS,#����	�א�:�Kx�)"]}�ýE;W�z��:aǬ\9����v��ZW1��w/�J�6�ʚ�/+7���C-��^��D�%�%0��uPsd{����[�,�~����Q�v����f`�O�[��m���Lm(%ʩkLz�����<�\I}�K���*��yH2)K��^��6�-���s��o��������#u������k��k:���;�����0�N��v��RW��l�JJR47s��s�����:hQkJ��h�������2��67�$�0�$%$Y�L�/f\�Y�o��D���̱�>�QdW�A��]b̻5c�����D�,_ٳ��ԏ�;�W����ݜ�B��<���^�BP�[=\��?uP��~��Q�yC�]���t�E"ɘA�<(�@�cK,��X�\�V�̷)������I��%$��ԴֹpW5.�_L���;�-s夥(����gl���)ō3(�r��;i/���4��ZI�T��ŊVE�f�E� ��u�b��DDeb?x���qiǣ��^������R �XIÝ���i�V�x�C����c��-�x�O�D����w�z�n�PA�w=O\m��蠻*��M�̺���o�)��0���S�Mq�I6x�f�`uж��Dă�zD�N��X`d�hp7��%�M���@���xg��.sFnnAΐnO�L�#S�~�����x?*l�R3)�M�^���D�5���Ѯ{��2
�x� Y��=_������dt�����e�u��N�y
Sɴx� 	�# ��&�8v6���d��R���&�T��6���>�`+�V�9����d�c�؉��0�E��t����ͺ4�Wڌ<MeW�W��<���������q��w�M�G�m�_�6�v!Nw���m���Ck!���Qs&f�#*{���^�����"����*P�%7�:6�U�%�����3�ޑ�2!}���jS���p�A�@�`U�W���.�w������~����@�$���	]6�$��&0n�潘�O�����~��z�N
�Y��6��>��в�����n�V�!�������#�E�Y8�k�x��Njz.�����&#l����S;g6'BO�MC�$Y�ۇ^��5�t�c\-���{޾Z�5):�=���YTm]����(W۹�!�D�w��}���X/|��޲w���T%�$y�5��`�@$g��*x���$?T�W��$���$8���Wnq5�7d9��h(���
{p�J�p(��W��6�A\o�6�D6Xu%�#����Q ���օ_��w����9\v��ts�q���~����^kҦ���ima�����zV�vudR?�����o��2T����Zkw��t~�xd�&�{��Z��+h~A�[�[�+5�f1���z��m�cH�[�6�Xw?�
�Z��C���7|-A��Z-�QX$�O��Ԟ�o�87�p�a$���Pf�j��{�vP�s����K�kE�� &����9v&Oв�.��[��36�>�_�rMotb���/[�^o�������O�󷼗�K�}����s$����2l�D�܀����#=ڊ�?�/��i�-�������]�F^�F�҇�'���1%�Xa��g٦M,R�Ѓ�N��5j)>a���<�[@b�2 ��Hw����lO�}_�k5�1p_,⤢��e��{�?�+�7�W�@��v=o©�R��%���*��5����n�OZ7'UU��߾�e��o���i�5^�;-��6
K�~�W��r��+��ޤg`@�cܴ����[���JI�'�1:�\̐fZWm�aD��� ;h���n�>4�m��Ԯ)��m2s����:�6Z�
�3_�O)%Ж	?F��~ %ͩ��|���C�IEF��~�����H�6��c�*`�܎a�e�6쉐�*��h�Ud8Hh)l���O���L{¹�y���F2oJ%�x�r%��ђ���>�ǣ��>-�n1V$����� oہJ��r@�.����@R�LdL��-�W�E��'�:���}FVRV��i��QP@	��x��o\���o;��Z~~:P��A����3�L
%{�(���%(c�SB�Y��VI�[E��m�#1�-
��8�+ܷ�'���Ҝ͝fݮy�i _�>Ij�;�۷���ۗ�̀�s�+*���|*!�Pw;������)o�k��h�7|o1��L�.�DzvyDc��^�ӵ�
�OR����z݀�D��j�'�zMڠ�Ŋ�8�h�T�Ҋ�����@t�}bۛ��/���52����n!��OC?m�����$č� }AAye�k���vs�	�g�b֘4��$�����C�WEű �>��C.��I�;�O��'8	<��wwwwwx'o�{Ϲ_��k��]�vU1�#C-6��M�rW-���;�tf���� D�_C��7�ԯ[^F�G�����gkm��k�(�*���Q���zXM�1��₇&��`����/-p-�nU� 0 ��p�b`x�"O��.��d�=���x{	5���
��g��f�H̦��Ƀ��l�rJ4
����~�4�.b�HR�S=�P�2���Vs'�,_�R��&��N���av&����L��Cq�Xq9q:�]c��UA�oE�U�� ���ݙI�z���Ř�]c���ٺ�PPi����2�Ju�;��BT��/�wL��6��M�������ԻM2�'1���;b�&���6�8g� f-+#�dA�0]K��Í�Z��%��i�r��o��V�+�H:����EX =�������� BaB��a�H�z�Oh�8����1�WU�]�*�@��EC�;
9Y��$ _�D���6���h�e�,��N<Z�O�8�ÄM�M.�ϡ���[�e)0�_��_��4Y�@Ȑ��zQ��B���\��z
F��7u a�^��\��Q�����򟣃/h�؁��aDAQ|�o3?Pg���P������� ������ᖳ���v-��
F9&e���		���:��c̒�Sʚ��c9����	AZD�H�Hu$���,���y7�bͤ�ʌ��1�&P>���R��g.�V\��Z��F�Euv��9lg
��|�s�^k��O����[Ps|-�AH֚$X�5��b��7[��vXvh��5��6`2�#���%ۂ�𖾽�iy��3����l��I�+�������+��&�-��.��v�u*�l��?5yTi���R,�㬊�=5���r�l�Cש�Q�p.f��?H*��h��F��R\?JF���u/:��&��3W@"�q#�� 8Ӵ����ޖg��/gQF�	F�IS��+���M��ɭ>����Cӿq��7�o^�YQ���3�6�ļN���#:�4��n�~��ik�r��ҟ"� 0E�t(<���*�ǧ�,�v������q-�K��ڱH!�G@R�q�� �FWB����V��|>z�������v�P�b��坾���I$�ۘu���s"�m�bōn�\�� B�ft%��8Ө}�H~Zj���ײ{f����γ6z�S�}@�����BIzV�m� �=Ɇ�fi-�W8��w�6R�h�\���qjA�ɘ�\!�[|���X:�H`\�j���ȋ�튲wop*i��W1Lo��c�M��X�pU��9�|;\���������'>��<n�H�g>/Ҥ���x��Hfs�n��E�2r"�w���d��b9�����.�Em�艐�������#�M�@�}��m� �FO�*J�k)�1����Gvы>z��Fi��������Wa�O�<J�6lDCQ��;�ݕsH�鳸n_�3f	�x�E-����L���O,<X-��[��Z��Ne�o��jJ]Y��qav�[�	�<�wY `�"�����!ĕ�ҫ�i��*{8.@�J��^d%Ό�ַJ��hGB�z����W��t:⇍ ��8����Ƿ�K�H~�xO���FӳH%�`ߣ�A �}1���+K�{@��h5������qW��Yk?a�G����Y:�?߄F�y�0�z��g����̤U#�����""�?Lm�9��G �qjULK*���[����%oZK�ᖱK��tB���t�ΖjA���v;悔�\n4����˧B%%@��]�J����a����Mo1��`!WБ�7~I���{Q厷r�R�]�����nw�*����u*}�2�D�)�4G�L�KF��B����^�=3�)}��C�L�����룷���g;�_���؟anm�r��5~�2�Y%z;|_Ɯ:Z��z��uJ�)�����S��:8���<��A» ]D��z���:�E5J~h[��n���5��ת �8�K�pb	��ׁC  qT�ʍ�p�M>���̂���T�Uܡ��Y贜1O�e��!��n�h��"_�-����[M�"߮,R�:���	��<����܉0A���7��;���u7\=v�TK����yU~QU7������"�	�
��΄���SE�y4�����{��c&$SP㳹-w��xbB�����I�����b��ȗ,��cƧ���$��cVOwd�ò�
�l���I`�ČO��[V��hf�,1�W�v����-�l��5b��x7Fv�e#d��RA��/}/����e�����$�D�Bx�-��^+=C�;�3�Ш��������և�
Wc�$j���K��k �K� �T7�i��_I�N��2�f�1�> Ͽ��?閃wK���D��K,� V�ܜJ]�[���W�{#I����y�c���E�9�@��|�G�?m�CA�4$��Q0#g�WҐD��K_�r�C敕�/�����Q���a�>��sX�ϩ�/�:x�ZO�P�k)���c[���B�������=hv���Y��[��JG1*�R��~Y��X�:��[�#�|�_�y���\��`Z����Tf�$z�l�<ʭc��*O��>`�_��@�tw\�̥�M�I���m�T@�p�5��%��\lzH�SJ�&e���خ����Rp�/����x�g�)u��u�s�3pʟ/�O�94���2y��ޤ*���'��X|}��G���Cڿ{)�p��u��o����q�͹!:r;�ϐ��ة��\�B|t���b7挬u�v�1\A�+ʶ@<����`�l|��_�3�=.&{�?��g�CL��J�*�k��B
�(q�fw�:�P�C�׵R�Ak;�r����s61�B.R��XWٯ���@���u8oib�e$/qf93 �H큡����;�rvV����?pJ$BJMƁ�%������.��$���wC�E;���2�l�F�;g%�c�m�)���3S�N_^��
W-~�9A�_��=�v���+Rg��Þ��'<T��ܾ�C��c�1�r�!nJ&#��\�g�;���XE���9���1-�!�� C�sD���l��7�mJ���z���1�A�CN�!� ���b#%�71��H�:�-Ws�UKkv�zx�NG��HgA;P��#P��m$s�Ԧz6t� �"����D�G�b�e��6��wS�'�W��d/�>�}:뜅�.��������@"�5�6�5����T#���W��\��5c�����(�� V��Z~IJ�<�O: �y�B a��k����J�$93�OY���l��w�f�u��d4���r���o�/!�.i�A�04��3�7�QA"Х�'�G+��$������L%�a�g:��ʴ�n��x�ڠ# !� �P�-[`�u%�0u������
'p�̀���b������{݀-nA�Ƨ����u��f�<�q�D@m�>X��ى��K�3��Dd0�3��:XXnڿ,���6�'�a��z�p�8m|�o�c��`��j*jEJ��������[��'�q��.��LU~�wFU��Q	�$��I
N���0��i���|pl��ެvD&��|���ҫ{�4?�x��ߊ(��� B��T�7��9�����K�}n~�ݗ���˝��/�]�V\���p����|3k��I�E.��}��Z�l�b�Xw ���HIK"K��z۰h`btsoY��򷇝&d�����t�G=���q�)�VU��,�$���������/���vK���MV[[���8��D������S{*�bklh?�o�F�|kp��wx֞��tFn����Z�p��Df ��|��Ch�j�d��x��t��PC,�Y��,��cs�%����c44��X)�+���������$�'N�`M;K��2���x֍�gAQe	��tW�u�*Dׅ��i����'a�kfUym_bE|ԓ0��ez�q�4'�d0��а9N�s:�mu����a���x}�6E�#� ̶�F�Lď��ٮ��.-�U��T�:�|�$���E��U��#53@=(S����%Yj=��"gZ��x��V��/�:�%�T��]�5a�X��+�Z�۝+N�R�~ˣ�o���IZ���c����>Z�y�v>��r�n�@BW
�@f�mٝB+��y��Q	Nu,+�2)�И���I���[�y�̘1���# �����?7��C�җ�9��Ak�Z��)�q~?W��7�!H�	��f⚈�I����IC�)��1d�9�>:lFB���dԊ���dA�>�6rJ�~��A�T�w|��2T*oTÑϤbsL+ ���]c
$��}*(���cb�ⴻ4�VJ��^����&��h����D�ͶӮ�6���� ��MF�+�J�.�VH^9L��|<7�s���V�Z�����0�|,4_M4?
��^7�aI�o��I�P.�2�L�I���w�r�gh`�\+����)��g�'"�0�7��:���cyH�T�|��B ℩����uCyQ�7%[{eT��N�v���������tk�V?�xj�S��o�O��zz#��q�X�� ���mJ��1g�$�+�Y	���I��Vn[��^n�^���uNJ���G�ȱ�����#	�ß��ß��΅W�T�ׂ�b�Y�}n��W{�_B���e�C��ϖiHM��5):'=!D��-�#$�h	�8��k4c� ;����x#C��6`IUE h���瘏�E)Hs���~�����&�K3�{���Kܭ�� ��_	��,����V�n��#?���I���& �j���x1��1ߎq%Yr� T�k~#���V�?�PR�����V���-��.F#�cs�����`Fy����������9�H���� ��Z[O��>h�����D%��UeCM�R�`���e�Y����v�x�7&����Z%ȥ7�ܩ�̫&8���H�oi���3��ߵ��]І�3g�Y(f_Ǝ��.r�d���L��ԟ�JK+�>pp���Ĺf���i�R����-�HW�×���W�ש����=��-;߲�JRS�� �!��Yw��$�6O�N�N�9`� ����S����G��_i%�%���M���M�\�/�_����X��<6����f_�ROupǑf�z���@�9)X�vU��e�˱��1X��))�;Q\�0����6\�EH�b���y�|#E+�h��"�$^��W�15��'/�x����ՠ@T�O��M�@Ŭz�RX��aa���!��t��:�J�XWtn��2w�v7E#�K�Ed�;C=f3b���]�e���;L�=:{t����v�n�����Fv��H�y�k7��&X�?�hG�D���a����z�y]�D�t��Q�Ă��Қ	����j5���π��+�� ��r;��ЉR�u����4p����a�l.캰��g��߆øy�����`t�r�!�U9�9ON��Xۥ(������-���ZƟP9Y\�=��J$��VVv�$��q����1�Q��v�IZ�HA��n����?ɫ�v�.��-3<��ph���_�Y�\�T:��;�jX/NyyiX/��W��k^G'.}X8�gllU+��ët	��a&2ds���>[5��s��������H�REM�y~�M*F�s%d
��e��j>w����aTz�D�q�T���*����O����.=��.���l���H�<�ޢo����᷃ò��~?f��� oZ��U��mG"�u�L�4f�� �w��a���f���0�"�!�bc	1�P�� ]�̛��ޢ>H�Hh�T�!@��~M;u،ZTR}���ǓS��w�l���vI����5�4%��������:�P��?�Ԑ��b��7ɺu�k��Ԣm �z �Mi^C��:���u81`[�}�+�B
R��đ�*������o�igP(�&;�Z\^�~%����=�v�ҷj4���m�"�U�\�`B�[�էZj��X�NO����"��*�U%���x#IMaY�;Ib&Vq�����>.G�<>�.����t��X��au��?���m9W��i�Oƽ�*<=�=�k�����U�u*
8�abK���t�M�+�P��ئ�gEĽ�ǻSe���b83�Xuvlj�4a�:�&ֶ�:��F%�5����<<�"�������m� Zj�lNf>��$�=�\E�{�����P������X��0�k"$WH7��EW�	��A:�Y�-W9�R��D%h a����܅IL��N��ȁj_��E�HBY!�nL�O�������lB$�։�Q�k�T/b��pu���ۿxPq�����$����K�<]MNO[�}�E����'�6�>G��|��x1qV1���L���k5v���B���qړ�.٣>�C�wD��64b�*&��t���^ ���|�E�׭�����n|��!*/a��$�׵�)'^����8�%^�dWex����=p#-��-���Z�W��ZbMk]F�ߋ�m�'@I���c���^�T�L��|kUHg��p�>_�`��M��r1�"7MG�׀�;( h�	П*v9ktY�gV,�ę��9���6�A��>Dρ���*���rҰ�C[�&$E�khIyp�!V�O�"v�RgS�ÔA��BMV���(J? T;\�qv,�ϑqF�ތ\�Ș/�7D��&+*t�W���\QC�K���ǣ���|'�瘶�d�SB�h��Cy ����>����5,0�Ač�2�ޭA 9U�>��\du�_�z�m�`�6_g�n����!	��y���ѓ6~	\�lM:-zȍ��3��..��Qmz6+���s��YQ������5ǹ�{����
s]���c��E�۞�b��0�����0�~�g� ���|rQk⑓�:Zy;��^$s~ӡv�\t��%�Y���M�.5�&����{CwV�x�;^�~�I-����Wt,}ٺY��~`�:l��j��PH���Sj�GXr{�;�JAå~�pTY��~�&&�w@Kq!@a�3�b��\����<�ZE+̛\�w�G��T��>��w�.��� ���ZG=��t[�!���)ܠ�-9��CVN��?8�vj0X)n��Q�*%U��#�=-}	��}#Ty)\�j��!\��4�����<�p�V1��f�p�Y1����/R��u����`]��)r.b�w�'�ޥ�-�t�#91`3��d�����".��W|�i�l�����S f�v�(f �~�
T��Q���H% ���p�e���YJkMp��S�$_�Ѳ�O��S�E	`�{[O�>�^eA�G��x�iC.UR,N��Y�V�g9�)6�[����hM2J�|��N�$-�گ�Mn^� 5�Q9�Jaȧ)|8m��kf���nw=�<+���3��uW�=!�|ѭ���l~g�Ծ;'�}v�S�-@��1�f����j��O{���ƙ���{7��23X�|�WZ4K#��C���+*$_(l��ɲ+=��x��G�l�
S֯P�uP��Z@'�.xt��kj'0�W��N�Y\��O�� ��4�up1�66�8�H�L8�k��a����yI��9s (	ʧ ��q�j�BZ �0?��$<�z#%k ���X ��~�Z�igt#����y qjG����y ��Hi%(N1/-7��UF=rC��3��e/�~�+Pfq��CSyk��R
n!� ᐶ�ODGzDG���.oڹ�|3uы��H�,�Ȕ�"��6kC���E,zھ���R {�I@ֱ���=�h~�U(��q��B��P�IYUR��RJD��4S2�
�͇�27�c&�<q��5��(�r�_0ѽ�]�< ��d�!7�~w!�Y�v��^i�h��r�5���Ky���|+r'�Q���_y���ԛRN�����l�Q�R'�:@t�ZQb����?ݝ��Iz��{��!��̩~�YQ�'��`�!p2-\w���t��A�b��Cd~���e\�ufw� @h�E�����hX,[�60z�-����[��s����p���Y-��vS�&��T�'���M�����8l 8@J��� �h�����>�x6��!V?u�౞�WR:�5�Li)�I�!�N��"���s[��H&?&T�!��/W�6�u�"-u"�.#�4�D�B�����p���IJ>�pe�&8���ji�zVi�3ghB
�۞=B�z)�o�=��s��1
?��(tn~�P��lzͳvP)'S��wvN�p� e9 ��q�7��̹aΨ�bM��?`|�z�N� }����a=�Z(�����\�ە���?%_�1	���J�?�^�>�r�6�o.S������\}X&G�uk�΢�k��֠�v�˺�0�?M�XV���U�c�B�C�ʁ��[��g�Ӓ_x���Q���zS!��|��t�0�.KJ7�a���W/U��9�]�SO7ǋč�Ѳ]�K�1���g�����U?�.���bW�Fgɂ@��ӧ��0�=�2�x%�b+�/uY�l�w��q1���PnnH *oo�U�cw�ꦘH/��"K0�r�~p�	m��>�Nh-�T=�T������B~��*cR�?�~�������Wʙ�)��U�����#�nD�I��j�'b�w]��\c0��C丘�Ʉ��(/74M����&�{��Z�|�w@�6�\���
���<z�v�}FϚoc%��E�w�ް<���X�����t�2�>\�$�n�����9�>��fv�|�Y������)���Q�e���39��U�ܼ�4��f�,��r���.%T�)�"&2ڧ�v�8���qg��4l�Y'��-f��zv�s�X	���O��"�� x"����O���{c@%ރE ��+�砓;!%H:9N��_��o��KA�(Tד��#@���+���no�� �� �\r��(*���ǈatEY x	�Tc�L����=1 ~�����[}q���|W礷�^��W��	��k���w!������A��*2����&�7jgWq���ӋJ�{���у�P=�͠Fp&�|ǝ��ȟ�V�w�2��;%CFHy-�N)�,k��(�7�>\����j��(��䓞~�+��e�=�aӇ�ڞz��֯��ܒӤ���r��+r���[BvO�Q*�85v1)s�M�G7/�)�K��֖_�ߔ��ˁ&�iیT~9,�w�.ⱸƌ�E�/�U�m�Q�!����g��XF���|�������K��E�����B[����Z�O2�n@W���(Nѝ.Q�ڑ� ׽G�RL�s�Վ��~ϐ�f 
Ё�ip�K/K�Y�&-�P�C\���u�n!dGX�sɐN�4�7�`w7�aC-�gx�v�f���J� �"*/���^L��?#���{"f%�� �^��@��������;rt�n}*�=�4O�����nv��@�id�S���,�樖��BkM	t����F���ؐGVt:�ru@�ު������W�SBE����������i��S�I��^��˧�x���-w�#'�]������DdE�c}�^����_�H��M/�z�S;ǆ�zz��Ȩ��y�u�������c��4�oro}]tX���P^��] (�*r�,�������9�y�MY����㺿())�Z���ї:W�2��bP�|%��(��m�5+ӏђ�"qY���)������􎔜�c��O�����m�C���Y����*K���Ob;V�`���1O���W;�����@=2��H���b�g�����W6�`���M���r1T�Cӫ������O�:�a��/QX�#A��$�9pR�M�;*�� �*�`��>���`�Ulע�MJ�g�9
�@\N��3>$j3U3i3�����2�8�i/f����o������U�#��Q&����]��_c�[cRJ��bu����G.z{�NN��r��y��u;��LJ�bF����X�W�=[���F�5�.�;Lʝ�\mͰk*P����cY,��5!��D���z-<z�����������B���}��Z�b��s���S޷�Dq���ťWa?^>��:-����=X����	6�&��"~4�5W�ŀȴ��XY�~ M/�D4�d�|e�BM�uP$��u�ir�Ԍ�r�+�M��J=�{q�I}k`��:`+�\��]�rR%��8g��N���S�"�<�I�2S�����/x1�(v�28T�a3���� �_����'u�ҖlY���}g�H�o�������V�LJ��B��g>gtSG�a�7�K�BOZ	HB�Ul&���p	=�!&�`�㹚~jJ]����H|,@��S)��NpNE`�dE5ճ�w>�۬�5�-����� �&"I\7����A%"�Gؓ���j��|��U��அ�z���8\	�M�O��B��Y�@bvC������vx�N?�qtI7���B��S����D�P����J�뙇�2�ym��;
��#��Ĕ�M�yj�T�6�o�WӲIe���A���b`8Z-�"i�����*jPГ��P~ܿ��ā���}UWyP15�s)ZUz�P�%��>��ƻ�0���F��mu���8����Ec���?�@aAPC��ۦ�[���}֏����Z*����X���S���Ć^�F-�U1�k9�W��]�A�C��o�����6CR@߂�2��z�h��K�mJ��>�KNT�597�Q�8�.�2NQ�ҍ:_��\�]�|�ʸ1pL��$:�"�\��J:Y��z�j5�##��%���z�3�ǉH�,N�j�	���J�|,���\h���ؚ5�Х)C-Z�Y����~vW�[�&.���]S�܍2��z�Y ��A߼6���=d��c>w�R�Y���?�54�73@;ʿ��`\�8*|�|�^S���h [
��˶CgHM����wd�K;��'ٜ��na�������I����\�@M���ba�e�D�(io����|�۷DU������PE�������c�sZ|�->���XT���Ӷ�^	����ff����6�T쒌���*q��b�����0� ��oD�󨄟1��Q5Cwë�}��[M��5-�a�3���������z�������P*O��_1��WmAH\�I�{�ꂈ�[��_Q��d}�:��/feƨ�*��=���]e�*{����b'@�ȋ��;���5p�9�?����H�& ��&���wE����6U�i���{�f����ۢ��i�OO	����H8 �b5������"���0�}7����W����W��k˚����K��������@��钁�n^�V��������L,�BiF,�R��4v��;�O�C�>�Z��K.�&�]�#>D~��"l3��~������
�k�6pmv-/V������-�����#�'ݵ�#tE���.%���x���h:f�zK�Y��$WYr[*1�i�C���5l�6�@}IԐ@̸,�W�/� A�ك�8 ��i���j��T�]/�萕P�0L�.cF�M7'�����}�X�V;�S��kϳ�*��Gg
�x�Rb/{���E�>��[[��z�I]%�_\K��:��)�i��^�[Z�X���}�)R���1��bS榍�ԩ-{��7�>���V�#C��$I�gZC$�x��gMԍ5���z_���k��>��Y���3"}�qR�e�x���/�߈��Y��>��Qk��G���>��vZ�P��Z��l.-\$k��Z�����^��'�e� B�q���()�.�֒�´8���RY�S�yh�k��n��}�_�z��O�q�fSI��4$E�H�A^g���`R�7Z�w�߉��t�����b����ޤ1����]8�nh8�{��y�^��&~ �GR8��`�D�XLUW��m��cAr���,�%��$����e�	R ��G���� �y����,&ɗ�E���6���pj�+8�i��� ��"@#Z0g<�f�|� ���SHc���P��ˮ����`6	HCI�@ݻ��x���d��-�l��V��|��1N�lwy��.f{��݌�&����ө.�.z~c/ڲX=�3ɴ�k�P,}�Vϲ���M���/R��w�9�~u+�TM�١3�9�UG���y�/���5/�S�L�}z��~G9�i���OBHBի�}ʣ���`�i3�}Dkm����nb�ja��'�ʦx��$
�$��h^Jg��a����s�EpV��w������Ũ�L�n��5$A�����W���C,�R�ʥ��1�,=�I�=|#����Q���b͙��o�\>`E��J��o���֧�y�j�ԧ��#�ӞF��|[p�r�3�ܳRwD�I)t�u���1h��t�7s�L�g��߇s C'[}��C�2�,��z�������h.I�ߐ�K�uB�yr��k��pT�����4��H�ba���:cT�b3_Y.+��Ōpk~�i�e{E^y�QП��O3��Y��Q��/���+�X3�j˪!��n� 8��L������*yFm�I�T��=�KQ�~�7.����bc�0���� ���}�1d��+�0<�9F�_F��z��rӭ��������Q�S�?�儶i�7o���7J晓Z�Y �LU����79��|bN;C�B�-TU^l`�H�[�N�a�N��l�) d��@}��u�� ��z�_�T��ތ�]���e$>�M	hM�'NC3�V�CԐ�)���~�|@DG� (���j������m\�ͪ�DMV�|��`��t�K��TD�6�	��Qn�)R.��Nk}��/1z�$���~�sX�����PJ�K���.䗡R}1��1���������A7�@߁��
�w=|)ܖ�mT>W�W���4�oI�h$����N� hK��H	��+���%>O�ѐ�ۑ���O�"���ɟ��a��*�_�G=��Tq�'-(8bpC���i�Fu6[��n����Qrp��� ����ؠ=�M׼Da��"��!�8��w�ގ;���F/������i���&�P"�N��R��(ߝ�a��7��}�/D}V�~.��d�aH`$-;l������m>7G�M#�Q*���d�?�m�Sm�GꔪXG޿T(�!����i�'��p8�FQ����u%����aO���m���Vc�f�O�X@������7��t�ZTv��[O|���c19�}qJr
Ӑ���=I�)�
gð@���Dqc�i�U9PhN̕�,�9<I������5R�x��Xn�c���XV�&����*�V2�J�^�'oY�O@W �n��6����n+T���_�z�g�-h5�k��\��-�:@ߣ׼$CI*B�7k8WU�vH�pW�YgEDřj����n���ؐ�e�M�'^a�"��rY�Z0��z�-:��y�
� ��Mi��b`UY�S�S�1>;��"+��rc.��(��_>S��'�7F!d3}&%&h۹�~��5�!�X={��>�M�>��
�_fN�w�sԸF{�.M��2-&��V��A�V��f���-�N��(�#w*���֎�^LT�n�h��^����^mQ�`����&����ҁ��c��~"��;Ue���,)��Y~ڄ�`7~��zW��b��|��叞v޲VQ�t�Ď���%��� 8��h���NjkI.1���h�%��~���x<]��P�r�4�ab�Pf}+C>��q^�INny�p��x+z��Ҟ*�������w��Vk��y���xfvS� `��e��]��F�s�Zl�N�(P� !k`�^ � �A`2<�RWFrz{W�w�$Kz��D�rWU��R�>�8��&�!���ۜ�!���p?N�*�.i�XZv=��!xo��oI�T}96Ej(騉�Q��˾{���rXN���hq�M�~��֑h��Z�[q������}#?�q��lE��[ۭ�+}�L;���!����e��7�EzgF��]E��`�Y�h癦ʏ/�[}{gh�
�����MA.�	�8����V
Š���2���l��!8��vd�h��_�!y�[!W�,�����ƌ������p��~C!�W��*�����-��V�S< � .tn:V�<}��~J�f�/�ym&�|sl���(�ó�BP+E����&XĐBA�G��s��Iŝ���o��Vd��:dH�8�{����V9澺�
dm�1k���(�ws�1�[z2�֜Dp r��ݾs��R4:a
�Q�)�7����T��8q�b����{�l��*�x���{k��<�ʇ[aG8�#��-�ڦՀ�N���P�W5#/d;I@����0��q���cF�lP����xJ��)��񶛸~<Ԡ��:����,(^��\��ͻ�'xۖ���ˁH�R���ܭ��g۱�[6@���1&�Z��̥�Z4~;�dũ�d�F� ��Ť�X&�Eh	���-͜r�W�9�m�-�Z_!��q���A��9v��`�@яխ����>-T;pC`p���{B��P�Ȳ��q��)�p�Fq�QC>&Z��X��H�_óIТ<ڸ��^[��tN\55�Y�D�@��K`;D�f>�I�D�$�� A$$�'��&#�'��<��C�~���4�������|f;֜l�! ���@͠�� 9��	9�Ujq �xMpv�RZt����U�_BE�����~;I�^Y���X�+��]	=`?p�X�O��E8��~�F�R�p���WՆ(���~�z���(��ƳP�Ed�8�e�Ax>���K��=�VH�M��{���B�"����M������]�L�]�<��fb�v8�ףӖ�)γ��� v5$���΋N}N�^��V�O�j�)ݲV��Ϫ]T�,5�gxKű1&(m�q~�Q0������"p�C��J�c4�Q��K���ũ�� �bO��գ���k���vH�6�FZ����Bi$h���L{�e�~����[U�����}u�8�$�P����s��S0(��g���	�i
�
����,D@��P�p��k�I���L�mB�%4Q�������7u��f�g�g��o��S��Y|�ea��
�P5k3PB�f�.0_=]�&��Ğo��	�ܦ�z�y���f�=�ȣ��'�[/�.�v)��^´��mw�vM��@����N�C��3�O��nea�WYe�mkL V�#e��S�!�����Kg}u����:"j�VF�-:|���7Q �*�=8���4<9��nX=g�:�������$$ *����Vd���gk�%�S:iI��=߿�k��۰��5~7�C>����=E�RV��{�����u��t�%�%�P�t�-�vL���y�h�e�ʲ�t�"S�� �tAbE8t���Iq�^^�2���er�әʊֳ`ve��a�`�e.8�%�b~�=��-ڷӇ�D7KA`�v\��������Y��B�i�(tF�8�{�xGv�S�q(�w��ߚ74BI�%B(.�0�	&�H�%�'E9�.�D;��C39-��;bCDjoaV�3X��]�h[�C�&��n'&�Ŧ�z-��m�}��$�x�W���~���$t��!�Lop������W^�V`L�*p4J!�}��
ct@<}:F�F6�Ҩ� �,�~ ��#��-�æ�"��ǷNF$�"�|�&x](��m�MRK���Is"�,�q�ﭼv��v˻�[z2(�ʞ|>�Ҝ�1�.n �_��˵��w����	���	��t�VI{@=!p���\R���M�mxSg��͏?[?��0��(6J�;?U�pB������E7r�~*`��ܲ���v�����w����N��W��o��{ٷ:~�^;���v��� �U����\p�׈Y՘˒��ы�Sч��Wr�G�{��S����s��h��4Ƞ�i�##�ob��D�k%�$�3w�s�.�z`��ӈt�wf�xa>Hѐ�k��aw-���#"s��'3[�G���8�
�ؘFI3����"�#��æc�:�_j`[�����{rb���_��lo��&��z�������MtRk;é�Po@�c��x��������S����6���(�$`�,>*u���a�tf��\������Nn��$kR���Z��퍒�w�x!�;�+/*w�A�Ȏ�uɹi?�+���u�wg�Z��u?��e�ݿ[�FsH�z��h��>�@r��~������H��c��$v#�Y�$��P�]�!�7D��{�.xшt�}�Y�d�?zYt�S�-qu	��Ug�eۮ�:�NiP��.A���q����A:�!���F�������߻��?�����y�ו3{��l��#g,@��.�R9��z��FߦW���V�'�瞙S|��@�xD�����9d�'V���f-	�b�]\[�7�)<,�Ѝ�')��L�O�0ཏ88�2�RF1/^�<�`kS��/�~�r����+�0�;�`�;��,�W���s�,�_�T��9��]�|&�՞k��=��lg�(Ǜb�Q+|��?�;9�+��$Ɯ���3�	wu��nH{t�]t������B���ȨO5��,o��,&�Wo?O�R ^�,?�,樂�A�T1����(u`��%��c������"�C���֤p���c�k��;�sip$���K�� ��8��iM.� �+���>�}~����TC�����C�B�=?�&P��!�5��yl<!���ʕ������Ƽ�c1���⬯��2_I�KЊmbQ=�6Ƴ�Sk��$x����vE	�<�����)ldܢР�w��qF���e�2S�)G;�6~5�q�P|�M<Q*,���6��U͹����J�c�6tٳͻ���y�;/h�g�u� �8��H�'�٥#�K���ǒ�^|K��k���%Z��W��&GW�jY����R%��@�2��*o� ��o1��U��9l�^�z	�:m�үW]�9���%�̜������1��0�*�ѢY��[x�#�J�pQ~t��/6Q��~�e�>l�^�9+e����z�zfQ(��ҒZ�������dP����c��&�%�#���PpW�A��h@���v5��ƀ6s[��a�R������F{�����}w�-L?,ػ���T��;bڥd@+�$>�f�y�ά�H�ƜHm1��Y�p�~�L��0��C
+���t�D�q�U��p�x�����D8X�d`��G�^VaJ�J0��/��9��:��W���>f�_խ�=VPT�j߫�
��/�~�U�����T�)�^�Z��8�����8� 9�`xk���<m"�����]�甜���ߖ�n8�r%cc����/c�३8���/�����w(E�RO�MWЮ=xY��� �r0�$8U���?�����pv�@��� ,ʇ��|O�C���4��$��=|�{n�֡��n�SҍEmIff
�C�e���̓�P����Խ��Jw%�1��д����P��d{>Q�IZ:���#�5Ь��_|N:C�\���s�vf�I`຅��Qv�ڬ�c��L������Ǳ� ���E���Du�Q)%�d��ߝ[�~�����T=J�;��h��%��{QV��LB�1no�zR��)84u�+޺d3��q͓S	*��1q�V)<F��ٔ��ƭ ��x8G�*W�g�vft\�+$W{lX���&�����c� �˨�p". � ��7��FMt�d��:���:���=ߛ�3�®X������y4+����s��ޒ���g�"Ro��F�s����(�{,2��/�i�D�o�Ƕ�����j.�/.����@�:��h�i�.�Q�li�!�8��~�];l�&��O��������AA��e�#��o�I���������H��$3��9mp�|�>�BDع����b��j�v�L�g[���2��s��-0c�����|�C����[o��ԇ��9����(F�	�x,�傉V/�� �8y��coQ�D����xx:��UEe��/1o�[��Pu���1N�x=*�������˅܊J��*�hѷ����ECI�(�6�����֯j
�Uv���F���ݜy�(=�y1H���V�6��J������e�X�#b-�ͩO��}�d���G��,V���^�}�1x�|��kBe�tNr͋�s�G��VZm'�#`�@�v��4�~�+P��ۍ������("w�dS�Hӣ?��C�|���B�_[Y�4ut�!�2�~�C��w{E3��{����4����ά�?�O�ߟδ`�pv��AlOA\N�XV7g���e=�'v���P�=��Iy+�Y��{�\S��\~L�B=��&G��]��F�鋅��0Sg�}l~1�^\����p�S��/�L8��1H��D�w{�����Ā�[d�0�"b��
!���7��e�Qnz1M�m`r�'���>Q�2�� .q>�un����*�%
�� �-�Z(��_��0g��4���O~f��$.�ʒF2�s�P�Us�$T'��HC�J�M��5�4�8,h;��#$�,�v�h�#���x�z�7{���<�z�> ���w���}(x�����r�`c=��uS��ѫ�yu�%|�w�}�H)�{ۀ��O��f0�j���6��p1�m�0���� p�;��ySim�Ë
s)�J�6�e,T�l�*�k�.�%N;KN�}˼������)���f]����k�q	 �*C�P�ZO��,j;|�Ti��wrL�#>wp�W�%��"�K^w�ݡQ8$^�&�����/����M��$�������%����~�;9�(x�~9���G_�W=�>SԀ�[&��f�cy���JU���A�z#7)Z��ek�6$#4�#���^
�{p��i�]�Y�E{��	����*�h-~F:1(3j}�xY��r����<Ua��'��΂$Z�Aq�Q��T�g�H	�������7�
�u��pA�����h�x}r��*�nB�v���ˈ*������9��ZZ;|d����gl���$x�|�p��Ȫ�nPT����5�s�D�I�r$������^5�lQ�+��}�@��w+P3��M[��D�Iɡ�A&�x�D�X��(v�e@�<L���vRNt��_jw�5�[K��O�Q[tޗ?�����Ψ�:��+�����qΟ�-�o}[��
��0�Y�.���Dz��6����Er�n��@�}�����wÂ��:��lڨ�-�v;�$ן��'�L���m	|��|��@��Z�V�#�%_�i������V����bT����7��;��e���K	2E+>��b�߼0`N%z�z\��ӣ|c-��F��'��o�%ÓOi��Qj�� I�H-ek��.��-�l���w�zgsh��}�;k&E��`��|lJ��tⷘ}Pj<���_�.��5������;Ƈk�L�.t�<��U��7B�����C	
�{o�\�@Do]i�ʳ��Mκ���2��5���(��;Z�:�V��o��G�C��b_���p4��ߍ�R�ː���zK=e_9� Jڧ%��(�e����C���9�6[p)y8�<��-uAQ3si�5��
mإ�C=l����D�M�D�<��\�����A��c.[A/i��'���lв�3'YK��g�T�Ԃ{#w��؞�+R�-a\m�C�q��t��
��t%��co� �5��OQ-D	�u��R�d�o�WK�1�1�È��8�
��`5-:ϯ@��o�"��
^����X��6MW��yq{w��X}1�Kц05Ar��b҂O�����p|�p��vH��n�ۥR��]��\�u�[�ْ�~�Jt��t����>>�q�u���
#a#&�J�E9ɉZ����5F3^��?�ݥŁ�!}|��e����x���,�W��x=M��$l�����Q�A�gY{��5%3Ֆ��L`���_��J~����u��ʶ��~K��tsJ�պi�������G��8Q�s��g����HAi�4�ᖸ��|��wuF��9�(�n]�D�z�cZ��6�W�N+|�.A��H֏�?Ƹ�v"C���2e7)�x� ���+&i�jօ����]/�8��E_�+�Jr��)^��x�M6GO� �f}���v>�h&|�����
}���*��i3=��#�Yޠ-�vX=I�]��ƛ���:�{�-:��-ѡ�k�]��hlGg�/vj�ۻ�B�75͈Jĉ���Ҷ��tۮTTU�<���F^O�K��"����h��&�F8_
��]�<�zy�����o�l/4���E��ӵo���ϳ4��QSڐD��V�#M�����և�y/km�_�1�UzpW]<�E�k�W��M�z,vU�?YhP1[c:�2��hn�6�C��ѱ�\EW3A!.�h��ؘ�θ`�MӍ´��_kq[(��_E6��2UD�b#p�xc݅0�^���e�"f�{�2z�3�c�R�&6ID�K����@�a�T�@?/>=�!��q#��d����7۸ѳ*uU�N���̛{l�m�|��%�˕�զ����G�3�1�,s�}��q611�F��)�Vs�����נ�~�.V9b"P�w����<�7`�n��4@�8S�G����T{t���ٟ����5Z_�[��#=�B�b4lŚ���kR��d`)jf-����n	��Q��+g��9q}��w�
�`T�]�w?��2�Е��Z`��3��&jld�l	X��������l��u�e�2�ubBh�d��:�x?w���{�ʢ
�~�����]>Ћj����,֯�;o.����{���)�w_�#��U)��3/�.o��TC���cTѹ���.�ܛ4N�kU|�1Gp�L�F�Q�3ϾL�݃�|]��_�#�:u�q�h� v�C)�m��`�*���\N�$X,��,_����ш�yO�͚��e��Ԑ�s�M��o�b4B�.�D��f}�����1Ƅ��&)�nKA��vw�C�j]�GWl�
���)wf�	_���<)�ޥ�W-�|�F7�����d>���u��d��=n�?N�Φ���p�sځ����� :q�����������/���<�W�p岧k5�#aj�Ȝ6`�a6��&�|-� � vw$@b���nw�A!l�7�y�G !I<'�9��.S���Ro�{�YV|�_�Q�I�D⑏w��&�W�0(���v���0�ٸ�d�:.t��I{U�ʗpe�,�#ŀv��t ̜�I�R��/c7����S���^��Y��s����m�V��X��:[g���k��>�v���:��V���X��A���2�2�w�=MJ���s�m�*���/�nd�@$%���Kl-88�CZn�����y��Jľ��hz,�K����೒?PGaΙ�м����yg7�tދ8D8�u}�'͂w��=��x)Ji�pC���i!5%��`(�B����P�|O�Q�G4�;Gc{�k"u���%Z��XX1��=���qo:��Z}`~V�.��T���N����Z�s�.Z��ӟ���l	�(Tot�^�N��S�`�kŞN�R�vDZ:����f�0'�j8ُ�.}D���l�X��I&�w?�j�O^~��FڞB� 9�>�Vc�]X�`�K�2�W��Sl5$/����.n~qJ��!�&J!.�?����y̅Z�����"�~>H���a��������T�����0b�'�f��~1/��S���qu������B%���+�*�Tk��Θޅ��6LK/|����#���`V?����K�1릅X��g/O�Q�,�q�5�4��ǌQ&����j8Dx���G�B��[�����)%��k��d�L��	�>��Ds�ܥ`[V��Om���<0oB�7���SG�m��!w	k���q���Y�N:����l�،�_��?��d�}��S#h}��xFn�M�=�b�ۊ�e�tR���)�t*����� �3�7@?��gp�����f!mW����v���/.�\d#��0g]F��� ��_<���G��i�fq*Ƭ:��捖��!�b����`�S,�k+)�9E���Щ0:o�C�Cl�2��/�_47��|��Qn^�[3v���xVi9�h]�6��(!	���ݕ�I:���q������	�"�N(|G�?5o� tb���Bj�@�A]�����v@u���9s��Y����U������L���ܽ�a5�����?tb ��zm� ��=4��+�(�ӨXM�q��?-�G��|�mCJ=�7��*kKJJ2�>Z$	�G�� �*wS<�ˊ�p�1��Ն/���3|8��
Iٰ�^3��)o�E�����hH�6N��-��肬]CO�z�0���ʰxN�'>nz�8<����]MQ�6A��㣯L�'�?����fB;Z�*�%6�! ,2���(�լ��vc�Q[��?�6���s�-�Zv�a3�rCz�g�D͟k��r2���t"�XȾ��b��^�R������d�2IƱ���jr3�}��R�&/%��O�4bc��Zo�"b�%�+^�}^�%B�t0R�R�J >����3AF��G.K��q��w��0A{T�J-\�T�mx������ے��k�ٍ���c�����E�tP	��������1���'��rç��')�c�P��%��2�G��!���Z:�A�B�W���f�h��G+��9�B}�"��x�����bN�FC;�{e�-;Q{��dB���IQ>�dW�D�<�8*�=^2Fr�f�#�j�ɭ�~i�1��> �J
iʖ �X�ʯ�DbQ_���@aQV�I��:R�7�bI����nf]����C8����ʫ���r3F"`0/<<P8{�_�}��"K�|QgP��4A�'��ϲ�|�:Y�<�p�r�b��~�k���T��78H`��t���p�rc�;�`B����5ύ̹3�V�<M���e�I��˵ژ��sN&Q��E�k�.����9�e�dq˳%����?/Ȋ�<����>m��{��p)UJ�����8{&�X���5�zf����;)P�f�s25��`�����>�=)�S�\�J@�큽��BKS��쭎�%D�)�k�GO~�.�+��Q~��2ٻ{nhU��r�^�9^(��T�o�z���۴�/Ù��A���?���4��x}>�}�'Ũ� ����&,(� ��k^����� vMVP����f��d6��H�����Z���W�n8!ҡQw\�	����Oq(��PY�Fw0Wc�H�1|h�լ�,խ��.��FA��/f.(�N�q6���M��s�B��b�7�eu�$~s��ko�4�o�m���B�m-�j����id3���(����*~<�Y%��^<33�Z{!���z.o���3<2%%�E�D�Vga|5GLlѹрd�n��B�����n|a�U�~tQq�x���˷��M���,�+к�H4l�X��ث|9��$��_����8��W��� ��͉#�g}-N�!E��aQ�T6�#�����0l�%�%h��T,~�T�Ex��rw�D����hx�$]�>$�%��=�_� e��75�Ǯx�xl��fʨQ�����Il6-�^����և�y:X�\��Tw�Ĝ=_,���Q�I��h��;�˨�j9�+��voE��#�\��HK�0���Jp,��S��g�o�`�ኺ�����.��N��[~��6
TȔ<�E`�9b����0�r 9dM!aB��p����[����KM�j朗�1`������*�y�fB�ƬTb��l`�K� ��l}�찝���*&��%#Tq;Yf4U�ކ٨^�/�!�v�n�gZ���#Ղ�И y潌~G��B��C�4�Z��?��x�X� ��8�ԯ�_jl:~�zy�B�4�L��r1�s�z62��_��6Ͽ�y2B_�L� �p�5�����X�xZE8,�w%��>	���6�[P"�#)�4M�c����}Hc[���pv�L�+m׆&��`3�mʖ�D��|⊷�knn��J���ڴIw��e�eӠ+�&b:�rUJ=^����^��,��n�_/�ю�8�F��߇O�ӂ�c�ԅ��GIL&1���ݹ6�k�p/ܨ�f��HmX��-r�������F����Պ��`���M�n+��F@��Aa�ůg1{(��m��P�����O]�g4�pH!�R|��4�+�h4��y[��U�Y�Oչ�3`���.�/rQ��p*Y}���sԾ�Z�~�<N"Y��:?��w]��<e�1j�C�_�����	�I�ޠ�h\��g� �R�Y�1
�/4 2BuU����"��)�����#I��)����4e��}>e�h��ɡ���w�H��V�8���.a:����/(�� ���ӏG8 ���/�����;Γԥ�>4�b|���+2��9��0�!A}l�_X���W�v�I��Y�z�l9�U�%��I�Ji�Aޚ ͝fp-�_�L^�0$�d���+$�\����bv.�Ԋ�8v�8���w}kIq1�\6Zc���(��<�g�H	<#�����k``]gx�Tn��ω%�s54O(g;��0m��b�ܐ���f��oީ4�w��3YS���
��Dw,�a��#
#�et^&�#�R��)�-.�:N�חvg7����&�k��ܖBY��aM���.��m���]��أ�+�ڷ��-U(2��7C�V�:v3�Y��:U�S]D�ׇ�G�!da�`��̣��9#q�΃r���ۜ7pjw>���3�HC���6/�X��_V��J���^�;i1�ŉ���72��H�E?��/��;�\=G#�^ɪ	���:�ƾ�e��*��A�����q�?|ې���O�&����':S��T6M��E⨘C�/�J)�:�}-�ZR贴m���mKH5E8�T���PCX�z^2w�̈ ::��r��fb��X�"B���4�~;=�y$E8���F�$�_t�'�3�Z���	��sߙ>8��l�@�<4K�A�Y��6͙ld+Q��W�7d�,�+��{��j�Z��!��4�@0W}ץ�t�J<�DB�.c��Zn�����!k�:��9���0c���q(��H��� (D;{��hw���"��`�55�����|UiŅ�6?��&g`�5vIv�� -��_<�O'K���3�d�N*� �w^�ʣ[���U>�.���}0_�D�`�
�����å��ϰ��L������5~d�f̕���'�K�4[�����F�J��2z�٭�˹��,0@�*�X��ࡪ������
�����f��w�0I|��^������Jv`��@_�x�0���'�aF�Gӈ�9F�M�"���j5[����]}�}�+�tCw���h�d"b�W��j�����'�"m�i�G&3��=*�Q��"�s�z���{��"q\�~�CU�1�s���@e�Ԭ�U灩ϬM��0��>���U�wΏ|L���]7���绌&�R�<&��P��-=��^�Č\�'@6L9M6���L���%w�Y2w�4�c�G91a.5Jʈ�~2��Q�R)}AB3��r� �N ��I_��,�m��sWJ���)����w-c6?N2�K�XEG��I��)���������"meZ��`v�0s��/M�]�~J���"Ӈ�[��м��Ĺ18�	?���^�s8\��3�XZ��^"L;���O����<v~�O}���ۦ���� ��uE'?���)���t�7؛��� k�My�~���o6Mt�,�mD�cM�Dݼ ��<�Fu"�ى����AĊȗ�SZ6�v��ʸ�#ܹ6u���4MI��� ���|ΩTk��4i�XD>P�Siں����cKz,�E� E���oOa������6A,��tQ���79�����@��ݲp��4�����&�j�r:U|�C�Ƙ_�&/����; �Y���|��l=J˺��]�n��°v-�H�}�C���&���o6;�C����Q:}G4���ḇ�vO���ُ��x)�Uz���������h�'�7�]2�̵�,q�?����/��ǍO�EH�`���q5�dW?ջ�#�cb��%>z����[C8Wm/ҟq
�6 �lK5-%�8Bl�<��Dj{g��Ux��?��Oi*�!�k�J�E<r�ޛ�'�S
�����;iT]A�4K̎����Ќ�a�a�?�~�����7l�<�F<-����X�(A�o<�h�������E�m[���Y�&#	z>�e7�Gm�ѽ-�m��ӷ��X���d{`l��j�!Qe�Ր���8��go����訮�N���un���넜��Q��%Q M���N�9Nlg�.����l�ߺ.���� �J�-3���Q".ƥV8\�l���d�Y���4��q7�ZG�u2�k:�v�����h3ފ��Rh��������s5��&I��r��.������g¯��[.���@_�+��wNL���@�3�E�E��}G4R�>qe��(�̪.K=r������C�6��f����$ڌ[�?�{_Ů�u��������:��-l����$���^�K��{�!nA���<��<sg-��AA,�ύ��ي4 ��|���$��d#2�߄\��d!���C-Й4�D�D�=`#��J�͇!��-��nHN��:N�o�]%'�k���?4
��e%kT��A�gb'�]�:{{7״��� (���r�5ø���H�̍�:���]J�>Wz��<O��pS�u��Qsp�da�~<
̬��=��e���E�~��}��c�8An�i�%'L#��"��I� �Ⱦ�s�O!��\����6M@iǓ�	�Y���^A�Z?b=�S���y���K��}}�I�A,�nu�<!�춲^`]�]�BL��ӌV;�f[��z��z���>���v�7-�� �
dޔ�K���<���9�gea�Y�W��vo/0�����D��R�/lϝ�tsFQM¦��!P�[=���;�چ�Z�^%�uԕhU��2{��Վ�������h�R�)�+ͼG�}��S�e��K�7p���R�eY��>+�_k��=�����~c��拐��v�I���&�F1�h���H��!k���r��H;ٷ]�j��5W������ >�a��4�[��D[�P�E�Jr�5f�Cr�>�(6Pڊ1(d�i��~�2$�k��*dZ���hI|�/��,{ɫ���R�p�kz:�.Z^(^��pf�9�h�:Ju.7ۆ0DxV50�Cb��%D�Zպpv����H���{ާ�W"zr�3ה����p�uk=��ޜ��M��x��=.u�k+��k[+i���}�sb� }գJ��A�\+�uI�8�?[R�k�F;�o������]�ݷ�B�'���j��
��+��w���bs�R�o�6�$s��r1��9��F��Ҕ\��HA�֒]�/��8T3E�#%^�A��Ժ�ѹ�t�)�WBh���ױLW�#��d�E|�lֳ�f�C蕯�s�����L�� 93�+�j�+��������E5RH�/�ԷC%��5#��C���S$�W�.��91(�m+l�M�'�c߰�r�w��[���N/_����J�� ?$���M����aQ�en�ൽ(ɦ�O�4o�1?��}�� 6����Zbs�*v�9E�]C�މr�%���7��wխ5�P�Z�R�Սm����sK���ˑ#�	�X�+�N�����/͓ƽ@�z9�=��::j%��H$��S�����B�$矏K5i����Γ�}�{���W��~�8�
~uP�+��0a���c�R����v�O�(i��G�ye�C�*r*{�M�XH�cE�Q�3J���A ���)�7�$�����IkC=~�h%�_<h�VW����r|�9����R.l0�'�&Xs�	�3E%`1$a�K��ﻝ���!���(���ц�f�A�9�k3M���GW�Ȕ�'�<5�$���-� 0�h�`^F�~�%Ŝó0� k	�������x�����έ>x��2�u���>�L �O��PGk%!�@�n
��"�p�B�Dy�:!^tښ��M���6s釔�����ߚ^��c��[����Y̯MA ��9
r�p�-Ƕ�dۖ7���aL�L��G �b�csEđ]�*,j�\��'�:al�K����΋M��7�c�5���L@@��vJ�Z�]����8�SwD�]v4�ķ8f8�7ێ���K,�;8�m36�hn%M�{.O[�;��Z7W�w��\\&t���Q��b�>U.KVl���)�,d�g����7ug�s�&��O��.���Y�����@�e��ۥ�at&�L+
���v�2 9�: ��?(<���MoW���y�l�v�;è�sAz�K,:�!��A���Wn�Qsr��S��Nl�x��^�C
����Y="@����7ϗ%��v��"���u��Sma���j�O�:�$��1��`F���-�ҋ��C:�V���,�P�e�v�����m;@HZ�)�Ŗ�^m�?�I^-,[��Ÿn�_�?���u���)����zk�`Z���e[KW����L��X��w��Q��:�t��ݪϢDG1ૺ9>�[�MY����@į�11�p���Nc�Հ%	ʝ.���E*��NhĂ����ڕ������N�mJyQ�h,�?�<&,[%���.�a��瓿�U�^�Uy�Q0�s3z��Hd�k�u8u�c��8S+�F��ߘ��%��Ս|�^�ő�\��jL:�n��_�������x��0
s�ͳ�,��e�\���baoHD�CKo�F�0.�<Qf�b�V��3Bh�K}��q-�HJ�)Q:1�yW#uw�l����+d-����
�4�05�&��p�Sebm��Q75���EFL*i�lQŮDxYk+bq��B��K�X@E��_rxEb	yW ��E�TG/��{����z����XKԻ#�b$�k@);O�qز��b��ё���ۅF+��4�xa0(��VH�^�M���:f�Ǖ(Xy9u��<��j켥�:�d�����=���8�b���Ȉ�w1������UH*9����Xy��!b�l����,���^��9��K��wm�(8�X�'dP���Հ��쳃��pK��kY��6����R���R�a咾�_!��3E?��T�Ź4�b�����ʥD���͔��faſ��8��#�=R��0�^����~$;^��°ќ�k�Epd�Z�qM��x���������r�$�\�n+���[���⇦�1��Ve�:����|ݹH٢�G�<&c;h�`T�'���v���N$���R~��
-}V��O;�(�3ώ�]i��i@5��Ň��g��v���3S?@�M+�r~h����ǡ�L��џt�F��3/���[���'R�B���|K�YE$�t�on]�y�Y��iנb���u�Mvk=1@L��2wWoVu"�!�]>�����MF��Yr�z��x�m�3a�n�m����FBݤ7Š������pC�V����� L�SC���d_�1�b��>�P(PB��>\�ϖ��,6_�B28-��$^�'Ŀn��6������w��:2+�]��� �E�h��<��,��3�9}N�������l���<�����䑬L�i�8yCW��{��@T�`Ȳ�A�s^�#��-,7�J��9�&}(��)���#74� �	7)��o��d��{��ŧl��E{ݝ�0�Q]�L�&�����-�"Q����Y�w��҈�P�� u������#|��K���n�c?$��_X�u�f��^�~�s�;�nř5S�m�ըk�z��c`ק�mθ���.�Ĉ�s&\�j)���s�W�\3��x��-��ZH(�'
ը�H�n��q9~^�3�3nt��c@����=����2DYmp'�p�V��7�d1|�w�B�/K�U�j�yG��S�c�,�X��$�����+�t����:Q�_2&���M�ŉ��y��Z+⹭��������ީ׬��d��V�R��ǦyPEi#EZT�Ns�V</�IZ������(���ڮ�ּ��ҽ��G:�>��w&d/���H���E�-��fxw<L��w;'`=�UR�R��"�u47Y2�������V	���C��xA��>����B�}���1M�����@�c�e�@�X���A��.N.�\6�,FjT���&�\"��)��}Ǟð�5ֈ���k��%,��S�w@��Zݦ�N���c�k6��fEo����3/�c3#�X���.����~'^E�=�9�:�F .W�h?!���å /Z��#��S'�c��$ʘZ�)�%Q�-J�>�zJ%�Z�Qu��1
�ބ�;pdS��5SϓìI1�mVrsl�x�MkS�b��1:|g���/q�z%�.�u��K8�-��ɀ�c�Xi�,���/����%k��r����읜�Z>o�%UGj����}��Qx�aɵ��8��T������!���6���R�9�J�?P���ܧ�oӬ��U�u�\N�,�!�`Kj(��(yP���Ν�n�S�H���@�M��%��1�'ƽl����؊3�]¯v`5��c;(D,�0~�
����>\L�����*<���Y:�C�s�oY��)�a��lnZ�.��RO��;&��?L<�w��l,��Dݶ:���`ku�[Ԏ~�I�s-��7���R�GO��>2�_��G�a�B�J&2}t#Lɮ��b�
<^�V��M�l{gW���I�n3�3��*4�uF�Lc7D���K6`�*4]�5�PR�M9δ��ܰ�3�i��t�}{W�/s�
��64H:�ڇ�J���>ޔN*�H�����y&9?�Q����9�Zb�%K6e ����Fb36��Z5W�����݈Cd�G�PV�g�A���m���y���O�`�_���@�ר��,��^�6`:
6m�Rʝ���r�zr!P�h>�-6�"|b�m����}��7�D�L��P��oj`��^@p��:1�Fp�-FMm9����]-��vɹ���͑��(!-OM.|#�!|Y�T�T���n��:X�S�Y�ϔ�1��o�]��|*�H'���iM�w��]X�=c��J:��
4�[2��O3z�TgT��Y�;��|/U.	}QB��_�E=@ca��S]�q��Y�Ye�_�l&~�N����+#�:���_�>n��h�:`;-��	U�r���奧�~��c���M�kC�$��wo�"�������(�t�	-��ߠ��U���*Gc�O����1��������Fm��iw����_����{��G��e����ot�_�Q"(x��5fT��8[݁ըF��(0�ro��vة()	�ަ�g��O�!8�Ħ@Ӭ�������aѩ�b��/uՠR���٨������~�o��/�f���]�.N���5�7�� �.�z �LT5
�J��Ԓm�,�77O`;�-H�*�kf��9�o.dv}B'���r̥����M��TG	y��x_:i1Gu�(�_^�ݯN���>�����||��Q��ԏX�4g��Rw�}��x�A��y-G q�8Y�y9<4hD����5'v�|�f���P�=�急��r*��[飳��/�:��}3�[��lߕ�l5�]+��i�O�q��m�j%|��GJ��9PK� ������?RtM���}wLx4��˞�6/���JX��ZUŭ��`�t0������TX��D��p1�uRB�T)�`�ŷ�t�׻;�32����G�M�8Fp��ּ<0gە�#"^4
�tt4BY�S�e8I hۙx'X���@�P�{�6� =���h��f�&\��د�>�ԜCZ6I'�U���,�Dw���2���ʒNs�B�b�z�j�'��C̬��C�4B��1�ڧ�pV��o�p*�S
q&��%WѦ8�~(K�׬��VC�V��Y �B�,���Î��:�zĥSz��^�o7��*�E8��n���lT"/]^��ުB7�n�����=c1��_��l['�s���_d4�[�r徒|���*Lr�����<|�+��7S�F��ɇMCK���l�羋jI^��ҽ��wx�wp�~��9�b�x	A��'T���f���ۉn1��{[���,�@����P�tz�M�t�m,�QKBU4����`}�(���a��Xn9��5='��Gc�.+W�KQ)��b8	�t�8�16�q��´�?27��7��8NȨ6�����
����h:zԀ}�����uԽ�����XS���/������2!��5؟��Fd~�����wM���~���p �C�v��>���a���L����+cB"*N-��������W���7�K��ᮏ���|k��MW�eeט>ܢÖ�UݍX�k�^V׍�3b�;}��P���'CI�����6F �p��[%q�/�w;��M�O!�#�Z`��
'����aі�F���{O	,�C����^I���r���s���\�f裬���ǐ`����y"z^�0��f(X�#2..�#W���$����b�2X�z8ؕ������~�#���w	���!	A�ww!��		������d �-��6����n�U�?��/�U]���{��=���w���$j*�˂A����97�m����a�n0V�`j �M�T��p��N�ц_��䤭�Ղ�y�\��c\��SY�K����m���WE_2\Q��ˑLVu�/���@�������_�!si���ʆ\�ZcN����dYT ��9�f���k�!�9@�N����|�س�97�"�yi�5�i��l	Ȕ�dR��m��t�Z����P>zt��x�&�r}\��c��&T�ws��d=�EvI3��R�MA��iΘ�����­�.**�e�*/���=*�ٗ2 ,Ӯ�7xP��~j��߫&yib����&$����}O:��i�Z7��7Z2�9���;�?��ěxJojm]�^c�b�B0�,=e�ڻ��М9^�T��s���8PG��~tK
��o!S�n��EFgш�Ȑ^��+��A��2�@�H|�Y.�E�;�+��JK��~�����+�(��͟��b�{��,G����}"��:���tt��+Y�B�H�G��e�)Jt*���qn��XښO�P��6c�g�i|k��������&6�o���8e�"���'IV�Fi����]����K8���I�,p��Q��?��'w�����fI�����a��|���$a�w��@Y>W���6��4��&Y�E��x8T��G����U8/Q���y�:�W�_�B/���!�o���q�u�w����?��ֻ屔��o�.��,�IpR!G��
�7@���6I���ט 7�<��-��0k�7�r$�ͩ+�̷��~`p&,��m�������ς1ɍ#Z�u��)h����!��E66�����
�k�z�5�ۣ���Z�xTcD��<b���V��ǳ9A�_��������QpT���9+v��H�I�I���2�,M�v��w�Mbg��KA�{"0Np�I?X�v����l�V'�6��DF@��_6�[H��ȿ��L��[��I����*{XR�F+d��k���0p���[�����h�8��b����oPG�����������!s"H���η�T(Uc8o(�ղ���&vR���O6^�$iÒKA�C�]6�۶\}|)�ylg͢�WJdg&��՟����+�V�iV"�S�Vz�o����������+�^Mr�b���Ǯ�a� �ʙ�E�f�Ԯ��|�a��p����签��D�4DM|K�kF��#���	�E9+��tB�`�F���LerC#���q�}��R�<��A��#��](]r6��5��3l��B���~3D(Z�GVI8y��!�:�'Y`j��?^C����p�0r����5	���Q���g��U��o��(T��Ӧu��2�S�������U���ުz������ӣD�
1�B?�69�L-��$K=��N��E��&��u��6zlK(����|g���ܰ�ʬ�6���7��s���3AfC]�}n��k�n��!�L�����Dxk��4��-�=�7G�Xg=��f6���jn@M��i��h�ٺR�ϭ����>�'mh��gy��A��^�?;� h�=׹N�~f��"��}�9?����v�'���Zn����=F��v�O�T�E����a����lʌ�n����i���b@�b� n�ΟM�1ƫ��������曅HId7�|�k���S�]?�r��Y��q�4�'��h��Z*��>mW�Ò������b!G�����q=��%�K�Ѭ^�$�̈4\�6�W�~#�ݖM"�ӜH��DR�(3-=1b��ȶ�_l���ؿ���oco2j�&��p!�c%?�gG���y��ɭ٠�e7>�te�X�V���=3�/lBn�x=cݬz���rާ���T���q�ο���i����ףw6�`48^�TE��]����'�_�㓽>��'A���@��a�~`��c�-u�C2^���뛺d/��D�,�{��1�!��[c�^I�Nɀ)�x/*2�`�B~��Zζ33K�)��+�G�O=�˄��~�*�'8%yż�c�g�t�x/���\sS��ޅ���>�T"A�Sh��t�Ӟrx*��@�&�1b�G���v��1q|�zߑ:=ڣd��\~����m���W��2��HJ>�'�/v�*:���UN���E�Rׇz����wF���ՎI��
�-�GC# ;hW-QUl��ؾ���
�9";��	�p�}���ia��?:����5�i'�<��[
#>��SL���n���^1���,�w^@#��~t,��xg�������/�2�ΰ��4�p�xub�ǿ� `�/��2�]tX��=��D�y�`8�����-#￭�2Lw�9g���7�Bw#6���n�n��؏ �P�P>��e���YP�r�qc�jT(3nRI� i�^���EVZZ{���.s�Ǔ����ao�7B�7?�bx1��Y�E��;�v�+�J�O�C������F��e�=��"�	"��Ϣ��7"�b,��k��|<��5&s���+��wƈ5�O|rg�O����=�;?ǲ5O�?�f�'>�/��/�;�#�ej�;�o�Z��X��w��8Ǹ� �`�yl�q!zaBk�}f�M����3Ml�7%H�O�`�N�i�n��I^	�a���.a���Um(#/\����T�؂��k�y���T��z}	!����*���_�LF~P�DW^��z3�W�I����t}"%KpI3Y� �ꍋ9�p--�o����ݾBfȊ�\_�ȝ�7�	HӜ�z*�0sz��&��ul��D�f�.әg&ݫ�E��/&�[�{�ySM���[�Ƥ��TO�+��7�,B�bD�d�Є}Ku�v׫3?�uV�IB�O��i&��0�SgC�y�#���fl�r��7F�/߻�рQ��U���dc��,7��lg؃2��O
�{����yɎ�h����E��?���{9����M
q[ ����cx�Qo�X^�:�/����F�q����8O�e��6rR	�̃s�}_%���٧���-�j�M6	;�AK6W��H��Dx�?�o5n�S}ׂ�@��R�+�SK�k)���)�y�g��
*����{�j- �����#녮�d4[��Ti�:Ƽ������6��� y��\e� �����x��`4�����dMb<�$p��1i2�'�uhs�{l0�p�q_�L��b<�8o�q�i\�G�a�>���=�_F@�	`�G��V�C�GKQ�Κ��~�����Y�:"��L�ޠ/�����Z�SfJ9�)V��Qޜ�i^���e&�IX6�6i��	<��G�마����S�eZdU�7�	H�@N��9UG��
�ڐ��?����֣"���B��r?���f��B}�jd�}�Zi0�����׺J�q��Y��	b�!A���-6�"|�m�xV ����)�``j7����EB&�S��&&}�gO�.�!��q�b��EG�B.>9��v��TT��c��`�@+m%c����
`����g���&R���w�u�/Kt^����V�t?o��#k��uO�2_����ʒn,���Z�}7�	9��9������ʞ�G���3�d�`��3�it� n{�T�� w��,��B���u�����ڀ�����Ƨ�9sT'�ֻ�����:���4�K	�5Y����6��;?(򴿠�֕g���Y��B��<ǆ,�L���V,����l1i��K�Յ���X���9�	
����?��9;>��P��O��6F6*O(H���t�`1�Tg�ǔ.�O�4�L6��t�\��XЧ��j�������,O��&�9���'8Z�n]�_Ҭێ���,��}B|�$��8��d=��À���*v�q#ǘ�]ܟ8�5ZF���|�L���������Mn��#�p;��6h��������8���sX�|Z/-5=��E����ȳ1��ñP$�y�L(\�,����ԔW�>x�E�³s�#�y��͇w�Ks݁Vc:�O��?�V@ܒ��&W.��jC -��P�U�	3�������Һ�_pV���zY^j$aUʙ�i�C# ��H�8�;���'I��޴4�c�Ϊ���Ep}�D���i��r�m꼶'��&{O�p�Ê�X�oi�=��{@T�%�1C�D"��>T�C:��!��{A������ �SyҶ{xGjYb�Q�#�xQ���s	�߽@�ֱ
#
(�(Y�%�y�9R�\vw=�C��� ��A�W\�I��ۙ}�Y�0[� �x�q��f�{(e*����lܥLLY7?�j�m���RY��{�w`����Y2^D�����%���m�=��R����n������}�ÉωPo��c��Q����S3ji�η8��F��N��[��Qn��X�G���.�jOj��^�x��Lե�/��_�P�X4�8WBGZ�ȅ�W��������9`?ZzK�P�Ȣ�L�4Ԯ��bϊ
��������B�DV��c.��0_�BI%Jh�آ *���7.�ƻΠ��U�]!o��ydz:�{��	���5����ʱ�E�x����t� �BH�[2^�8�J������#:��?{4��N���	)��p�㨹!9=�hW�Hfx��7���/T@��1Շ?s�J��8� ��e���Y��N�s�H������I<y�.Ʈ�D��q�	 ��g�a�_��t�H�.8u0DC�Ǔ�ۻ��`鷺�+���G��m4XLAX.$2y�Ya;=�;@�,���L���K�)ʲ|���탠�7�$z5�ܶ%�������%�����D.g̴3ŰA^�AD̳�]�>7�P����*�i�m�\�o���צ�K�!!a�~����J�$��X��`���Ri[w���TW�ݪ��R(�pkw?E��㙴Y 
�q��ֻ��	gAnn��k���9ՌD/0�EE%B�/)��ӌ�LܙӜc5&���t*}��GiUb�@+�'��z�c4@�S��񌗮G��}@��%�[��`�C�#�1�K[o�fO���(
�\�`�}:�V�<o8��0��Uz4�毹��~�O;^�����2�&��.��=p;p��?Ij��1 x_m�[�$-��]�������窙R�-;���i++�����V����G~�ӱ1����%�.7�rCBk��ڲ�}R�-�1"�`쀠���J��1D�Mg�����ěw��G�Ù��)J�IO(��#���5y+QM��5 k�/^��7�M*5�WU�-O���jO��fX�1��7	 �{��WnY�ˆH����i�'J�U�'sv˘J1��iV�h֦��wo��?/h��SCI�5�C�#t[�
���]R5��8��9��xq��^��֧��Z���������O_�Y99�>�X�����i�B\+��w���,���E��l,H-���uJf� ,��>k�;
ciP-S<!C؅*�NTvǽ�Ҳ����:u���0=Ao�]go���R��}�>CT����*�e_;2ș��9����̩ò�����Uǌbx��VՋrIQ���_�T\�@Ac�4*y�d�,�ХV�F:����e����w�/C�Ϲ���ow���{S�\}t�غ{��3���K꺫�g�P��V�ɝYn��m
��Q&%>5x_�
`}������q9O����m��bzz�۫�p	�s���;��ч��l��s����4ݫ����1���1�v�N	��'��a��1J��$=��Y"nϒ>�w�L�bGn��T7gF�?Z�r��Ǎ㬠X��6�i������Όs��T%3��T���g�P�3VƊ��� ��;�Y�~a/Czc�`��u|��~���jd��l-T|'>:�����|��!�	�/yq�@�O�5��A ���B���`}C�����	���͜hɧn-�T,���O��;�`.��s����N
i�78�7�o�v������⑔|������Q���c���_2�'�z������.X��Q2��,J0�* ��b�aDɵ�e���ʮ!���$y�F������I*�_�9�c��we�Wy�r����~=��(~��'}��?���<��*p�=*��!��� Jy7���q?n�g&=u@��Ǭ7�m�޺�ٳ���ğh�d�>vo��QV�a�yWcw��s��G44�����q���K]�9p��2������K�d3���9�8�=� ҭ�Nr�ǔ˖���H�H�x��dfMeL�?;�Yf�F�����5��x��}�|xA_~?^u��n��b���%� Q2���?�ͪ�{��%9E�&_bk����|S@{ ^���Ih�@��g'���7�C�dkB�N�e�Fע��j����XoM|�ϩ?�r0�:�@�O*�4]�`�y�EV�1��f[f.�NDc��3憏f�[xS?�-�ۭ}<�o�!vM�񄓳��	�nŒ�'s9
&���6g.%.�b{��{�H�E���Q/D��?���A��-�>�o� F �|�#6d��pmm-mEv�(���N�.�Iم)�н5��լ3�~)w���YZ)�|9�@�_���2j�2y���>(��x�<((�{�;�l�}.Ogp��M#&� 3�$lS1;��̐e�E|���"�6��Ĳ)3�Ax���ʒ�4��/��{��Le �x�@g~1
%ZC�	��}��78��6��Z�� "	�M�b#[dQ�is�${�6y7����dΜ���y�N��&c����ŗ�v���l���c?X�ƾ���.�:�EӣGd�BkBN��ku*���'�9��dA���z�ĻˆL����	��w����k�S�3��[5sr%z.���gWp1��Y
�>��q��m���/�y:�����+@��$�o��O� (�E=N�X��4'ù���R�<��s��}]�Rm,}9Œ���Fe١��I�ߙ�M�C/�^�Sl6��tV������0gp�<��"����^�Ae�&��������7�RrTn��/���%u/���H8�%��+��x��f����q�b���L_6������ӝ_{�s�񿻉K��(c��7W���`�������>Y��`�L�z{&�$����%�H=�*������ ^Tr.��%�/6��e8ش�b�aq%ҩ�Q����[�C�FB�	e��W����1-n�c*�����H�s�c�lR�~��t���~s� ��C�D�B1]nIk������'>h��,�:�����Ί��F�>�����m��Ƽ|0&!Z��J� �}[��?'�nw�E)����~=�i٥�V�k�	[vmM%M��I�A��ɤ����9��mx���>�Hg)��P�%X/x�\KXBBA�UZ#WƉs�r?Q��F����Z�������N](.e�پ��*:+ȟ��l��]�9����$�����U��� ^�m�YɁ�3���ڰ��`����V[]�ϔ2#y��i�1����lh��.��P0s��?�����E�y,��Wa��� �JoX
ȣ*u��l	���� % �>�Z��z˓�m	���[(̘R��(Vu~<����j=����H����m�܋���?�R?@vLH¶qz˖U��F�^:�jz��������q�I�^�k��g���I�o�ي�$]��¯h݀g�o�`21��ח�;�]�	eq�,�p�Vgtbt6��؂�u*���dF�f�؈+��U�s��t����jH��@$k�Q����+���d�j:�I���)}rI���}�z�܎�?����=��&��W���E���'�
f��:�
�nD?_`�n�^�'�;�g֜�^�&3ˁ4���r���f�-d��Y;���9%P&=���t/XȆb��_,q`��Z &zSuQ�,��Ƴ��x!�y]朡˓w�8;�uz�.�4�7,n��w.�a��(�I'R~��7�APE$bg���I���0�>�ߑf酅�r���G�o�`>��|��ˤ�>�K��m��ɭ1Kyz�G*,yDV���i�3U�K�lE� d&�7De=��$y���XRpi/o��F�
P{�'�kz�Ͼ�Ԑ_�+|$�r�y�xG���:F�����.�Ym��R�l�AW�����/�?2���.d�xI��w�Qb��&�p�\7��@J�T\����5`��&��_Y�	LrU��`�Ɠ����@V�ǎ�����BG��2��d�B������FMv4���,"v_����a�}�ED�Q��4
nK�~����a��%�ܷ�feA�o��a�����7�h�Jr^sKFIC�ͯp4}����4���/�"�t�t<V��� 2�8Ǥs4�� �[:������U�*���\���m��I@O��ne/�8�((1�߰�`T"��}�ݔ���W�$B}�tS�wV�w�+�y�~�;��g�����d�\�^��Ӽ��x�
�d�z��<!u
��5�E̷b�_�N3��z�K�����)� Pnz�zIܑlHh��H�7 �w����;p5��z(!�����?g���~�0�>"%�}�z�+�E�����;�E �/S�I.�v���e�[�4�,�����%�泞�Ϊ)V��q$�_s�2���t�-n���o��pV�9�n�"��Q]���4�t�#?q���S@Cr���i*'�bV��Zg�ፅF9�8����U����k���s�����O�2�TcO r1;�Qo��jD-�2�s���Aw��t��K\>-�������ʇl�JX\�ٚ� �m=/9�\����]���}p�ԭ�';�h.�q�PO�uz�ڋ�n9oi- T�A3@?ڵ&�}�a�%����Oچct�`D#�b�Rm����u@�J�c�[T
g>4s��ZqĘFr���I�"��o�k?hN��t��u ���;Q��(\�{�)h����B��w�3�f	�٬8�� 惋��b~��lA�H��]��m#n�5������5p�.I�x6���b&�n��/�A`:iX,t��(���@ز�{�c^i�X�O�ʅ� %瞟b� w����b�-�}���D^����Y|bg}:���L�φV�̗+��!��,�.�7�)�*�4HӅ�͙v��������z{���Η�x)��`�l��\8��x�b>ЬA6��_O�Sאv��}&���x�3�M>�g����:�][�G��e��@����[����������C� #�Έj׸�����*_&k�PK   �i;Y'(�5W �@ /   images/4737cce6-ef6b-4e79-82eb-dab57378d86e.png��?���?��*�N�Y�"<)�J�q)��+�9/9�ͩ*������i��"����ls�a�9nc���~=���O�].��?���t�^o�wL�=  ��߿� 80 �<t�w'�#ĕ�c��]}�C�O�!�������[� ?v�{Z���n���<�{q�>}��B�
n���O�;+@^�?�5D� ���~Y"}�~J٤��@\�,�m��g�;�o��]Q|z� EC�J���2q�D,�۬>�Xk���i�_TO�h������T,��@7A�}½���_ؓx[+��3<�������9�X��,v'�W�K���R��2���W���&��0� ��ِ���MA��+@]A�3JY�`���=Ɲ][h�Fq�M�p	@�3�Y���>j{~����;D�oy��s��-��y�����'���������߷��o���۾�-' �o�����������Y�w���9� ��2H*T8jfVtðKݠm�촿�h�X$��p�Y}���03a�H910�aUv�;�bg�"�gC��wf;21�m�1��m��K���0vTss���t�bbf쒻����|��F��C_���\7�.�2�%+���Q���}�Ȫ��dVO���7Kj-ڲ�v�S�o �>� 6{H��@��|��k̰���D���Y�>%QO�Kߚ��;9�ܠ��ܯ:�E��g��"�4TfIW����^�m"�ck6?[��;���qz��Z򧹤w��� :(z��P�F�:�G[\�'#�vg�#jKKʸ��Z���W`zb��+A�쫯1�\~(�J>�T%c،��&��ݐ�N8����_�h�l~��}�BU6�2���|!�`�u�OЭ]mz�V��"�����"��ձߪ\nC#�M��E�`�,��OV��H<���dP��)�����t�ӕ����E����O�.9a�q���:�bug���(�B�xg	������T_1c`T���Wcɟ��jܺɉs4�7k@$W,y��.�h��<^R�Wo�!����|(��/]�{o5Hn7�ǔA����4�//�蜿���%��6̋�)�J�6��7�a�/(N�˻@��wмiL�~�[�SLi�$S��q.�b7�_*-���j��Z]8Dj�'�^����cRe8��_�=+ZS�N����X[��MuF$���I/`b���=�nboZ�A�z�����n����42�����3��9��5�^CQriJ�>t�֖�q崽�j����֞EsV��,�(��>�u�w�8�$1�L�sd_�s�3R0Ոn���������r�bZ� ]߅�3�i�w�?��,oީ�����R�Tb��4)�@�{��u�GvލZ��GL���^>~ڥ�|u��,���Oٜ��W��Ij�̈L/|^7)��d�̰^��҈�	���y���	��v`�_o4�}��;[zoå�\B��fk�4N.������s����Ы^k��nH~�p��"�!gb��T\�{�O�L��t�K�Iw�����Rdl�d��B�oR���e�m����D�����h�qC�����Ҽ1.�*�>Q�>��c�8�
9�#��DVB���o3�mI+��5
mT� �hR�2��a�L&|Bn��^;���nM��}hq�W�΍��s��*Ʊm^A��xy�ڐ���ã�_u}Syk7q�	KeΜ���mC1*"Sw�&���(VT��-��>E��EW�t��ԫ�M�ce�.6{I�H]�sl���9�עQH3Y���KϦ��*��.Vj��g:rb$f�~��	m�'9���S�Z�Բ�(��2�s�,����_l���I綧:�J�B(ra�����l�.��ɬ�h�������H�v��/	��´"�8
�u�O��A��3V��3� {����|i!A��WNp�Ah��0�"�����yC�Pʾ���U���.���ه1�9IU�-�v�_��|�ɑTwƥ�0���۸��Rh��љ�±g�ckt9��OE��Uֻ}c��M46#5�2�����s���3�wNp�d���}-g�'�w ~��+�_{���UZ���\�m�XiI�7�r�'b����d������Z��'�t����5B�:Q������ti�-ܧӔ��0 ����!�ݎ��#G��ǧQ��5$�KO.�/��ԣ�P#�Ẅ���1z��]�C�>Z� �c���	��J-�ʺiZ2�xT�����@�>��Ӫ@��$�Gكg��on.���;y���Օ|p\W���E7�R���>9&��j����)�ѩ}5�$^xF��J��
�P/H�����a�w���ͪ)�q���Ie�G�
�dq�]��2�CBv�f��?"������U_I8�ڳ���4�R��� �}A�;-4S��j��:��t��<H93�O~|�A���M*�&�s�@����"jq_E/��1+�_x8���T�S"L#�I*_Џf���;��T�d�MSҦѩc���I��hj&�#�~��L����C`tk�� >`db�7�x�2CE� n@�Eq!�@�`�8W�׻'�w%��Z��<�������vw�>�,ͷYd��P��}�hy���qSǐ7-IXg����� ������R$g���l�^�|�j�6"�Mi�$,d�å��r���\�ۻ+~F�B��M#����͉l�����,d�B�k�G�^�ɂh���]���Z����q�Hx�C������ګ��f��nC�?#�d�<s)N�2U�RX�g�lWz=!.��H�^a�ח��@O2�,�����:�6���\g~�	ix?��z���\b���6��.rRU�u��Y�t"s����ya�4�����H5O�)`m'��x�e���n��fF���%ڪ�������(�{�7���}�L󻠫�)
䘱��9J d徵ΦtNr:)�=�S��xBN�[�9��S���
B�L�6�٭���'3@fKe�0����?��_�1V��L�����j�!��#�b6�>!��9�i��������XO��c����/�~З���eb�nj�.�������ey�F.���_���+���H�8�-!~.��%�C������9]6lt1ьh��-��B�D�݇;u�\d��]��C`JN�Q������AY�X��q���S�Ry��֑=���$ ����#�o����T���F�T"��9������i̦r�5�uٱ�}7�}T*ВM�q�Șy����ـ����!\�S^��&�)p�´E�<�_8)�3�i��m���8\��{i18W�u�Ɓ�M�5M5/f�Y�a��~wr���;�s �Ҙ%��|��REټ�#9�W��㼪�?3+�2��z�d��#�-'�"^��������Ra�}Ϯ�j�>�w�hI���lB7����;�V��/$wv��=�>rRK�
s�3�	�宮�œE��,��k��x|����,�w&$�]�W2Z�׵dD���ywEwN��w�DX�aN)��F �*Tca��m�.�Y������]��I��$�}���=¬ _,�F����s��Yj�W�n�>R��LMϋW���=��MYP�B�|ٜp
�I&�I�z����039pp4b��2]o<��d�`�؞Тg~n~�����C�����j�Um�<��pk��;I-��͈ȹϱ���."��/�o,}�X��-���z��;��M��sQ�zl����T���I���m�by�hz��kqv�����<���e���%�0�'�^��BN��� ���5���@,�v��n.C����hf��Х���	a]a���Iޟ	e,EO9�b�`��)#b�]���7
f�.���}Fl�H))t�)2�.]���9櫻v1W��m)D�2��[dow �Yx|�vw>��^�>f_��]�ߙ^��s7>�va�'s�ŝ��{1�1�4�ЏuW*���$��L]�>J�@�~A|��)ז
׵��A�~�[�\� ��?)'5�̗�{4{h`!�1��^����m�	�{��AeX}1"�Š/�����[ooA)����}r��Ŝ�}p�i&A]�P�Ik�F�F�`k�����RXx�T���X�i�X���]�^д��k�1���s�����3�5�u%�T��u+B����a�V�x�m|*^�^�g%�_��K���vֽ_��aR������h�����y~$6 @����k��{�~�%^�xb�o�����V2c�����9�6M+tc̦,3���M�ww9����.���m+n̥��B`=Y��bĶN�[$��o��%s/���a-\HqJ���sS���(Xg��	q�F`.e�x�������@�"wܬB�m��|�.�Bv-�_,���~�z(�_���b�������č�Kގ-��:��'�C��P�J��D;�Y�ON��)}/@o�xQX��t5ؔ�P0��u�Y-8;�EN8�*�F������n�>��ó	��x��ƌ��srZ
uHX*WJ��:z6���K�g��ɵ#�V�ZI��喱
1
�ea�e��j���c���!߮ ��Q�����AD��!�����_ת
�G��R7�6��O��,����L>�i����^d)O�s.ډ��MJo�����gh�U���;"G��bi<��$*�2�E�N��ԤS��}��@��`Rv��%͑nR����9��chU-�5���{GWt�-�$'�=��"����ǜ�k=��Ij�ɢ� ��J�ވ�y�~��IY�[	��/2��R!|��4a��?�����+éO��x���Z�G��_^^ܣ��M� O;�r�Ơ�$�X��c�{ �N��M흌Ɋwhi����<��s��7��1o��~�����'��S����!���:���ئ��'�6�7YM�!�
 �F��F
��4���o��"x�Y3�"U�r����i�݉�oOن"u�c7��m�����H���*�A]SN��<�1vh�����)�=1�Tb�������������Y����v�֮�m�/��ɀk�������m����FП�c>+{		��UjV;/��sx�<�8v�V�
��d���/�Gl�*Z�C�|wがQT""�ioTMء�^��Q�;<<Ί������X���s�~�ǜ*y�~'7��N�d����Awm\��D��+周�e�ɉ��P�z��C�k�I���\U�V�Lu�~5$�K#Ex(�g�%.s�o����S���\�F�{|�cv�����n�^\�69Q᳦�54s�����1ƣ�9v�o�ho�ՔL��Ȕ��|TYZKl��Kd��J�WC�%wY����c<��ؐQ��;6�����o@GK�[ܩ��߉Lr��h�(J�!usD3�����s��?8~#yg��t���~��Z�̫49$��`��KŅ]X~�O��q���.�<L�V���,��ǹ�J�.�-���cvn|���������ƞD�����>W�E�YQ	�ח��y@�ƪ��D�����p^N.�z1Sbu���*���İ�U��:�K4��h�ac>���m�۟0�W���ZbGޯ �_�ym�#qÉ����X#�=wnb������e��M/���v	?h9�N�!���j�i���=�7_��cby�#7�5�џz�g�gy�95�dw��'����CJ�S�/ic�Ãe�� �]���8y0 б;ڄ��S���t��A�icK��O���V�*9]��曖0��q³��;uY��3f/�1!o ��V\�:�z�^S$���)x��Q����
�UL������|J��Y�����/��sVY5G����i�^��*sL�J�q+�f�\«�X�P�v�6D֯G*���!kI���\�Nl�SŖ�zΦ+�_%0�~����R7�&#�7�y�oN��t�n�=tp�x7[�N�C���h�j����F��Iק?�)ğ3b#��܁����W4����O���d�Tս~�2�s�g�p�7f��˱IY���f�^�N~�݃����./*�:44�)T���#�/�<�/y�'ܰԢ�� _y���i��#.�n�^�9;�F,{ȩ4�=�����.{I)������r�4��(CY���v��_�<(���/s���'F� ��ޟ?N�~��=8w���r�z����I׈�'X�6u�~�,%m|���sҜ�y;{w�X`��O_��bҁ��VY��>t�
��skŨ�f��tR�T�e����|���`���49��9���2�^�~�l���ˍՋ���ٷ�q����%/���w��R�~��Ϲ�z�T/mp�@��w�5j�~�y�%9���H�O�f���Q��و�P��T>r�7�����>0x��8�:?����r�&4Z}lI(��$6I��$��2р�|4�;��'mt6����'2�op��+Msg)��jՂ M|����	 ,|OS�1R8!@8�-/y�ߺt�7�'���-����I�;�.�OK�C�a�jw`R���vSM�DH�$ԑ'�o�vQ	�CN<�_��h�A{��A��XU�BsG�B��bHY�9�rh��.�����.G�b}��)�M����S�x.y��^1���*y���3�D�ڜ��9ިj��f۟g��鬻%�,�1 F�|��Xp�b�u����s�2���� t�������hB��8+�좀����y%�Z���.󿑀=�^�Cb��0�#"ě͋W	9���OT����� ݗR�{��")J1&�T]j�J�aþ�l�)?�?����V�i�ɦ�y<����'D�*�<a�d4���GAD����r�w��-Th(:�"����"���)�uu�ʁ��[��fM೔ӥ0����]?52��-�� x�u���������}��5_ͷ�hx(�����q��;�
�Q�\��	h%ۤ�(��m�����3՝���T���s������H��+��Nq��M����ˣ	m���G���(jE�gy;���7���'`�� D8z��)��cw*C*�5]Y0�|��r��-�9$��Ϙn�i�.2�
Q)��uv�(���\�Gh�紨l���o뀦�)4)�\�o]�r�@U�Nb��eZkr�(�{������!�?1|�{P���d������)���kdF���6.�H�lZ�����W	�����	9x��. ŴD���?�봀��T%א�,ƆX�����ZC��4R��}冑���ť5,��Su:97!
B�hA-nQSיMAs�ugjlO���:h>�<�*���à��C~c�X�錄�X���O��X/���_]�L�3U|���|R����Dt��Ӱ� ��g���������˲m-���f�u_�=�i�ꋖ.���
Q�	+B����s��J��~�n�-���;��r�p�m;1�'��D;3��jEt.n�� �����/_��_�������3'���(���EK��$��í,�����@��z���fQ0�_��>���?��0*��<"z�� <[�'Q��^h��w�c�~(�L�����\T��{����~�a��N�f�Z�2DO�֗�RXJ���N4�R6x��"�e��Զь_+�9�,/���}����E�Ǽ��m?�n�q�ո=��!�a�}��6 ��=���fч'�M��j+�P+O�j/)4�|��`�4��U�!C�����6�C���ôl��LCO�h��]������Ԝ4����6Zo��L�b"K,�/�k����Ł���
3���_d5t���fD�(��6q� �+�`���ol�^U����~�>O &�/y�ϵ�w�V�u�y�t�nο�ؖs�Mg�T^�Rӌ�NR�����BBdiZ��Ρ�$�q׳�[M�'���C�ۦg�����Aҏ �ҋܗZ����K,�*y�f�syM]�
\������R{(�{U�ȅ��Ë+B�R��*=�ۀ�O�A��'�(q�z'z,3��!u�Q&Xp����c�����$��s��n¾t��O?�_Ij��p���`�v�j8���1#�bWL�}�oK�7L*:.O �o�׬������$t����7$L{y�=86}�v�bb[�RK�KK���+����];��sssWh �����;
�Zv�Q[_��_Nj7����R[���7:p�*�#	�I�k��&��]S^��2���:%��9��[��J��H2�^�iVONd��1����u٣�FB6}NU�Fmp�!YKTmbQ�1T,����iX���%*�Ol�_W9�an'S��A�4�P)��7��Zx�1O;3�G+4ޠ�?�ɹ��H9��s�1��2~jkl{Z95j\�O)���p{qj���
]
Ny^��d��*����z,��9���?��~����{�Wݥc����8#���Ps��՚߽&:q �jwz<R ��Y�qW������˷]q]gQ	���9&O ��o6�5R��|���Q۩k�/>E�e_��'2'��}΢�<��8S���7�f_�,��sW�Lb�F�ȥ�z��MHc�#�:"=� �����q1�����X`@�&hǩe�V�Qҽ�钷j�K"�fI/���� O����hT5T����>�9��^O
e��r��K )ó�ьMqz�EP�v� G� S3�(�q#�̞+U���9
��}j[Om�7��Y�(3�v�{��ot^��;9*�q��C���G��������ĕ=B�z)?e6,��X�Z����JS�[I�M(�`�J�ɭ��^����DU6II���0����w���_�c.:��Q� ��L�"пbc���ȑ5�w��>�1�X�*����c�ڃ���WEed����ࣗ3NO(=�F+��\q�bV�d�~܃�e���RѠyc��H��L��V��P�^�wi^#�����m��̻~�@!G��PO�٢�N��{�~6yY*?)P<V�Ut�va|*a-v�S��a�
;m��i��3x���}�n3CX�Y.mX}�Zoc��/kd��Z�|8��􇴯�s	M;w��?�W~�����������Ww�v��%����Ň���|
?Q{miz���'�Ow�o�y!6�t^�|6_���lߧr=���B�����9o?��g�8ROդ9M��I����Q���g� 3M�֏p��� ���A���s�7�m�0m��L�0T��CA?�rp�|�d����)iTg�Ͻ�	���r@��슢��SMXN��<B#,>Q�ˆKp��\�L�-K���G��d�1�$���q���ieaj% ��]j�o�-�Q[���K ���
�9^$�h��2ΌF��������_O;t�6������� ����	�>�*����6~pD�܇`�`�=��ƕƅ��28�J�p�!G� CI�������s��ǐ�zY�?�<n
�A���:�z���|,_��Ӽ-��#�@���>��@�m��o�.:rH�G=F_]���p:g돐�+x##|�a�^˖�X6W�
nFo'o���[9�ƭa�u1�vWX~ڰ��  �k]	���r����mz�79_����N�k�j�	w�� #mTO��ZȜLH��(N|V�Q��dr�����9�~�����AaxM%-��[B~t�A��y<l�P!����Ƀxл?n�  ��yc��!,�!��ȩ�N�����I��_���RW>g�8�*��K	=���>�8�㈱�i5Gٟ�dv.�n�2�Ȟ*��zO�G���\`��W�K!��[6m����,��K�v`���]Qȣ'd�yq)G*��.��.Łjұ���A�)X������'bku'�"�c�2؝
�o@����[$���Ƭ�7�-�+���.s���"<�u�����XI~�v�mI�1Dn
,��^���^H�{��]Q�D� �����
$�{���݅�K\ V����BqRp���i���B��5�	�s�!F`+�{]��	�7�(�{4���H��7���Xb�����xf̽�yfο^��OAV
H�ʁ�a���P�0]�z*�=��2�""�}}�8�Z��㴑J퐐�E*���e*�֟}aegg'�{�.~����V�ڿH����+��7S�,��5s��@S'U��L��ը�0ݸ���o�?����$�
4Ʋ���С�'hz:c�����C���Y�RifT�b�v�Ȧú�~"��<�ӊ��b=�D��B6�1Q��Ŏ4{��I��	�����E��>>���M�M��V� �W�\��O}�r����/�>(�RW{�3�����x+*!141�e�����7fR���5�^��kuL\\xlͮ�LN R͗|��N9\X�`�#µ	���Ek��THQi��=)�8�6_9y7��f��r�>�g#����?g��3;��i<ox�ܮ�������XH�����cu��H�������� �-��_��}�j0�q k߲L����9�\\��^��?G�6�zL@`(�%uV$C�>z�Q:���Ij�=A��DƆ���"3EJ\p^]g���^_�'5A_�Uu"�-Жg�·�@�;��>��<$s+y�	t������sg2Uй8���=F�m���|#��ǎ��rV���My��|�i/��	@�����^��,l;�A0_�Ryg��v@ߡ~��u~��8�u�b��%���/�}�.6c���{X\]�X�K�����U��\Ͽ����?�)f�1�����^��NR� qE��G�����<Xg����].���N=R���!ja��o*�e�R*L��������[�rj�=�P�[TT�)x�|?Ԑ�^�?D���(��Sg`�ǉ?��j� ��ʨ�!���[m��m��_��׻!�O��ǧg�C=��3�(��o�m��l��
�I&&�H�#�i<t���'��Ŵ�0	�W��c"�$H!.��<v��|��0v��6!�����������.�E��}o����g`Y��i5غ+�G��0�e{��?X��Բe銃��a	����x#gA8�%��0)��#�dO����S �p>&�恄���	�-0c>n~��� �[Ӂx��7���&߅��Co�m��,���#�2��)2�ou����l�qy�m�Ѕ���O�<�-��Β���+�ˌ ��EQ�#4x}�|E>ux�D�s�'em��F���:���*��l~�Kl���P��(����ɪOOW�>*�<�(��'#�/xIQ?߈"��G+9�_�}=�j���-����
^�����ȼ6��f�bx1,�J:�(��[�S���h��X���Ƚ�F�_��7Cu�	��̧�����e�}^�����JjRUb#�'��� =�Xz�v�,)�Bح��s7{&�W�C�}*Z��aצ��2$j��ޱ7�E���� �����p_H�v]�ZcN� 7`d���!z�{����8�޷@s����k�?Y������������|�ʤ�o�|�?u�W^8���O4����3�o9_��h��,%��j~A��s�G4YF�,;���[�_d�7P���
�.����PRR��N��Ø��/_��j�?HB{���BK���!��:%iQk�W�^w��.f�ܲ�Bim^ck�{�?v��*dD��|Hn�A{rkg��TÀ3�"&
�S�3oV�4�4�`�XX����ٶ�Q,��C$��8mg���$���؍!� P�7q
.�eK}�񣖢��$	$(��'}0|�7�����{��l�o1�q����j��#�;}��"PT1�)ͱR d���A�f�N�ɰK�=�G����Ğ�P�5"�:��=YS\]=�^5Ը��˕c�!��b0Z��*¤��7�)u�Ch�<j^Jr�-��C���T7�����Kd�(��Z룇�������ۿϩ���զ�g�\�ޭ�%��g8͊��#�M|U����&p?�wu���CZSէ�,Ｖ8�.~�r�i� �дy��эO��?���R[*�=�	�/�l�]F���m����z�`���ʶ
p���5�fW9������'������*���ڍ��~�0Z"�A������JG����Ɲ�rj�ֶ�|�/y�Jiٚ��*�0�2i���
tS�92*�Zz���ohŴ`mxI�,�=J���mQ%+d��L�^��#
��N.��.w&80ŲyU��ɘ�G4��W�@�e�h�T�?�O3�WN�;W=X�|�.���)_hX��,7w�H۰�!%����H�tC���ߢџ��ME�q��S��gK,�4n�K��v�D�[IcJ'��={e߳Ί���Y���r2�0�|����E�?Q�,|h�l������G<��SF�+�D`x��	�*�&�0���4��+Ф#���h��D/{�x�	o��>4S�w�{�<��v6������7=����&<*.*�}*�Φ��20RL6_�x�Wɇ�_��.bP�uV�Fj͸�k�`�SJ�g����[}}�f[����t�U�������r�2�v���O/��
`桩��'	7��S�h�J�GD)�L���K�e��g�1%|w�mN��u0��l�i�y
�V���t<~e�˛�
n/�vJBRC�I$R�o$`19�^]���o�T4��d~x}��ώӻ�< @c& ����%�BXt(:��7�T%/k�2k�a	��@��J�
�]���!���AK�Ű����\�B[z�!��o
WUSU(������zT�TИ��� ;���UL�"�jb2,��ШQ0k�\���)�m�e?��6�a��I��B����ꋇ�R���J�}��НL�����+��ywd^>l�	��~?��uJ	Ainv�ܝ�.2� �x��t�t�uɍ!oւY�!�<�
�X���PB���*�K�V��"���^m�i���'y udȢ�0L%�Q�^����Ⱨ�6[��عǨռ8��3|�3c��zN4:�
�ߘ=`��h�D��܆tSW��{Wc�s�!Ý���ȗ� *����h�I=鬋���dK�%��~��{ı��%��www������(��z��n�&J}���Fh��l]p��uʕ�w�Ԟ��T&I�����?��v=�}�iYf�>xB���se��To�/Y��Z��ļ�dMZ1�-��p;Y�?�A�1�k�I^n�ɕ�vW=�[��*P��wX#:An����.�t�Ʋ�<7cE���wynv6�_�E�FZw������?�e�p�p݂Ka��)S:�gF�r��ᓘp{R��=�6��u?w����.���i?G�{��{N��)�����FM�������_���\�Ǝ4�Dߔ*�:~e&�0M�K,i��y�m�du���só���>Z=$}�lKy�ְ��N��6p���6�w���J[037�#��s�civ���(qK�U�A�ST�.����*X$�P)�7o�{��n�eh6OĮW趒�+ӌ��oT?����U+�nL�~���$I�Q��鷀����;�s�?���\��lY�49xk�W��---[�`���U�-c�8��F���3>�tujsR���ր��Xy)�	��Ϡ=G��ո cy�Q�שd����R<o��ϽR#=�����t����[�Gm5��VVZ�ɗ�Y��P��;���`j�����;���(��g���&�h�3NM-s{�f-,\P3r�LQYi??)˦	N<z�P��tg D����
!f+��fR�O����)��pc��EK�k�Xf��&��1Fx��Hoↆ�V�4�@ �G{�2|_�n��ȥ#K�&��+ޮ"�ޮ���R�����Z:O�ڂ4�Z�:�[��roI������{�n��v�`r��m�����PR��vwX	�@y\���9�k�4

"���l�ձ���ּ�6`�K��-����
S�U8�2A�9�7e�sH�q5���p��@J�Y?� J�F��e�իW����`F���S?H��t���$�ݾ�ߴ�:0��ѵ��C�nD���ɐ�kw�����o�q���J�@�_*�����U̱+���Z�A���4\�K�(U�"��=hg�%a<��>M��@Q%���U��'�$�XϮN:'�hΏ��>�2�kg����}�e`3B?��]���Z�b�����GWA-�U����BK^)
m�z�~��)�2f-"���x��<N��	��|}}Kȡ<&:Dg�y=�
\�����q�����~l�}�Q�V�^o�a�j��� ]���jJIf����f��������pf�17�pV���F4����w��CPڹf��:�HJ3A��`s2%���X;5���h���C�vGs���FDR���@�֗^E�g�
W��w���4X;[.��wp�&���lc]����a�YF���,����XҌF��Dť�p@��}�ۢ�dd6��M��I2k�~ސ�B%��3B��4\�.�]e���
\~_�XF:�P��#����YV�)z�%��k�a޼�U�ߣ�04z9n�wG+���+�����%���rؗ|O�?�r����Pl}�})�BC�zZJ˺�q�R�dg�Zw������c+�R��|���f/���U��C�yn�`Q���Kz��@��H�MH�OQ����3�P�{j�X�������b�:��߃���nR=:8ܴ�2-F�����Ԩ�W�"�E�"��]�/!U�y/�\���U}����'�u�X�Z�\�|@Y�vh-~�_�x���
0�-|
��qJ�o���E�w$Q��i����R�ȯu��M�_Y�ʭ6ɽ;Oge�۶�B��RQM�5SʴvN�ph���!��vm���_c;�/C��j������8�G`�<
�򱃧ԑd�6iL��,uYb��B'��\�VZ����T�@x83�b�jkj>� ,�a��~Vc�f�7/�a[�WK�|�����V���=������TC��iÏ#G�ի�"#�q�+���9��C*����>��}@�J����!S�%7b�̾2A��S�];�Py�~��|V �gY�~�Q�S-��� ܢ���ȑ�{�4}޲�I����Qr�Қ�?L�9����̀
�%�;�e,�_|�N�2X��߻ #���6��pP��}(B��4@�������h�VeS���h����z'�i^��`��v�O����*�H��Kaas_RC��SZ[�9��.���Y��:wR��T_�L��E[��C� ��A�X���@4�a�
���`n���U�6�=O�=-1W?����î��^��6=
f�حK����-..?�i�eA�;�"�7(�ÊA�*��Wx��� 5��8;�t���{�qur�9-}�q�_ݧ��N	ol:*~k�􇰡-|�"�ţ���� ؃W�Y���rj���j e8�o�˧_s�Q�ي����n��+l�	�n�ƹb�F������'k��Ƥ�W�s:$�I��'��l`�`U�Vvl1��6�^��"$R��az���CXicꈦ�j|/{��#x?1�4��l%Y�eETh�eʳ�,��n
�y������uK�H`h���cjf����l�#�9X��J0�3;����KS�3��Ōeo���e�k-g(g�,@Qd�c6C��.��0Wp���P8X
^ t�5� Q�'?_��q��q��]p/��N~���}�y���z3k�AB��e�gw9Ws�|��g`aI��MtD�m�fj�� 3n�F��:�Q�m�`��5s���t�cu�'��?���q-|��W����͝����VI4fH�$�������St{Rl.GC�o�(p�QP0���4�Ԥ�w/u�YPūqovӑ�-��ձ�N�X;0TJ��X���0Ib>�`�a:�d�����-�N�����L���H�fM�����9�/J3�a��`^�I�=�N��y��P�����;�i�Z��2jӱ�H�O������`-�S�؆<�Q<�z'��q�~�~�wƏךT�֡�O��K-r��e���3�z]�� 㼈�O�ѩ/0�O���ơ���U�]J��!���ٗ�N�U�!A�?F�+Qs��=��j�8q�/���	~1�v��l��QZ;�[�Sc��L~�# �>�LK,\�0����A��TIH4H��&V�����S�3!���j@�W�����kN������G�/V_�?iK"���[��غ���}m;��c�c�)� 7}��ф�kRhƏ��%���@E��M�cZB��b�A�j#������-����j�
:ʚ�YL��O�$���ǖ�j�ۅw�mvH9�٥��v���%�}����*y���)*��r�q��[|��"�8���ݏa���h��s�	}���N�Ci�{�]�Z3�K5��mz���L���d*��]���ׂw;�������#Fd�7����g��,�=.<���+ok�j
ߴV;�`S�dV�V�6�.��z�x��[����`������*�n櫶L��>����<�����/濎j���RX�
Y�Ⱦ�w���m�
kZ㦻�C�ST��9���H���K�k���e��Q����N�<�}
Y$����S]��J?�NO��t�PԷL)[�Y��L����1��qM���8)��%R��))"�"���0:�Q�K@0�FKI�1F7�a0ꋯ���x���������{��~�$��"]im��H]#Rj�~���^��mk�2L�I3���q�G�T�L��=��CD����hM*��>_[>(`����Ŋ��HCOc<��F�7��Wu�Wq9h)IGj��:�Y�)�!Ă�rS���MvV�~��Q��tM�%�=W�Rg�����������5�V�x}�{XMܞ���B�z\2æj`���=�;%����IxV�[@5+��Kj�K? �\/8����I��!z�1���M������}�=Ǝ=����bjS͋샺mD�T������38��P���/뻳qR^�k��L���tS��p'��P���/� �޹�7b�~oi�"��/'&\���0 Ǖ�G���%���շ����ʗX�^j4�4`���ĻV��f��ӇWJ&��z@���1�G�1Q��t!�Vg��>sV�����k�D;Ƕ���]�MYh{N��)_q��6|r�E(w	�k�'%�*���v����N:��\�dLg�g�O��>ϗYLQ-�V��%�œ��8��e�͢���.���{n���;eʻt���m�= j*�cfw��SH氛�几�����.-ޔ\Ej�"M�Z}�R,��5��nsX�$V�$˷4����yz*PO��L�X-��{-�&�x_e�QB�@�ȇ�f	��m���;�h'�:�)�X��=�=R��|��gH���C���7��/�F)u�2M?cbZti�\»��m���e����ˀ�I��ȫ�|� -�6��׾�R =����1��ߜ3v��mB�ކ���\���3�i�Fm��n��=��7"� ����8��y>�Ɓ��Y4��t*�{x��8�����c�g����4��U�"��j��iT��s6�R�8
�q]�	��U-�.A�����5���C�r���=�}dI��zP�������U�͍�`�ۦY}-�j�G��7rO6�{plνl�}y�� �:)X��sr-�r-A*� T�rf<� ����!k��U�-� �>��I�G$8��s7�)�ڎ�+vi�g�w��Q�����Q?�R�?�;�Î��4�*;/�>�}zt�n{�%�tySFEBok˗�l�e
d�^aI���y����(��Aӯ]�b߷��2�>�`���7�?9�OӶ��l+�Z5X���خ��m7}�S�TMX�v]7�,[���b�ٯ�w�R��)�����n����ڟ�#*�,
IIМz�����U�$q:u��,�F�Ļ b��5I�'��:��!���v���4�3\ϷZ\m�I�Ȭ���I��q\�]���U|�r�Lw��J�?9T�!~��a�;�׉��	Nr&{Df�d���.��v;!��{�	=�f63�c�P��(�kDy3,��G�1���m�d��)�j�X�̛h7�?`B�[��&��.zze��~˷%!Yf򋷐i�8 C�{���U�E��K�7����W'��]�^lPFz����q��d���H�+�A9ی�w�5Y�-��]n�P��m<��W��-#L����2F7��#s�o"�+ey�x0Q��7i ������m	g����״�8�6�ac�؅��yn��S������7�V�n#�$Gv��|���s�.Ur�3�9��QUԀm����T�z���z�"��(cN���,�.6�yߧ�+��z��9γ��N����w�T�qZ̊��)�j��Cۡ�̯@���*s q�
f�7"�~=�6�O[��˻�^�{��*������@$l�~[m=�L�/�Z��M��}_	��_��4'o�P^	��`� &��(+Y�6��Mf�D�y?%O�n�ch�_t�@�-�
�%�;_=u�X�%��b�7F����?�ݖ�O�a���F�2D���\k�O��ϕ�k��^��y��{X�x�r�b��|d_�mM�9���G^5H\+���\/7]\�4�f�~ ,��e�3{n&���*���j4�ֹ*i��)�;�Q�c��ۘ緋��_]��C�8W�st����}���A:b-�|i[s��Y�ޟ��B6DL{K�}^Q�.	��r�����+;�;@���=�����4�L�m��D����M���.�Oze�y� c����6격3�)3���z(;�'''�J1<�<����bX!��||�&�[҆&�#h.?7W*�����g�pX��B�w?T�8��rrdI��X�̨������W�+�q�,IO�"�(��������T�_��1��2y?���7撑N;u�:���u�p,r)���)AP~�_f*H'���zUWLw"ڤ�� A�w�; �^��Ҿ�j/�J�z'���r��1���4ei4`_�*O�����LN�?-��ѷ��Iy&Y���#P�� C>c�6��I$����/#�Yȟy/���!���Y����R�|n�B!ϲ���k�0�l��R�9�ِ�{��X�s���m�iJ���̏����Cn5�9�*����)��y��Y���T�FoY0��Ol�A�!����ا���a���>����Ͱ�:\�" ��~����w��=����cYx�Z�1�M�H�6�ߵ6�����c\�.��HF��/���?�{mVz�Yfg�{�z����(�mZr!�y>�(QǼ��L���1+$_O@��p2h�@��.g�CS���{�w�H�!>aT�.<z�'��%Zuq���J;kx"���b�XeH8>���@�5��3ļ�/ۜ+��G��ݻvxw�c���:���阷&'{nfO��t�(e�����n�u֘IQ���y��z ����^�RCuu>_�I����;��[��I�A�5x��y/�ֆa�e�?�����<g�_�R c1u�U<ţ|t~��ɘ#�*,�u>�˗�a�}��s�n3�2tINǅ��!�k�m���M�I����F��-R��с��W�u��D��u���F�������-��xMR.��YUP��>�S&.����o�L� �oW�a�뵬
��0�z��E�m���4��3�xG�ti�|*N�e/5�Iǅ�����6�1���T�����Nh�uq�\b�|���Ad�5t����:b��itd�^�y�3���e�aT�2��B�o��w��.���ר�c3pBd\85��&��U���"�2!q$�� ����u�_�}!$E��`s�~ Yu;����*����g3���lU����x�HY�7���1#q��{�^��Y����חQH)��uV��!�&�6�lZ��M���&��2M����+G����c��H�與fn�Pa��C����u^�_z9�]��Q�W�I�Ǵ�E��>�ң���3&Gh\
�H_o�6;|�_�0�uq��y�%+��O�ڢ38R5�s��jcndM��-l�,zCP6�VF��.���e�`f���p9�Z,����>��vk
�YЍ'�J������f�J�Ϛa��ڑA�7�2�h��K��z__ΐo�e3��xL�h�|�[RRBc�5ӧx��ڕqQ�S==��y����CgO��M�m�H��MB�k�6���s��'�D�L,Dj�e�W�иԠ��9N����~5C_�����7/]�e�0�5:�����I����3��%�_�s��%��pq�z����w
~ʛ�M.*�1d$+�lRvx�Ej�C��U�Ł��^�s� g�&+]��Q����Q�R�%�т�ҭ$6��QB���x�dVG��5����^Wb�ti��oy},����. Kf#C���^��g�č�N�;-���5i���s27G�����y_�^�{���k��߁���eQ;Nz8�S	.R���$ᤍ�Żv�=n�L0��-��;����ׅ��g�!�a��J��^ ����	!v���Yl��0/}HV$i�`��8�y:ZKЅ?�q�!�5����{��� ��:�h]��1�f�������u�[L���9�]0yF�ޛ_��YP�@�-��S�(�&�v��E�3bݖ���~@��nm /�Z�N5 �b}��ثS�3i9�r�}~��ڗ����xjF�V�ϻ��N��SuEmaO���RvP���ݖTS S;,�^�H>heۜ|L�<��~5�(�7�>�G���Ʀ���h���P8Wya���	��I��;���YL@0"�j)\�6�+mn.j,��� ��0{G	��H�����/�EÃ� �l�?�[�k���������4�^)�V�"� Z��L4�����I�̬�s�3���9���d��)��>3fz���"��ȇ���4���&��)b�%�S�yp��%;#Z���V#���k��Z@�Q;'|x�s2qkV`=�ǪU�Q��!-N�7�S)�2&Zk�w��1O�C��#ɻ���=���4k;͏���o9�$�:j;r�N��q��$��'��i*h׻��O��(i(:Ư~~2"��v2�`r�C�~�_FKyܿI\"�y��v�+}&c	�ҋ�>WJ�-���S�#�������
S��9oS��{'�����(5s|0(�S���i���{�K|@H$2_�sz8��ڨ��D:�����w�xٛh;����i����Ww���"���M�ڹO��;��&��;���)U��E�2�Βl�&:z0����z�K��lu-�!�#m�ô�z�#��]�o�Y}]OWS�8��kK��2<9��穹��,8s&�6}TЬ8��W�p����Wk~
�wQ��N=��8o��oI0�g�
Z���E��>�rs���
��P��s��"��=�P6��zZ���c0f52�@5�pJX�@����	Lh�N�Ɍ���-�s�>�8�"P1��������� ��7Mƻ��
�� ?��5<���΅��NY�F��l�MP�̭y��5��y
vx�7Kɂ��s˒�,�?���y�i�Y��b'�Y��>��и
���<��y��{V�w�:ۥ�x8Y�^)�K���dn[��z- D^Jj#g�J���"`1\h|���U�&�U���n�b�c�3��V�K���%�P�mv�ٹ��|�v�tZ�c��HXR���%l�W{Wo��4u#&C�0D0� SL^��/;��-;���E���\%�vĨ���lD������f����6�7�*�q�i������ў��D"q{e���lB� .���3B��nd.�!yNQo+�6�N� �b���ڇʭ�X�Z	@Ri�E�Oz�'m��h��5�2�Eb���sT�I$\����C�_��9���3r�{�Ag�������!JH$>�=�c� ǚ��.�q��EH���K�Ѽ�vv�������s��"c[���E0cx��<=�������-�Yi]�/D��f��S�[����gIjO	0�$��)�+�iî����m�n�U�3C��f�� q]�U��l������S��g[!���كW��5>¦���b��-���U�=O�|��Xy)i�+�st�٦�D[��{�{!���I㠣m��|䳑�Y��sS+!1�z;���c���ov��I�B+��z�~������G��:eu�A�1���/93i�^|��>Y��d����� ����.:�����N�=9�Y�ď��`���m��ϔR�:D?���}
�0�\�r�/��'�x�[�����VK�&�/߃Bo�>`�8�*��0|N����P�4�m~Ox��j���D�M��dKhS%�6��
�O:�K��D��_Q�����A+�:IDHasE(��p5�f�f���8���}�r��)��'����ŕvAn:���"a+>��ig��4,\ml�]�W�J�{�0r�����%������ϟ���á�S�<�5�+�s��٦�H�8��QT�����3��^X%�XE'�r*�B���t�h�7O�e������:�SL��|��d�b�e�������D���#�Y�R��pM�������7F��_ɅDoE��1HT?)l�� �~�l����-̢��Ha`w�IC핡��39k?�tn�Ok|���<�V�O��ҩ���{��qW2$Ș$������0�Ձݒ�,<Tԝa5en/U%�P+9�m��Wdf9zӞ��T�� �ۣ)3�.z.f���cgc0(L�mFy������w��z\�oU�蚹*[&�7Җd�v�,/� 	��M���%��^ p|u��a����Bj���9$�]ԤQ�9iS�.�M��H%�}�p<S�rᑝ�\��G����9�%�E��%nխ� c68� ��n�����N��&���$o���U�C��ڣ�/¨���*"�W�ߴ�J��]�6��쾛�}�&�$�*�Ϲ�yk45�f����lx&qv�
)��%~��zG�h���H�G�ܢQ�9ܡYq��޳i��N�g�րm��Ja_���V,��.ز�6P@���7=���T��^��ɾ��런�ݝ�.��:G럏��
��*ͯ?�f۔����z������ŞLz�*�sP�Z�ZD��*����+���S�!�n�HIoFZ�}%��t����w �x֒�r�/��3Q���݈��l��ɠ�'p�'��a#/���x�x#m1�ZHz�����k�7y��w���Pk��ů���Zo�S4O�����(����b���o�R�vTq�"�d=�;��Mu�.5,T����O?Z��i٩_fǗ)h3���A����J�d��������F���B6	���PH���֌)�q����%C����?s
V%<M	�R�4M�	(�L�2R�W�E8����Np��>�6�|ʖ�b�W��P�$�nb���bVD?�5����W�<�#��N�G�҂���R�=�VFF��A�{!>�V��	�x�3Pϴ�zv?�z����l��bY�e��e���3r��@��*��]ϤM��w>�Ƃ]��NSS�5;y������G9W�G]�ȸ��=����(KWAA��Ӆ�;�iaq,�@�rL#�7yS�|�����۹�� �!����M�����$;��Ë�E���Lo�������_�f�av~�[w��4.���4��U��,Z���'r"�"�څ�8�d/���+y�ȩ6a�l�|�<b���a���+?��Tv���p�W�1�2b������.�li��6,�󋜄LU��@g�Kk�=���h�]z4�}&3�� A�FC�.�"�oV�aȽ�#�,�ܽ}j����]h�E�>�(��>��J뜜[{�L| �c��>@=CV̹��Lc��|6���_�c����I���lǧ�u�2g���b4�"�Ԙ<�1>���a
���cC@�d���XL�GO�7�+2Wg�%�n��c� �Ii�dN�.B�F�_5EO�L)- �9Ae�LP�W~k<Rd��PU��:���	�W�[&���
���'�x�?Ak~�������A�7~"ծI@!�V�s��@�9��y�s־���ҫ������;��� ��Q�V
[��8/A�5o>M�V6�2�bڐ]���x	��n������O���ގ>���Z����M����T2H�|�ۑv��L�8���i�y������ylz$`:���	D��/�mя\k��~6Y&�A��c�}&!jQ�r,�뙴�H��rز�V�����h[�N���	?�_���Q��EȑH��Ǥ�p	�Z�4��A��>�tc9R�g��맛����*��n{:�-���*�?,������� 8����<Y룢���(���"i�5nQ�7��)�n�2���>]�@�O�\������Ԃ�����踳><�ʴ6�JUԗ-.�)v�`/'�[���'w�&��fd��~�<�^]6��4;|��^fJ�>���Y�')�33�����b���<)�U���~ŷ9Q��93ɗ�y+��+6�_��̾�1Q��6~��_]����U��2�m:C<���r�|8h�*��0�7�%0���w��(���0���Ű*���{ &\'��Z3�����ui��+��!]�&R�E먀�ϸbg����ՉpK���*����@���ŀj������I����.�#�����,�ǯl�=��϶��zc��B6��0	X��;��o��yt�i�;����b\h(:�I���>�K�Up����[��n�LJBY�?kq@������|�On[����A��"��,�-1J2%;*&�0�rY!_rs>�.hG��Ӄh�w�Y��.����vo���3j#XM�x����12�/�oX=�Q5�ߙfO�'�@tk���}�)r��#�铟u�{Jm�0�����l�v&��q%@j�/�˚��*�mL��Zu��E|y�Q�9�(	�Se�tK�~-.y��&s��kf�5���Ռ�'�uJA_�\�����˺��O�9C�Rs�*��|��qئm)h�on��h0�zz�y�d��\w�sl���}7?��F��� �r�H�ix/�rd0D��=/�\�Z?�!h����v(2xL0�з��H��~E�~����p�NiΫ��2�����%Y�ۚm���^�&<�C�ACC�������/��N��Ϗ:d�$�nI�5�_��[�������!011�k,�gAfI���+L�i44������@2ᓍ'�O�Gjk��G�Jn�u��|�q�Glb��b���)�7ɥh��W�=�f`�:;+����37/�t�M�{���XK�M��H��[�7W��Wi"�m��[�A�X����WI,���O�H����6������;���⃚$A���?=
Ꝯ��\0?w�Rڄ��~�ԉBƑ��wXE�J�{_ס������N��y���6J�E�`a4>Ʒ�e��?:�)�҄�� �R'�4�g:�TA9�|*�^ �r��Ls���zK�j��	 ))���3�g��^�(Aw�L���؟R�۶ʵh�l�+Y����H�T"���Ѽ�� �Js{�\�#ONN�Y0l��qԵ��ǭo���Z2�AR�,e�ǮH'��T5����������م�X�Y������Ϙ��s]�WX�W�pc7t�>���N�"�׫u��X�h����/���G�E0�K�骈��;Y��c�T�Nn߼uk��S_��<ޓ����n0``��|idC�i�Ѵ.�?��9�̷c\\_e���e*�������*�P�ޤ���}O1�Â9�����%�y����»��@s��J)H3�({]�r�qBD;��Y/e91
>�Կ�n���q�|ً������&�_�8E�ggh0�u�߭��
�R�+q^��E���w��L��p*n��+�<]��!×�&��B}�����M\�Aں/2c�f�m!Wl��Ni1�>���c�vT�z�o\*'��Os�(�����IK�8Xl=�h�\�Q��β�W��]��+��![�Y�W�D���4].��R�]����U���l�V��=va�GT��&�	��C���T�]���kpaƠ�-�U�V������B�υST�&	T��O�O�L��"@`�s�fx��F�l��U�
i�4IJyi&*n*�D������M��FKV��μk�Y�,u���33,�)آ�'<"�¨~�c���T ���M��V��'�?y���g��-�h�!e�^����SƏy�8b�������;z��D�oF5{�<v݁���fˢ�w��=��;���X���?4Uh�N"���{�Uvzf�[G�sR��Z����Q�,���B?��D~�iJ7�mɥ�x�ѯCt���ă��re�Ptu�b���)�ǅ�~���SƁ�:MQ���������젡�z�Pp�tt�|rڟ�m��\�Y����wл:_��:)��xF��!����Nx�g>BN,{��C�л�L���J�0��)�H��	�[՞��~��4�١�9T��Q^[�d�Y��j|�|8��n�� ��E �?G��<7,b��c܄dM�gLOw��u���ӆ��ג�f	���Gj��g��һ��Ţ�]�(��]���5��TQ���F'�caC< �΄@+�{�I97��H��ޠ�>k�ڠ�56g���XN&�^��ˁ���Q��x���rR0{���Ѥـ{ò=��>b#�@-ǆ	�z ��K��=��\���������:�(�,۠�������'aE���ܼ�:���]dß�� �k���'b�/�x\@���
�֬ճ�������,��O%8X�	�z�����W��&Y1��Y�����î�H+�����^�8���]wQ���;�(��/��4{<�Z�J൙5���H�]]HQD+��1�T缷ک����!��g,0wW�T��v��o^�ރ�v8?�0��5O���`��������z'���1k6)|��-����������i��I��2"{�5�V�_�ޫ�bYȨ7���6�M�2��m�l���<�pRٯ�-�f�#�D����@����k%{�\K��n�N��7����힥IjR1�}�6�at�j��V�����P��N��`w��t���P�ʿ�Ʌ����n�f�B�����bg�O���_�J�t%��[���R���x�ػ�q�����}_tM.��jh2K���ėe���}6��xp��L�q7�xЭ�f�x�#����&`oD�ۚ���Y]n�F�&1Sā_Z:��`���Y!���n�ǭ!�Y��'����Jׇ�R��Ҽ��ge���f7L"�.u���$������}������I��m�k��� ś��)v�����A��!� Tmɕ��ə�����+��,ꏓ�����%e}e�zo)�������Juvg py(����+�QVsS�d@`�g��io"i#��}(�XPk�;�U"t{��R���W_m(�ݽ����v�eх'm�b� t��qҜ�k�N(�K�t �`��=|�@~����J%ʁl+�Wj%�+�(�~��<o�6s��Nˑ�3 ��t��~�S	_-Z`ɻ��"��Y|ڄ���#�=���-���@����C�C�9�����2�qsȟh���o̾G�H׽V�n�� �5����V��H9..ߎ.����@�)z�?z��`5���ɡ��z麟#�$9�7��dJ���쓊���S�n�	�\H����D���Q��9�6L�jR�ν0o���s�es�8���{�7�Ǽ-H�"�@����c2ls�q��<���̣�C�y֚�.�Z� w��~�:V�iB�k�+�ř	��u����wq_�_��ij�R��d��6�_�q���b`W轿�Wb��}ŧ|��hm���H~QY4��Q��҄p?|�����W��m��<@�+�>v%_99�Z��uҘ�+2g�B�ā֨7x������p[s���2msю�,}����dQ�{��Z�`�E��Ϗ<���T�`����s�wR/Zeھ��1���]D�5D����=��B�(-���[��Y��=�����Gr����;Y��K,_9�C��[q��PQ��ܶɐZ0��q_޳�1�$����󛃡~�	����
�J"%���9D,G��Jǃo�?8hIHb��0�ha�s�&}?���}�n��Qz4�����G�]�X�*��@:�9���]��ځ�����iv���'�j����'���1P�d����	�K�+AUI��7�����}�t��5'0�r�%��7�'���M��5�^�8�l!���5,@?���������޲��f���f"4m��nŮ��VZ�
�R��K�uI��Q�bd�I��ݻٜ,�F�3�\��e��0x[L
����l@+�M'@%�����Sg��6X�Y41��'���h��s�O�����pL�@B+�\� ��z������ۍ4ȥ���������%ϴE�5{�'֯:��Ka�^0Y���/_&�a�n���aެc�~X� ���ʗV8!���R|o�״_+�.�7!�a�w���P��b�_B�*COK֬-��5��y�K�@ɑ�/L SEoJsY?��'B�r|ʔ�MB����՛%�?�<R��[Y��)���!+B�tk�2\)���~�1�r�����G���&_��[�7�n��]���
���%��s1b��A:е{�J���'��#���0�6>���#+Õ��Y��e^�AiZ)i��Q�A7�wTbc#ˁ�),ݭ^��6��@������jm�(!-=}_S�b��Y�����ϧyS�e�x#Ekང��Ox�X�繿���=uD��-��d�o�Zg/�Ĕ��Mu���mut�����e�潆�l*� ���N��ȵV�4<�����7i����b�$?u�i����c���Ƨ(���,x�6Yi*ΨL��Nȿ���%���b��rt�/��v�I}��b��fM��1Dv��J�~^����U8c�KtR�Nq޾���&8/Wu��W�~�/Q,I
�O�M�(ǎ��>�I����?=���h>�E�'ᩡ+"\����c�Բ����[�����U�՞����w�_���H��I�8�X�E_�r����eܟ@5���EÚ���w�>trAt&&&TTT�ד<����;'/eo����clp� �����U|��r�^�`�bo/���r��
����fX�{��B�Eg�\��QRQK�^�Q%����(A�[���v`߬ѓ�}�/�:�Z�M'�\�jX�-ʺ1׉Z�aP�	I������dZ�_�bēy�P�&����+o͓��`���2`�����*�jy�@/#��*����	���_���Fq��)72$�(����L��$h�h���*�}!.Z��4;�� g�tz���/=��b�ł��n(r��H��bC��i�k{�����xؗ$��Ό�����Zz1[RR�/�Ӊ����N��j<w?�76�����m}O�(iM�$c�4lv��xa:99]��u�nmm��T�Z�w������PL�	�ϕq�5gI�_7���m�}���ƴW���e��ܕ=��K���c����Cw�,�aq| ߧ�`���2�y��+��i�䜈t��t���t�&�� �~ɱ�Lw���I�'�(q�{-0�Ν�d����oWI��B��p��w�6GֆB~�<9�Ώ�C!�X��o�DҢ4��B�s������X�wAHC��{�v���+t�>��,Új���r&uglܺw']���G����\}��ި=!�&/� D>A���ߧJi�*U�a���/�8�D�ar�ÿA	_��K�<ل�P���K��
X�yNN������l�靏�+U�t���U]w���\�^*o�¿a��/z0�'8�Z%Қ-�%��y��2�߽�]-�ekC��Ȣ��ȗ��!�!$97���gg�H�e5E
_��tϵ�~���]f�-R������`��O7��e�ɥ�4�T���9�ס<�����Ofv���e>�fs���>�5�10o!��{��\1I�&ݸ�a�3�3����3M�I�������y}��*���4x��h��bg�5��y���!�鋼�P�����1*��ôP�z2Cզ�JԦ��$~l�䉳�k��z��s�M5P`9�����;���U��n,+��w��k?'%�����e�6��5�eS����i}�;���������-��B�@�-:�***��I�P�I�2�<�28��r�>F��M]�w.��k��Ƥ���+�'�T�Dh��l����UT�s��.�z�i�b�ҕZ�����9�;�:��\�N_|5>�AV�Qύ�?�{\�q�o��f��UD@bY�-͟v4=re�U��p����?��c-n`���A�[�/�7�l����DԮ��KJW�A�U����L�� =��U�����/�Uf�M�$�q���'�X�;!��u�.}���;g�.����Aŷ�:{�N�L�7�1�=�4�*��h��m�x7�,IÚ���7x��(_��O0�=;�xѴ���#��m���LV��Օ�_f�؇���o�!l�3�ey����ϴ<6��p�[�G����=������dct���%�vҩ]ME~�l�x��d&"H��6��f/�\�0O��"H�r��(����oN���qa;�Fe3�����فi3zΨS�Cam�c�[o;#�$)�;oK���{�rk� �E��B�_��.]%#�Ր����op�b������w���`F�XUz,d�d=Y�MA��U9,Y��
�i*����[��
?nE٣����l�&
Hgt�X���dzr?���YT�}5��$�,�jK�q� �X�0����9�յ
ʊ﵍�z��#,8������[�}A��M2��Rx������a����h��8�����t4+(-�N�q�TkQ6���t'I�(��V��u�o�۟@����	�����1���%IIII�38Jc:����6?��}������S��=�$��}���>% ��|{a��OK�ge�
�!ڃ��Q�:�pw�(��+�����6��6"�)��(�/��;�ے��urPn����D��)�Dn�����b��z��B�Sb�VDe2?u~�+���J����!����$\"\�Q���ř�ր^��j�B����Ʈ���ꃜb<�ޠ���XK�}E���Jc?�cW�}�$��#E�=��]ߛ�n��K�MK�"�	��nO�E6E�'���
���h�Oag��s��穤T�>�y�ƒ��JCkJH>�����$䭇�"��Ի��Yn�>�.�r�/8�V'
����;����3��[�t���w&F��[�?�/��e�öb.�ޤ�[��>�[�-�
� ���I��.���	M�,B-6_^o���L�#���kЙ$!#9oiE}��'.��-��g�$* P���m�z��  ���/�!~���ET��M�:������F�� �ae�@B�ٻn�/�Zo�ԏ����cL�M��Z�;M��P�/;LS�@�F�*q&N۫��S��s�߄��b�M�6��7�\_mG��?}���.ķ<��̌;b{�c|"E���%���1��	?w��k3���@:��}��v��[ca���rK���1Vq�3R�D3V!��y|8v_��q�pm(R��;�!'��_i�h�`Ӊ��u��6��!p���VVB|�
e�v"�\�Pw��>Q_U�4ɖ�����4#�����ᓖq��
&8��Y��4Uz�p	^�����U��*<�u�᜚e;t����C����
�����j�$�~�F��T*�+Z�֮�J��ܷ�N�o� N�ԏ��eY^�]�Ԛ~�ؘR���`ȜS5�/����FXklf�S�������Ӏ��Ml�/�Ы��>=��oMT��l����r�s6�Hh�(Y_�թ����"�?�5�h]m�?���\�Z����o�Ŗ�����*�lU���ϐ�W������,��� ��4��.7��)�)�1/�ƠUtQ�
����C*�#���=%�K�P�'G�,��/a�M�Y ����lj�~�l9&�l��MV��&5:�N�ѡ=_�}$��Nﴣ1���_��7��Y�F�x���|O�J��:�k;�R���������`;����66���>���`7˝O(^{��<�ۓ�����U�௓��*�B�^�q��9�����N����I73��u ��s���|"���NM�c�ۨN����/~�P����f6��ÛR�LC��A�Y��*����G�A�s�f�����e�G�䌱�h:�?����9�5c���5g���%�W_$d��N$c#2��h�
�DX\���;�>�rĚ>A��Uq����:���
�頝|� J����Paf�����'���*�*��c �ٜ�	�`>���f�F��憟Љ�����g��·J�����@��瞥�l���Y��dț�D�;�d	ݼ{���� ����o\��4^[�S���?Try--�4>�����ƵFAmm���{F�?��F�vvw˼2a/3eھ���'��.­?$�Ey�r��±�x2�_�;�]��Ѝ�/L�h�~��[�����f�z�>f0:ϩ��L�]���my^�a�s�,vg��}=�"±���A)&����#�jP���uv���Ez�p�Y���'��:[s/���.=�p�E��=
�q SRhQp38�3�I�͑SZ�q���%�9�h�Xô4�'��up*^�R=��"��r҄P��^W��h{�e/�F�b���Ks��*�o#�HRE�s{o7N=��~ؖ���I��	���‛-��������8QkzN��٭	��d6tz^v&�`ܹ��e~p@�X[1gX׿= �����ޞ���?����oq^�%f���V�լ�W�߿������]���������S���1��Qm���8�)�R�w
����wEw/�)��]�C�νg�/��/�w��=��y�0��1Z���u,������a3X�����:٨��O�^k��솒��y�����<�>���&�d�A�m�C5�nOş������J��T�B��CP�_-f�CvZ��'Ũ���I.[|P�Ķ1v�����d��#�#bC<� ��t�	ۓ*�<^�Z���M�ԌZ�����g�$檌'{����{�`�����D��,�k�?�F]M�eFw�.d'DC�I����@O?̠RG:+�T�
)���h��|�w9��}����h��u�umr����>�CJP��J[F���[}����Vp~��l�{��ٶ-�����]�!��Z�������_Ҧ5����/f�m|÷�u�� ��Q����A χzs�|��z�*�O�ը��,7R�����D�[М�`���\^�D�Ed�Zzѭ|����/}�����������i�8X,��>t٪Ǘ����4��%���m���	���Ĉ�]�8�$6G:xLXn�xPE[�J���b����Y�|2����Ss�Z#6���ݩ$�+ڕ%LW j]�0k���S�~-{����'f8�mE�f;UDw;�:�[��F��`3�N_$\3�@���Jwu����2��y0dc���p?�����,//�Ɗ��2��Ӂ?��l��5�[�뿔u���]f�T�, �OA��>���v�d��&@w��O1�C������WU�w2wJ�Jc�gTy�<gưEf��g���%��=T1�{ԑN��\,�9��B6r�Ǟ���q��ݷ�5�_���(1�V��W<E��ր�k8!c-a�h�	�oa��0R�nK��=�%>�M�w�f�lV��S�Y�]9�f�#�`����{�ScW��(��+֗vq'���у_c�\@^����h��"]2:16���
�F.�'1yr�HZ��;:�^��VOT-!O��JY�{��\�Q-XB��/6���	9�����m��[�6����<?Y����r���-m��Ym;.#����Ûy��f�|rjJ��C3���F��;<?�I&}1���)|ZT�	����X&����VA��=#b�W#�Q�;D�4�k�ċO�R�P䲼�:�6::�ҙ���`�&��bm�ɇ���VvW��v�7�Lȴ^´+��f�ؾ��C��]���G3�"��n�Z_�>�uu~�: �M�$�o�=ɆP-�ʙ�C��j�Q�C�Y��5;0��6�� �h�ƈƇ���xH
�t�����D��� �.1s�H/ �\~ρ�L�03KGܵō��xiGƦ3kU(��w�#wf�s�u}��\�)Z_$0ͬ�Ӿ��\"a�8�����mxv�̿�b���x�ҍ�Ņ�������k+���^��Uo��7�9��_E� ��`�������/��8;c#�>i�ֽAt��^�U�E���i����l	��6��=#Fsd$>�RS,�_I��gV��h��m͢]�G,1���z�!���l����lܮ���9�3�~��fn���z|�����&I��X�F��^3�Q�.��I���N�|R�c9=�i����V',�@� ����PG������n��g@��y�K��u�����8��z;3g3�����-�\��0����׹�k�;":��cv���b�D�Dp��(;-D�
l��]�0��ҰG��9�S��xƌ���r�ۭ&V )�c� ?)��U󲽜�IEbO�*���6v��������7_���������J�}��{��Q$<�2~�

�kO��зv�r�� �]���/A�Zo���{U<w2����=���E�@������%�Yh�����z�����B�x0�3�J'���:&~�ݥ؎c�������+�@z�p��f�Pn/��l���%fr��	����l��}���0;q���Ϛ4�e�Cx���Lc�LB4C5��c1Dv-�5��j#R2~�m���ɡ����?�;�4ֿ$�k��O�h��s�Y�����:Z�}���'�uGO��>��x���jmsh-G�]#��uz�+v����sO��ylw�ܨ���u=X�v{�5�B����H�������|qc;��?���tg=-dm����� �WPzŞ�{+[۾��o�K��U���	�"�*	�B�w�xb�����Ȱ�ȭb�Ö\q1'����b��9���Kو��XTn�@	�]n�w�L�;�Yg��q��1-&���ӗ���]��p^�S��kw�Bn�u:��\����F��]&Jt���׷���qWVr��ul$�u�d%��sI����Qb~kw㘗�Q�:��L�'�Pg�=��i@Z2�v�O�����ǏbL��	��m����w1SM�A�����G�ߩ�Z{|j	�p��"pm�|�}t���I��G3x}�C�V�T��QV�Ħ&��NX����
���������WB?|낕̎�E�J�v�Ը�M�3G�̓r���,}�j̽�a�Y+������uFGGk������wܶ�n<ݮ�93��l������]��f���kLGGw>�r'����v��#�/����:"7�K6g3�(l�6��s���OZQS�"*H/�c�Rk�nP�|�1�XK�-|Z�O�� �9X�Er�i/.����m`�~����7�|��y�el�I!�����A��웋�2�����cy�-�r(�o6��8a�Zқ��՚�M��ԛ#����Kc�},L�bs�ab�y8D��ƕ�r��%��r#���>�L���ݩ���gPt���s#��gvBpi�t��r,\z?����K�}�ݎ��Tk�DgH�ߠ
�2���ʫ�fbN�½����P���Ԯ���������mB���v���e2|��`���s�*���ƞZ���)`_�j��A�J=�Hʱ��&��ˣz��ëX����WNN�k�f=�%���B�=�`����k�����:�?����1~������쏡x����ZL+�-F䙗�c�=:��d��d)��^��sdt�Y���Q��]����ٲ�ak^O��G�Tp�PP;6���o>��@PB��C~��=���U>[C4��p-�+Щ���kl��|��$���~g�%��~�d�T�#��1hD����)�t�s��m@��*IY�9���\����cF��jS�7�]F^�tur��b��KS/����~b���c<�b���)2?ÿ�5�`0�M���zYR<H施6}���*�9>��ǲ���(v<��"�P�S�润k��C!�v�����FJv*2�"�R�^Tajcm��S�+l�U��}�/.z�jQ�#�_�M�+S��b�]�߰y����y�8���6ⵇ�hq��Nq{�tJ�>˗o���U+�e7��/2׷ �)d
�^W>�e���+ͼ�玦�l��S���<h��⯬���B7By�n���K�!]/�NV���t������@
T�frIgl�3�����>�Y3���!*&�Y��[���?��cf]�06�����9u�pf������� �Z�ԃ�^�Y8���1K
e>A����Lx&!�7�b5�E��KGh^.�ƍp<�{7յ�@+)�6tϲZ�=��h��"B�Y������qoX��WOk��щ ��!A�=D.X/����¬����3��!��z�Dwr��+w%��rqg�`�������-8��oQ��ɤἝ�>�`W4A���e��x�q��S�O�MT�LA�iY�� ji������Zy9���:%�Z�f+���w���������u�DSItEm��$���j��6����
$�rk
d�6�N{f˵'gg�\���1��8/)�/�V�W�%F6~�\X����rN�-]���b	褗��A�Tb�}PEM�]��A����g`X�Y5<�nCC�&���A�C�WA��V}?�z���%H�m��%$"���X��U����\A���|Ꜯ#B̒v�|Wzʠ޳�e��^S�� t�#�U��٧9R[��[��0D6�e�>d&��a�ha|�x\X�x��n��sb,��7��ǆs>;�U����)���+fC`\��V��B③a+~��=J<;�����p�u�6�F����E�>�����6�d-��� �α}���˴��4{	��y�)�)���IݼQ��B�l���ej��w��.M�6��ZS�΃n7AK��[Tv�@��2����ȶx\�|kp��tC�>x�6��Lɻ�kΨ�=�]"���v���"�5�
��#�T֤�5��HuW�ˆp�(����J��������B#`Ygҿ�y6,q����r=�j��M�b���w\F��ǋb1\�/V.:[vE��3.�*��*Cqy�F/�m""Y�����MY�����
�f�!
�y�Xu��,��ˋ>�V�o��z�=�	9~H������a�h��$Ѣ��p]�k�|�6��v���}ؒ��?a��J�`8x�c>L(���Ɯ�.
��9ݹ|���S=���5wM�U�5���PY���ExV(��/=����~�m�n1�$h/��0���I�c����B�c����.�ZZ���1'T~�3�*�5��V/�u�>fp��K��) �a�m��a�ƙ�&ۛ�68�a�`�ה��M����� �E�*`PC�ɒZh~���;)���`mԥ���H�\���qn%��4�>��y��S ��t�<
r��=�Bba9�?s�t�)����EO�0+>�F+�����n�����|�u��4��3a�௥�q>�1��c����Iݦ�>����F렙���lF�nn�F@�^�)v(
���T1��sv����i�����2=QGG�(�ޜ`ͯ�bg8�D //?_m���}!�|y�?=��薎[_���;������Ӓ8�m�8��!2!�d=f|T[s��VR?k�eӓ[1:��'�i�xqs�8��(8��7�\����F�\���L!iNO�=�s���VH�s�2��~�U�������(,�8:�݂�z�SO�s@a�����/b�e��~��tˣ��mi�i�K� ���,h��r�4���CTe���W���1�ќ���-:���4|�#��㳌�zZ��ŀ��#�0�_�dG�j�?EݼR��ѓ�����y�b�ع�"�h0�L�b����a|2Sr��|:y���>��������`��*����1�_�0Q�w����tކ���_g����P�ڱ�1e�X�&z�r����X��MS�]g�nW�曝�1W���� ��j��w�_��.�-###WۭuX���L����wd�d)��q�WZ���/���n!%ǣ�77��k���'����Sē@!���1��'j��j���+a`��;j�瞾�P��q�6����"��Q���r�Iq<K^��0uw��n ��
>1�Y�NvY1�R"�,�Y��zu�@S'3��
�/ܼ:�x�~V��J��[ƞR?�$[3�1|�@��Q}�{�Q��;M����V-�iq�����ؑ<mU�, �DHxcܻ�I���ϕ��ޗ?�Tvo�k�Q7O𡒟WO&7F�\�A�̳*4�j�ko�a���2�\��ۯy�b���t$h���Z3�=�sV1�x���f�x*i�[E\�ϲ�M@�;�CW��Ӻ��z���B� KΣ���_�Ɇi�P�I�o%�;pR?�]�5R�^z�uT��Bjj��k>�2���O��d7_�� Uo�$��Ap�
��	�\�v���Ԋ�Z���X��[�r����imKM�W�rMBY
����L��}�8��QX�U+�v��=j~��C�!68�ĸ�������vY§��^�������)���/>v�A2W(�,����>�tA�iv_����AxR�U&opL?;�p��M�5!K-_�Dk�8]����zr�b��G]�<�r�6��19.���~��q $c��FOE��peQa���iC�`[��N�>��}���n|��A�F�,\��of�����ӆWU������G��	�,�f�k��[���n����-���(E����
S^�-�
9�����B.��f��������Ɉ-�Y2]^T�rvd9^9�D�1�}�v�#\��;�$V�>;����j;���I�^�O=�� ��cc
�WE"���_hj�}��Jk��t�k�q���C���wGR$�6��?v\�n䄒�)**��\�	�2� �4�i��!/�ȿ?�Ujc�j2#�������Q�_�hj��W��'1T�d�;����A����y��y�PS]Y�\ۑ����+zk�+��+����R��|C����Ib���~�����(�Bw�Xyj�BTհ��ş�D����͒/B�!�E�C=��^q@��J�Œ?'��VYқjxEQa�F��7?J*��_%�ɉԆ��y�z#o�-������7���(��a�`��g���Rz+��W����l}5����u���0�E��{e{sȋ733I�),��e�kb1����A�U�����/�}�����@%�>%�c^6�bT������b��>�Vi��%���hRx"Щ
�Z�����q�}�x��)��v Y���I>���'d��S�X�pg(�8��u����~^�n�)33���?�6���rr�5~X"�U����K/;�7=�HX:|Q�(���U���qBN�:���w�+�RdWX�3?��'�Z���ua�?� X����Q�7=
.�hP�tH��E��nK|��� �H�
Y�Kq�&y�����^y���~����ѫ��A�A������
?<>(���m�c3)������
�'NzPMa)"¢���n$m9�/¯����}cm��4h���G���[�r!��~nN�[�a�͡cS��g��;��I!AZ��W�w�6B�950;��\��;�=ŝ۱r�z��~����y�xo���)�ԆQW�7X��N5�%t��HZBlؕu�+��\�<e�!��VY<8�{�+�5��ܙh�q�x���K^��Am��F(E_W�h��^���&�@����ci_�s�I����/��F,燅3͛{zɮf_��x����a�2 ��T�$8\�R's+�;;K�^���	l%�-> �U�;�j���0PxU��p�(Ѱ����7u��$�k���k�R���}�bB�L��������O&�sx%����R�^�b�#��(��x�{L�k����/�>�BN�[��w�z�'kvWB�+x���Бm&�z�L�,���<�hI#����ŋ��c9���
Z��c'V���oS�93b� �B�ho�hٵ2�4+`"�<%�V��B��P�M�C^��B�{��6�ЦE9<��X*���/v> ���A�3�|�YKm!�J�
y�o0�'�95=`�����}n��PL�d����/���2�'ÒN��sٻ�bn~�p�5o�ג8z�\��� �EQ!U��Q��K��]F��O����f����3��G�	����� [y��g�_?/��xu���x�wJ�R�z�?I�)���UhRps,e�Rc�S��)1u�8Bmĸ�ټ����Ä�&m�nOs�&R9�C�hQ�&�>a��v���_M���ry��{��.x`iw��ls�w��W�|���ؙT���{.p4�.�[�����s�'c�����Ly�'�8�{]=tT�b5�k��l�n��)��G�xŴ��a���8k6�]���cz]�o�h)���v�Dz[oTVD�j��5Q(�-8�o�ں$��)Eˢ�턎������&\@�Gqa�/a*�N�#Z8��c��]���ʩ��Nz&���)���K�.�z������� �����1�RQQA�+��1*�����gR����A���;����ۭ~�g��a���3��{p��B��+�y#���BK/Y��ͥQ��p��"{���!5��0�2�4|4$,�-�Mâp�|Sp���(�Y2�>Uk��P��]�ݝ�%�_I�qL�c����R�w-�2��?0��o����W'*J�Z��cM`�H�(�
>otlm�V���[$�$uM��T*���ě��$�՚���n�����[1b��F��&c���d���oȄf�7��ʦ�x�;:�EI��ѓ�j�Ӽ&e#�7}�<���wg�Wh���;k%�ύٝ�=vw��3K�h�k�81<r��0�\('�Gɻ�Ab��Ko�3a�9�r�P;Iu�9�BT���#j�V;��B�S"�k��uL�}&O��~�?��s�&_o�5��m$�&��hr��v���b�8pMu5�+����|<���?�JD���75e�ե7��y/95�ʙ����ֻ<���}��в���bC�_՟��g�\���#�o�&&9rKgHj�qo#Ҡ;`��c�0��Z�T�����D���,"��ē��>�g+���n�	��QՇ���BDwS�R��p�H�> �����v#�{����[/ªKO��<&ˢ��:��p*Vy�k]V�~��Q�`��3�U&M����j�0�v��9��$b�8q�`��X2�6lL��FsU_t�Z�R[U�g�8�Q�	0PQ����P=~kR�[���+#�N���OY_�z�f�=WQ���6ml<K���ey�����K����D:Y���è+><O��h��~W��%����>f3���\���k7�4T����>����a�E�ٱ,���gB������.�-��]��X���'%��I,������q��c�|���{�$�7\o���]�j��ɤO�� �4:�ǆ_��.�=�%O`Y[Qs�J��J���攕����AB�L0�
H��Mа�4�T�G�W��С!EcK�,<� ������N�y���oZF��9��IRqµ���c$A�E����^Bg��b�U|�ZpNI���}�Ksr��j�P���5gn"����_s�Y���}Q��1��D&�gm�gjI�}���ؕA�zsE�Xѕ_`N����8m2�g$?@w%��X��Mvdg=�w�lKQg�� ��%9��C?7_���I��-qJ�C�Xj�~;'O��/�W�n�O��l�5�C��D=dEA�k�l�v�����E�B{���H�\�?~�*���"���n^�Nb����6���.����z��+���5h�o�����W=ł�JD�ՎGdff��lQ�>P���'t����B_SJrKE0��}Q%��^^�T�5�5u�W�UrC�������p̢0>슏|Hߏ��^�����q���Ý���Xn �݂��%��ZF.���.�=�wR��[�<k�^Y��=��[���^k��ph�2�{[�8Wo�q�K��fl��P9�Ԩ<S����U]ƫV���@��!�8�ĘE<d��w(s|�/�;x�d���n��U٦>�T!���R�lƁ�q_V�l/��qTB���O6�ؽ��L�nU�^p�?�u��	�LZ�\n��P���yY����J�9��$#[N{�i���<�� uE�$�PeL��ӆ�}"򞅤�.9�g�ڸ��Y7�$\��n��g'��yB����B�b=�0Wa%3���	E{�b����_#�[1"�G"0&����s�,�c�g�	/C��X���&���y�&�D�{�V�_�2{��_�VlR���}3�C�P�s+�za�6�	�G{��V7]:^�4��#Å��D��{5� �ʄ'T_bHqB�����h��#.k��JY�����������������?|ĢT�q�Y�Y��{�Y�̬�T�.����*�g'#�Ã�`)ʳ�9�P&hw�%�����}�L6�w��]�ID����Ҡ���ZVғ�*�/��r�ݞ�s��T��E��#��;L�4p����50k�إ������!C�dQ^�a�?� ��S��f��6xX��$�sz���ɭ��)9H���>&�fTK��h޼$K����;27�m?���s�Jִ�d3�`��E�W@&�^�A�8;b��$�I�������~��Fxµ�_��c�;��8*O�K������Я"�p��UH�=~�l�U���K5!�q�>S�v���jpN�I���,ڊ��]�՜l�n<�ϻ�Ӎj(=�9]�p)l)���\i"��Տ��-�H��w��`���ZgC�_:X��Cu��L��!^"4џ�/U�Ju3��˵�Zwq6�c׌��?���,n�3Q:!��t�)<?#鷥W{Z��+9@���M���<���_ް�?5��i~_�W̏�?����q���H��8�n�k��(+8�
�V!<�ŵv��3{�$�+���ր�v}���$�x��]�����1��J%��>�HL �լ�^�0�E:]����Vp�--X�����4=�,�?��֮�y��{��~;S�K�N��`��ER��wz�(Bcm�O��D�]��]�ZJ�8[�������4y �sq�M���|��Ō���o����(�b����L_�H��{Pn�~�W|Q���.;�B���"�E<���4�=��w2e�*@�`�0�'{�!�3�t��ki/�'z�N���?�)���&|d��A���ܾ�L��8%Q0ti����5�5N3'r� �Lf�Q�`������L����R�_��$���y�E�����?Ʉ���\�J��O���"�Eíp�ȵ;b�|�U�	t�Շ�hw�!ֆ�׶�o㥗�B#� �p*ڌ��{����)�Q�{1Pu����R���9I��q=�g�3��4C�ckVh�2����2���C�i]�����?rn�|�3a޸����͕e�e�	lcdg���i9b��f:���I!SP����~�ӞB�vc�kYz+k+���z�>>>����@!���xe���4B;D�"6T�E�N�U2���U��C��<�{e�l֩J�h|v��g�L�~E겿���>>$�T�)��y��u�l[�<��f����^�"�~���]��:N8�3��r�_�^E0�v����d����ѣyHVh���e�8I�b|tkݨY��j���gϪ��*R��0�"]t�;G�E�#�>U<��|c���;77��{�L���(��7�,�]�Jf�?7�;�M	��w�;BGr�3m��1v�.ܽyL��9k>ܠ�(����O1����f����]�d�C�xg��� ��扠ѕҪV7�����Z��'�����5� �i�~��/�������v�	�+7�T~��&G(z�YJ���"���y�嘀�Sl-x�c��T��l����&>ׇ`�t���n`���eZȎ~������ D�ү s5���L9y��8���5�̔E��߃��+9�Zo$2Ђ�%��u�$���
�3�ӟ�����ۡ��d��VRD-)8Ṵ[F�᢭��ߏ�
�k������v�,��L1����:�z2���5Va�f�8lF�J1	����d�[��MSq
�y�z6�x؆��*�{�_6�}���Ղܡd<�u	[.@�;���c��x���ƍ�dY�|�������)���ћ�Z���-)��,7�#*j��j�d��8ݢ��g9MD�[�mK�VO�� 3�ls�~hx�o���I��m٩Vț	<x���q-��2p�$��!��W���B2�cO��������?���j��&�}�a�:���f"nkg���*�'3�/�E�t���I���p���̀�����~vv*�Y;����|l������	!ږ$k5�;@��(,[��14����J������:�(�M�)G�#�АV�B���8���	oE���y�\����g�Sq"j|JG�	�@3RYo�:�g	fEUeO�)OW�ʃkʱ�DS��Њ�����Ӑ�GG �%WER>���^/�pK��h�LWfY�e�%���?�b����-}���A�a�����zAe�h����! 6��ݍ`s�s��Ƕ�̦�����n�Y��p^<�B��'6�:7yt�)α�GGq��}ٶf��z���fg�*��!%����X��/:̾�R���̢��f�t0��r�V�����&�I�:����z�dN�0.>&_g���O{)��c�Ip�l�ަ�B�1T��R9~���8:�'T��wf�,o��F�M�߫��'��A�֩�tl,���1��{MGnn, y^^�`����#}�׏�`��y����l�.W�khJF48l�����\\�?.�b9o����A�;�����	8n�^�����j��)�4/��R�^��Xji���U�	H�y��>����,P(S�����><��{e��}���wv��N�6���f�5�ݮ���O!�}B�)s o�R�o���n�o��i�]��JM�
����Y����U���'�`۱��gqO�u�m%��>���5�Z�� EC`x�v���ό2䴱����:��{�h�d�ٰ,?��)`��r	����A�G��em���#�\<N��#�<?Cl=~=���4� �uDy�s�}|&����1�l�W���Z���'��/槣��[�@k���5eqV��u�b���O��բh�w�����&�:����j��+đIغ"d<M�/�c�!��P���:l2DN:��,�j�L���v��|o9)��T5C��������i�y��4Ij����v����x% �Y���sf�ݵd�Ð��Ѯ����`��Sl���{N׍���PR~'�F���C����cC�W!Hh-Q�~����x����`��鬾n,��ťF��P��<ֆ,B,��E���ڗ/��8�k��{��1W@��F�X�Z{��������4��l����[�Z9��X�~M�b^�}-��<��'�;�7�:��O�<��k}��B8��m:%e�����\��Qj���o��� 5łw4��f����4�P�}��|���]��GT��{1Le%��X��X<UNx�5���!A����/����(J��y����|�"�5�2鸆�n]���$/�s54�o�Z{��ۺ�.���G�o�Y�c�X[-�\��py��ZX��c �0�mR���o�`ܦ�ϻA5I��u��9lOj��O��v$���/ݑ0�g��1���!v.��������k�h4��p������L�(�L�]Q��CE��}M��k(�=�cwX�n��:���}W\�_I�,���R����Mm��I�v�&��@8�Ҟ:�`�&27k�>H:6�XB̈́>Q�ZE�lգ-W"��|��Պ�x��&�Q������G����vޙO�鈙��ښ�%p�%�I�p�~�}��<ex�����-���ک����	;S'���s�C2��S���@�����]�։:Y���^�;�A�<��s@oݝ�����@2�g�4���\����]��]u�kL��l�v^�A"8{P��1��R�⣰�|w�_���/ޜ;e�{�f�1E�v1{U�Yp���Ô����ddLR��{[�t�3�\�Y���)�*%�����O^ݠ���X*�F6���	R���5±2�e )�LJnM��3{�+�6O"_�xj���zs��{��Q��t�7׌���^��oq:�ͼq��W�E�~���O\ތ�ǂ�����-����6���d�PV�%� z�z3�1�b�����	�kk+��~�-w^��2a�?��wE���v�"�����(G�4c�I=i2~���d4���1K�l��Xk�m˱q���ON�xh�2O0�_C�?U���bw�k\e٠�����o����'�
r]R��dx���bA�
VO��G2����N	���� ��ss3�=r�V$Q?���w���/��W�c&!���;�eFjFB_b��P\�K4�z~P��w�^����;�	,k��M�0�m�B�0���-�e����I��4"�b����xu��֮b�~T;B�o�n��F������3^��]��ݛ'�ڿ4�ԓF�≙n�oYF�lH_��r�nrp��՟N7S�Y�!..e�Y��_��Ζ��[w;>1���%�%@!I��ve�B�9P���}ߠ���Kn�L�3�=��FԸ����=o|W����[�Ҧ2���g�_�t6�@� "B�K�����y�����{��{��M��m߈�ea`7њ$TOL ��5|����}���B�:�Z�.y�a�t�>"�ʕ��
��>>Rͥ��XS�߬r0=��И�T������[)V�j_��o$z�Q���q�����oH� '<fF���d�w4�V�CŐx�qJ_;|oV?��y�\yo�λ����@���L¿��+$��tZX�����d�CZ�u�3h���*W;Q���T<@�4�o�z�M��VU�`ef�q��
��'v�X����.r��z�A}�.W*\�c��Ј��۶�(:�Y�v����h��;�_��ɆN8)0���d/
�thyt<�O^ؔ]Ԡ�so��m(htU�J�*j�T�%��K�YQ�T��E+n�/�V�Xq�]}�f�)���� H���5~�xh�4	�ǧ�h0�ģ�8�P���Jf�T
�J�Α�Gk>gpdC�����	ŕ9����G�u̾�<-OHBB�g�v�V �pӲ����5�'�歕�E����i���-,�v�*��qm�Vc)��YF��u*�Pjݷ��&�V��(�()�%���(x���iF���Wʷ�߶Q%���N�Q�۰)V�]�9j�O�%��R�Y�=~��2��)r����"����B�72l|���s^���\<�{HZ��&TZ8 ?�H����v���6��}�#w�i� &pO��,-�ߦB\��;A܊��k/l,y��'��:Y���[2��Tq�<�7�=�e1�0k�뛲vBd/bT/�ǮV}!��O�uԏN������yp�rձ�$�=�r> ��3��ȼ���Hjw��h%t�G�vt��KLo>N^�L�����8���{�a0�L�+#Kp�;b��a��sU��Φ���7tP�����Wm���Uj�� �?O¤)Mg�9,�4��F'�u��[\���0TS�/W�O���a[�0ػ(�z��|��\�Ŵ���5�(���`��r����ژ[!z�����bp,��zI�P�J1qLM���r��u�귣�Yw�Φ��1�yO��  �.x��g���A��q2�o�u��&������B���=̷������#�+�+�S�wK�t�{�e������b=ac�	323��/� �S)��нt���{��y�1I]!8.��^Tc�<E�)��|�ꊻaz�5.vP�A��cp��L����g;.�tܶw�?�mL��v�R�����:�����{�����$v����Q䢪�;-�v��Fz�%��|��Of��.�V%�V�/���0t��P��*^��h_+*'T�8ˏ�qu��.����x1_ΨW�8�߳HA|�x\��mĜ�Ɋ����fW�.GGk/�g��8�j��{I�~@"�d߱�C���.$ҹ��q{���bZN�;�/쉼x�8�r�Z��%����YS��V�����&��<v܏����Zt���ܷ[��	�DPk$n
��D��.�� z3��Y��%���J)h��֣�K�K�ŋhy�n^�������|�c����w�2՟K�g!�f��ЧD8�;��be�����I���x�����CO�2�|��^�Ѧti^��a.A6�2�:��US���^ɖ ��S�hG����龜��O�/�~����Pb1��I��8^���z³Iwß���-�l2S��.�$�$�)����6�����n��R2��'n�;�z[_y~/�<��Ėe�=��׻h��/���yf+a�O�\�U�+L�P��T�
ʻ�?FYHkwk�m��It�g[������t�!is��R����M�<��[}�3�Y�O<�;�����X��C��7��KK����c۶��fcӐ�L�Դ��~Y� �/%���Y�-�v�]q3������z��/���^��	A�4���;v��owq=q`�aht^�n�gygɀ�qٹ����'�&�����ީb�H؋K�ÚG-�
־�1${Yi�Oe���Y�^38&Ѣ���zVń���=�{�t���fS�iT�hO~�H�e���J�aQ<�*	u�}ы��O��4���	$*�3��]��M棌�'�tj}�3ro�ɊG�ݩ�I!}�b;�֌�,�?��S.�X���B^Hg �ubZ��QC�4V����
�,P��q�i��d0�nh�����}���GU<�MB�^i6��%B5/��9�Y�����^��.����}<[����q�A:&D�m5�cJ1޾�V�6B�I� �P��;fc#ҥUOL��/����2Ƣ��ǋ��:��p}��5��SS�#������q�ˑ y���Vȿ���G���nY]L���#%~F��+�C�0�n���'�j�S$��Q��C��*6�^�}�0D�3��۫WP�6�ar/���}�f�$���%����	~L@�ג�B�Ĉ���;�;�[����w��E�"�D�ѣw!"���{�=z'��[��F/c�}��������-���Y{���>�L�z�	ŭ{6��.?��R͐f3j�(�4�\�����XtP
2������q+30p�"R���,=��R����LѮ�ZY�T��ʿV.{��8Y���_������d�n=��[�f\��ֿ�l� ��צ���Ƒ�9�ƽ2�h�NW���ȹ���n��JW�,>)<oǛ?�{m��feK<+cb�nB�_�38���m1,�Y~��Gn�a�{KⰐRF�'曞������3v�'���&�JmseS?����r��ɏU��Ķp}/&d�[JԸ#[�=5�dzWfF�=>��42(���ڨUd��9�����ӻD�M�K��ۂ$C�he�N�g�L�`U�=�ȏ���끠�ga��~�EY�E�݊���`���ۯ��t[�����d\ĉtoe��K��/=�B^n�7��� O4�O�Nh`{����B������%Ո�3��J�Q��La��Jg��o�L���|M/�}�\�G5����NNƒ�� ���t�*�|U�μ�1;&�uM���Vs�l�g����N5����1`���B�z4 <8^��\$o,.�z���wk&��z�'�_�[���P�z�R{�<����u���[n��U��ˏGl�v����I}�i�y�t^g�lp�Jz,��Ĩ�����Ϟ5��=�nsv��|���x�CJ7�Z�%$�"�ȁU5��4T�g����@��[�H��p�PH( ]�!0�E#�l���eY9�b����m���WX�ԩ� n�������7�z]�#4v����~��4Tuass�ig|VE˟Dl�_���n�����]�r\��n�����t<���BC;7pGS�4���|݈�S�N�HĂ#�#68�)�ڐWSE�E���b�J��K������c ��
��������6��d��H�9�B�Ĩ-�q��.���tI��kf"2l�te�G�A���"��i�Uj����29�V0�+C���!��&���&R�gMLLp!|H��D�68<.��z�iCd����Q��Y�h?�/o�n�9��{��$��(L ���3b�\֢7\Hf���ڦvE��e8��G<�� y�ҋ�ǻ��SX�eH�d-IA��yeͬ��2,����#WS">C�v�Uho;�}H�bUC�T	�e�h�拴��Ԛ�.փJ�U�4�o�+u�=�pk��@�^�%n�)c�5�pl�n�"(�n@�%���sj�(,�tu\)���
��[i�����������3��y�j�W�b
�P��op�8�m�"�r���v0�*����T��?�p��\���|�}��P=O���c�����D���^1+f�����}�?�v���4������ٵ��}ruРi�BE�cD���rSx�db�k%zsY[i���^��6õ��4KϠ���V��sł�ym4��D��v���H�T,��E�(�V�4�Z��ش46���s�~3F�,k*��^s< ��'�&!!��keOeUdx���eW��\�rQ�]I�?=y�?��b��o	
n/��t�fT���7^{��T�T�jN�Q'�4@��q�����`rH�1�_f�����Lv*3�- 0�឵)�q�@��֓\�1��q��ZV�M�����eVsᔑÔ��՚��X�v�DĜ�y��gdv�n?�*�I��d|�vv�~9�lXx�s@L���ͤ'9$�M�5��Hз�])U��uA�6#���Mo$q��,�;��sʇ�.�ί�ƀ��O_7��`��6����@�h�6��g���[��T#��>��x�]�vx#
���߼@w�K�Wgu��7��K�vu(*�f�_�7�o��?`�b�%m��%�C�W_��-^�gs���胏t�-u���o��rB��T��sƋ�qUʋ�}����Y�����e�O�@��H,3�՘o9�����Q����+jM���=��v¸U�V�N#�O1E�qw�w����}�	��-=<���r��n+6I���^�s���W��I���&��H�lOd�?���Y�9R)*`�艸�b�*��P�=�i��l�LN���B��I�)�YM��[�]�I�-����ڦq�Ux�e�z�|�'+%p��P������4����\��oД��lLc�Ot1(��CI�X,`�x]�.�ۺ�?��+	��4�?����TE���s勵�0d�D�[r�`�����o=tv!�Jm�Z�~�~gE*婏5��j>�|
�]yj;ln�_`8Ϙ��;����n�F"�W�t��(�-i�1��l�jBU?Ł��l��3t�}_���h�*�����R�$��ɐ�-�z��+4����|H?���mD��n-���Ǣ�%����31*���6�vb;�kb�Lۈ�-�����e�������\_Z�촗�c[��I	�����&K��@���C�3�\_�i��dҜ����:[m��uI���50�6v�( y.�h�rٵ��A����ӥG w�	��I��V�_u��|��  ���h��(ea�#�C�ɱ��)C��F�Tz��Һ����ֽ@�h����
�'~�/e*{k?ҡ2�B���S/[@=��~܏~��2)�^������4c��,Z���#M&�d�ճ��A��HNw(��c��J"�}��r�����A�FC[[�j1�`�F-g;�8����?Ɂ=�_��nZ�����҅$�F����r��d(?�Y��ډn�֩gA��ԇ�䷌�;=�J��S�'���:v���0-JSo����~���������������I9�2�cC�u��G:q�}n�Is�nO�l����5�J#�Ȅ��F|8gɇs>\�*�~>��&p]klo�"����I�Gƺ]�q=�ʃ�����vC�D���s��Ƶ� $ �S�� ����B�B'�bj32P��F)�eD�ì�g-�wv���>F7�U��G �Y-zn6�<����0��[��#{�>���Z/V�A���o�B�:�Z��鿹��R՘���:�)�m�P����5�����O��5�����^��I���a�,��VJ8ո��
�b��J,(�y�������J�V�����ż��6�)F��H߄��4x��J�$��?��o�y�(=m���f`�^w�>:���b�BwD|~ ��A]P_���, y����V9SkGA/������0�Ӽ���È�Qw�+>P澠��� �8]�U��x���T�L�����i�oX�N-����������`�.��0���k[���'��O���.=�~5��������=�md���Q�U-��y�_�ʵ�h
BJ�6�=n)D�G�Yq7		�ns�}y$�I994�x��)e" ݝ����q�����ɱ�ѭA�#���gjb�uE�M���ۺ.�dBP�#�[��S�:����h�fO9;�$�w�]&No�ѹs�:�9�?�j3�I���[Ѽ�����C������&w|���X��4�w�ݳ�i{%WIwoN����[��}n	�?
�Xl��iOt�4�>�{_���f��؜��������24��a�5���|��e2����pL���!�)9ws~�M$QJ�VO<�@���q#�d�'=��X��bΚN��Y5H�����I1F~Ό�x�K��Y��-sX�8�KD[\p�G�X?�i��NH�/��uH�ʿp5*���{k����ZZ�l2"�Q��s��$��|�g&~x^�W��5���SXID��]6��7��� ��㒹�D	>�P_�|Z�0�|��^���E�8u��X�]@k@v\�l�ȗ�:����U u�2�Xw_9ġk6N
S��`��Ñ7�wwv�l�S�k�'��3³�s�k����+g{p���qk�N�ұ|���B����U���f&��蝧�~Qق��p�&�&h�p�
ם"]�����0��!f��'��d���5����Qː!�՞���9c��'OwQ<:�:o���z����ٹ�(9� h���K�ګ/~k��%c_H��+�?�\L$��%�Ӹ�`֍-mb�"#.3��f��;��ll-�Pb���~!�>�3���È3o&\�㗸V�X�-�o���eLvr��.F � ��IO������B2�7ݡ���";��|���z��
l7��򚵂6p���}���V��?)��D< b�\��:}4ҨdN?��	�*���L�K~��h�o��	61.v�4 ��� X"Q[��n}��K�:�?��^��zR�\��D����6O^B�AM5U�)�,P��)�T�Q�劜�NJ�n�Ϡ��`i��������4/���啨��]z��a��� D
�;��IQ�P�a��%h\��Iۈ�o��� �4�n=���y9x��kva�u�M�� �Q�އw����+�r��X����e�l�:�`���~�a��AV���	H6�he.@���>stw�^���o#FE��K+a����;�&�_HW�[�ܪ*�����2"�W�P&	LT2/�/kg�N����L������H�������D��T4�v,)��B��Ue<�+=�����޹��%��^HMd`d��S�0�?�ʂ6��h��y��T��ʝtk������uQ�c�v`$�-ٟ�O`�fP	)���(���Y�|)������!"�dp�F5>���]� �m�K��߄'ʰ�v�����a5P����`O5����/ҷs�S5��M�r;d�+6H�(���v�0Qx�]3v*]�Ov��SUX���+�En���c�%B���}Vh�rb��ڭ<�' �T���⁛�ҵw�AF�M=g߳7�.��y���D\�}*A�##������/��O�V����-��z�E�E)9��m1�+�1��`�v�F7������+�Mcc.�,N�rDY��
:��5Ʀ���8�x�,�7�̒�9�|���,�OǍ�EEE뼳�+�m9( ���-<��Tm�`6�~�:sN	�Q��ڵe���r�Ly��pm�c)�E>�lr?'�=�o4_��H��a�ʜ��l#�)�*d �7ӵ�Y)e�Z�v_p�i:�rH"�.kH��~���]1WX�|g��NI�	�̢w��S�Wr���oc'e)�x�[�*;B�6�,�y���DH��mIm���#�{������T�k���T�>'��Y�4�{��15PۤE��ҷ�~_�������Q�+Sg��fS�L!U-OC����1�D2(曢�L��7�����iL��u?<��i��6�R���:�hJ�Jګ�0^���AH�6�
�C�`JCkHx^t�Z��OM�b���Ѭm�C}�/ck5F[���3�t+�<��}
[�5��Wn���_��ZO0��H$��W�l]爹p������b�񢹟msmV�n,ck}�,c��ײ�<���Q"�O���ta�"�c|�/��(�D���Ϟ"z��x9�[�o�!�iu�wXX-��Ӑ�����e�k�oCεr���{������dܳ�?���B��P�sT'�:i[zQ0�տs�\��*e��9J�A֦N���GY9�S/R�>h���w��qx�j�M�dC�
�n�������qe�$|S�Y�5���_�So��	6}��{5��䰖�br�ӝZ��?� �_FD�3g׾�]4瘜�Cש,mE]DR&��8%-��j�܊�m�����sp��CW,
5�J�Z�)'�ͭ~tP�/�k��;Bޝ�����-�)+�z��T�����-Z5����#/M��K�JWf`������g�z��K���_췮K~���4�i�9ih�������# ������8���ZK��#}���}��CB�>O�v!(|�(e
�@Шe}[��)�y}ޤϠ�"�?�d�\��Ǭ�)�'�p[_z�@�X����;5|+��ʜU�W��y�M���'�e0��{�>�j�(�?v���&����֪E�R�R}���T@�t��R�B����e2.%J��A�2��,�XJ��,�Z�.�o4MR2�������R�!���G��]��M�Wj=�Jl���6�]$�7}�'H�4bԖXR�[a�X{Nh:	L���AW�4G�4x{xE/fS���Z�ڣ��ipØwPYڮ�*~���l�M��c$~�D�XO�;ZKÄ�9&���z�J��q�	_��.܉h���0���а�j��-"A�!vqܹ�q�P}��|�+�<�s#�_M�}
>�9nɉ�2�^4�Q���,g�G�����H�ո����.x~8�o?�k��4�JE�
�R�2>'���u������0?��$| ��R�_2a�BU0������.vZ/�u}Єe8@�O���O;k��G��?=�}�w��	�h3ř�w>�	h1�KC���4�7��-��q|t1�!���w��[u�����ཟ�%������2f��(�{��b'X��N�˵�-�x�b+c̸��H��,�\t�6P/>.��W�kf�>�3���|\s$��g�g:(�0v$I���@Ov��5I%TfՆ�Oz���^���xws@�'�|���e�W�B���P���X�� ��$���]s��?SUIJ�.1��%���X�,Z�\���x �y(��F�`�WVz�|W�Ÿy�7+�/9�n��j)i>��t�݄h�w�TZ~Ͻ��Ѧ�w���?�Ȍ��ޚ�i�&�-Ɯ}�'�ݠ}Y~+��z%k����_��B+�I�R�+	|ph	�9�䋌C�l�@�N^�\>�X�p8�o�z��D@�ƝT��T�������0�`!u4rβekC�6�P��w�	�L���ս͸���Ƞ%��y-�OB� ��`�ѡ�-��n��2��v�V�克��xc��ϔ��=S�?\��B���61��V�zvQ�q¹x��oL����tG�I��-^r�����F��H�e�G+N��Vw!I�YzϷ��76���S���� �(DQ<_�圁��Ӌ�bf�P[�D:Y� Qo;;���FcR>�һ�
�njA��f�fK3S���84t�>s+���$�<�������w*�n8/�~��b� _���K`�*T��=+D��$�tm�HC���x�\�;��F���~ya�B�,����-v��Y/�r��z	��{�9��׈E���q�Df�=���B�Ɛ ;Na��B0����kA;	\��?Xm�]>�� �2<�]��ą���c�LI���H��ľ^�����r!a��W�.��$k�8��AiY����x��d�.�TDeV�!�����율�o��S!;�� �_�|ꆚeJ
�+�ѱZ9l�_x�b�����S}'��<�����B�H|��u�G9�����;��X�?]�*���jy�'Z#��s��F|MzS���y,�.�j�Ԩ�r��C>'��Yb��0���ۏ�闏�/�����~�
Z�J���+|���������	!f�J��q��=[�.��#���!�����A�|�> �8��C��f2�gZU��$W���-�7U�.[S��з�k�N��t�����" lkT=����cM����~� ���AHh_���F��,��ZzN����c���ٚ�:���_�ݖC���xX/QG���������n��EE�����F�ꑿ�:�'��I��+:��.�|��=�����/��Z �h|���ى,���|�Z��7��7Ue�}��4�<��N��}�z��_���E���9d8� ݍХM2x���#&W,������Ai�?>�Q�ώ�=��&6���
�V�._��_b4v���d��k��5��S�"�޹{�d߀ف��d�
`��)Fj�i~zr4Ƹ
�1�ݷSƙ(������O�Bd�s��nB�c��"�X�O�lTE{���+i�*IV�\�����_�7�ͧ!�� ϸh�/n�X���͗G��u���Z:!2{��Ih�@���A��������D�o�vç��� �6.c��?q�'�Xtp>����Zε�(��M�X��J��V�QZ����r��&%X�)ɕĸ3f��~�/����������d�N��wך �y�+;*vb�r�2�M	�|v��Q�|����R�^p?Y-�P�6F��JY���!~\Ր6�>HÕ`��l���4uJ���Fv�'�r'5���nz�a�O�ō��R[��������W�L�3�ZV#8R�$�ָh�j�T���:�q���{Թ�y�r���K���_3���礦vLh��y��Vt��.SJ�� �4��"�DЅ��a?���2LJVS��W'V�p|�z~oA/4A�S$J)��h��.0V�Yh䊟�Wq�dO�F;��8W:�a��=/�`���\s秢,�fW�v�	�e�{��@19�ZE�Jc���Q�i<xV���띶wvQl����/�^����\Hy�@^��V�Q���j߼W��㧳�M���V�oSh��T�/#\ͼ˘Z�E����c\}�׈h�����ݻ��UN��0��Y��� ��Xl疷q�X��o��;�	��s� +RtǠő;�D�z�(�hs��b$&i���XY$����T��}��ئ6��O�Μg0M�5�}$��N.���0��ߘ!�j�)G�������������j�ڶ�LeMW�E�ܾ��鍾TP��f+��;I����E�>�Є���-�E�a�������W<��gs:t�-�%r@[4g����' ��ʙQ�qk�'k��Wj��������b�m"Z�j�b������f�p_���{.�	]5�v$ǣZuv u�)�-�*~�����ܚ韜v�'W�M�w�4_���d#Vl ���B-d�-��6A�}���n�������ߢ�)㼖�Q�k��}�^WEQ���h��c� '���Á�6�j�����~Z�+rN�Y�W�Qywv��-��w�)� �֗^7��3j�C����52 �^!5�
qG�	����������{M�3�²�7S�K�$E,U�Γ��{�0EHn������N,�W���c>�~�my�Uل��7UvZT1��у����jRy�9� � ����0��ΦCZ+X��B�\.�+/�k�E\�$/;��Sq�_A��O�h����f�tX�bmYo,�Cx�qgj��+f�</��p�ĘZȧ3����h#���Yw���gZ<�q�����)���Os*�g�)������֜���5�ף�P☰R-'�h��7�d���s#�؊z���)�u��1`���k7#w����g}��K�f�Q�'M�3c�b+MՅ�H���.�R��o��3�����0��V~�7aK0#�P!��Jd6�$cPj�ġ�P"ɩz����?���{�+�E0�z���a{�-�!�pI��Q<�%�?�m��U��+("�+�����|6��"�����:�����U�9\�6��ߦ��b=l�t�a�ә����8E��\1��#�$0vp>m/��~[{m�I�d���g,ݝ�}���p���ݭ��U~����vۯ��H)��;ۦ��[��F�+�k���:v��N��2-Rƛ�����+�j8�ό����Zdה�G���>��0�Z�'�ɝup��V��{�$�B�?�ep~rx�,cb1jюr��W!#{��=�jd��xM�,{B?~��D�tFW���g���co~���m�vmp_���Ђ�u|�o{�^	_���4 ��m���l'�2..�Z�U���W<{������y�Y�-c�oa�Y���q1�j]z�#��.��ƙνJ(�͟,!Ͼ�[��>�:SDW�h&���<�^���X����/����r�̡0>�������Dم�ڃ�=[ �<k�?$wS߾�Ly<�\�t_�>�#�}����gC�4���ю�,B-l���� ���MG���)�D��9��?�-S/X<��n��& �S|ۺ��6�����
433����N��<���vq*&eH�B������G)��!I�]Q�er�ڨ&J^�M���3�7�ewL�ٚ��t�1��w&1��-�$��{
�5ބ�ym��f��	���S.s� �yY>�xOu-��=+쇳��]�Ęï�tE=X��/i�#���U]�gJ���g��{�~�k]X{�Q��sYa�iJ��^�&�B:蚦g��k��!�F[X���K��q�<�aܪ�A�^f�g�5���G�������i�6��"U%`��'��u��蹵�+I�I�s
�����@�y�F5��-�T�t������k�rO@?���qyM�U���e���F��P8�S,�h�52��MzAc�5]����(˻@����BӅ�dh���D��6���y#r����)������(�*�>�vs�!bV��w����Bu�p����`Z��"�kf�9dx�D�Q$y$u*7��f΋����E�k+(�x�8�t�h�*��V��h�?Y���c�;����$yeV��B��j�i���Y�^�;�h�j�o�n�V�liޮ1q})��
ʇ�zm&�]����Ō{�y��+q��N�-�=Fz�)/�q����k���ȍ��>�q-#UK$}����|�fNkk?�֜匼=�O<�vU��۾RbwP�Wl<�HE�PG��ߏ�S~Q�#cףtLf�1���F-�\�7��K
�sU*�F�{j=Ł�ؔ��.1������G��$?&����'�b�o'�Z���z��6�����[Ѩ��~�n�@4�ܱf&��Ѧ`��?�0��wNEoyq�әU���v�[<\O!��q�7�U�(���p��_�#9t\�#�VR��r0��⨻����З�)������s���S��������uQo�������Ep�6�wm�2�v1�R� Tf<�q�k����9l񳫆�RJx6E8��s�ra���b�\H9L�y�cQT�u~��N�݉������*�9p�
l�I!�K�-S��q�hق��et�4l�Ҏ�����>��4�Mcщ�~�����R�G�ti��ݼ����u�V���_ż���A3�oe���Y%�5�5���i;�\�j�7E�G�";�����Rߝ�����v���\��֓?np��;��dv��k��B/߂�&_Yu��y.Gql;���߶�Qʳ�/�g�OEhS\���F�N��\M�1�e~;���2�g�k��#JJ_G-Cjʱ�4�/��~.�;J"�g1�hz��$c��J}L�:�o�a�b��NTYy�qL5*_#��� �c���Q9Yq'y�ǢhV�,�ϰ��S�� ��g�oy�(#3��w�9���v���E�s����=ǉ_h��N4E��D������yF>�����.��$Ei�Ntv��E �K���{4~� 0�T2�k��x�C��[�ĩM�0N�ߡn�3���3�;��e ���� >å�#�_}��dr�ᮖ��He�FEDR�)]�����޺�)��-�	B�+[��hֲ�̿ �Z��T,�����e�b�.�0�-)ꥃ�fk�ʜ6t8�9���*33��������`�H/YmW�Q�y_���n!�KϚ�~SJێPR}!k�O��MU��s�+r4��待��5���:��i���͡���t��^��W���\|y�u<�'4-��Xu��gF�ݲ�?����?XZ�C�`	�kC@.�w�4��s�%%��������8J���߬�žMp��hԶ/���ۆPh�;��V�I	pb��Y"l��k����|ƨ�<�pe���5��cDX~^�����!'��3����l��:@"���rؑ�|
�D˟jg��5��oXI�ڏ�38=}�W���%6�%�n��d޴7΅���ϞL�j��������,�mV��,N�lj�a�g�g�b@���3�M��Lj�K��Tm�>�\PO�0Y<I��[g�b5�pC��l����W��γ�Y�EQ�����o���/���9�2������������	
�Ʀ�
d����M�������:����5����$��� �/�>R�T�ʬ΃s������`K՞����a�0����}_�N�i��#��q��J��j&���`!����?`nF��l��
��N�4n)A*�@�,#X$7r����y-��;ڼm��Ͽ�Qn�|�4C�D��q��>C�R������Y1%���{=��NQ��=�&�G��Hs/e�oCD�"���t��dY�@�����o���q�L��!ô�&)�d��$��Z��O>J;���j�%?�V�2���WK�G}��39U�$b���7��J�K;��3�*J���0���d���0����ѧ���ҔUɣ�|3��Qӧk�=�J1�a����b��kM�>Nۣt�35@�*��a%4���R�?�j��o�b��қL#ۓ��"��\��Xr����
���=n>O��?Ua�[~z��������A���?&�����"v�5.Q���iGgaL��9B�֣��������������ڙ� 9��ICߢǜ�A��u�;�{9�[A�����%��_S��l�Q`�~��<��~@ŐP^������ރ�|�>�-���0]j�V":J�>�1�D=�����zcWi��J*ɢ�?ev8��x�Ȟ� �܋��~7��CţTv]w��ǼBufrR�3݊$�:�{ު���%\V�Hx��>�O��`�W� �Fy��3�t�+v�r���^1�V�X�=�������K3��ip����9BNhJWo��<�
��̇)����;�\��~�I��ʇ����)�,�S�F<oob���T?{~�B.#�r���U�d�͎	G��y.궸F��IR��C���e}�nt�T�y�b^�̪�I���x�H!�u����+�U�t��h>I��5Z������U3}kQ�"�r�*@VL������4x�-��v�ٳkK�*Z��F'5��g�~ɟ�UZ}�B�%��lKx��^ϒ'T�k����%nDK-��:��X�4NK�#5{%2���J����D��-3/�{N
�g茒�s(��Z^qMv�;����Wq�7f���r�V�27��ˤ�_�뙮����<��Ԫ���<BR�H>�w��VP�����L���{�.���e���f�'������a;-��+�}���|s�
�AVwg,�4�
���b���bn�*�m�)�~AՅ�2)�\��1�61�޺���z0CE)'����X<��>���`/��i=.ģ��tSn����8w�t���Dx�'���%��*�շ�n�i����2��8�Ü���V��D�
��n]1��V"6��i�om�!/�[��.�JI�)yn��v�2��iQX�?��mV��L��G��J���p3iS�c����xw2H姄D6��Y��]#��KVB�Ҡ^LSxrày�uD��.�L�������ݫ�ے��MLx�!�k%��%Էy�)�ft��bFxChVƪHG�K��dr����8�Q�a�K�J+��2 ��_sq���;d��gޙ���r<W����eO���pEI��>�b�آp�ĉ�mW���(K^���Yݴbҵ+1~pL�c^�{ʫZ>c�'��?n������v�=��4�DHJ�֐�a��Ji+��nZK�_�g��������BAm��_����~7�F���)m�>M��+0GNӨ$�����VN�.4/������oWV������kCj=#����E�.�!T-N�{�Z��E�Z':��������.���ǅ���%gh�%H����,*��D��8�}�����K���� ��S|�o@�B�ʔ�c���i&0e
й;�1~��;.�&�*��^��}s$�;	�P3wr)+�0]�g��IZ4�s�Tkxz���ϭN��������c�[����p�8w߷�
Y���]h���4����I�J���hգNك��i�I�������G"�6��2�ߵ��=��7��e�����W�B��0�9��7;�x!J���QH3a�K�	�NR���G�P������o/��D��$�)��=�L/,Z1ʕ��(Kۈ��(C�7����HD�=«P��85���9���VU)�j̮��&1� ��j����FCo[~
n0>s��������v�dq�ܻu�Q�N�AP��7��
������ybب!��[�8�&*h�d7�5�ػ5�!�gL��z)�ϸfx�#�]��5lԪ>���W�[y��M^�-/�������\\��y������-V�v����>D����,'^Y�omܦ��UzVa�~$R�Plf�DA�$p��#��k@��}3!|���#�>n@���S�Z$'ٷV��(z���TJ��@����]�	r�w�gM�*#�`2���~���B)�Ce��5V��nZҢouY/��t
�gn��>���Q����������G�Pأ)���vz:\�M-�Vs�u�;����N�j��a�ۈڅ����A�V_�M����V�cة�hZ �o9��݂�H��RXg��$(�41���rz�Q��C� ��~��G�KK7�2_��9��sLN��7)�y�H��c��7��wC������yao�خ���$k��y(Ę�Zߏ�M��g ³�#7�=c���o	��5#�͎��a���5�6L7�hk�k��WX~�����Y�3qgm2>�0�ؙ���!y����u�83֌68��o��{���6,D�L��r$��|�< U�|���
Q�!�>�7�G:����į�>;��,y֤ăX��r���j��4��ΰ�����TV0�~#��^�+���k=]�hoԋG���f@&���J���eԔ�h�=����~5��O.��ᐼe��1^��y#m�H�{���N��Ѐ	�P�����	�U���B����\�3L��Z)>,���眏W��%�Q^+��X��������k�V���̄����$NX�q-��_�g�S�&-=*1è����%Q�ä��z{x�x1r��Q�w�l�����芡ꮌZ�y04ؗ���;��^9{�k������[����&�H`[T"9]n���\�K�o�,Q;�t��M�iY��¨�n/&��������"E�z�����;c몿 ��.H.N0��C;lM6;���Eo"�e�����|ޓ�l����o9��
�����, ;R�H�vl�[����2��;�9��g�Տ�������3�X��CCN��Q��)����5W�f�>��ǩ�	�Fi�$YG_��C��s��BQ�,�v>�w��)g�_s*U ���aΝ��:�/�S/��^^�NY�;4���g�,;���
�m.NR�K[O#�� ���>KO�Y�];�Ӟ0�l&ȹ�g
���Y:P��<��^E<�H9i5���4����������~�E���[wQ2��7љg���n�υ��͸L`M��7�-��?���&8+���o/�0�d3r��3��̓K�_���'�y�ˠ���x��v���rl��s��O����ވb%�!�B���w�CPB˲��/U�q���܈.�dTS��RWbՠ��._�u��9w�͵d=�J�i>��p=��4��4�<Oȹ5�G���$`�<�$zjl�gQ�����q{9���ʉ��M�3���!VG�t%�Jԋ�K�%�7"�o�ká�'��֯�*Q�~`��[���[�p�H
bU�_?���\+Iu�Y!����4}굶�<� r����z�8吤爋U ��3���ڍ9O�#�6�>F���A� �=1�`�^�cxV�0�ү�մ�QD��ȑ��P� ɢ��.��o��vL��0ߓC7�J?5�BC:��x��>$��c�|��>��Cβ���?c�U5!p�N���B��ܜ�[$�W�W��?��ۢy��I��;r��̆8��k�7�uD������}1Z���"��9�1�O��sMa�� ��zz�&\4=%�A�H��1O����������^�z��߄[�k�2ȿT�C$G�N����֋�J1W%�qՇ���*�FvP�Q#'�r��
~Y~,R�#��;�C֍Σ�sR���H%����=��`)h�Qf�,N?�Z��_'{�/2�냝��̂o��f�O����q��Ak��"}���/6���X���R�}�"�of�Gz�����S6�I@#�\��K˽~�I헕6b�=�/G��JpTX��וk_WnI<�,�+�o��$�sYQK=����,�F%���u�x\��s���� ;kB����ny�em���^\ y�!�Z���U+c��z=��P����~��Kh$����֒Әf��%L��?Ը8�i�6�o���w#�	c|8�Xw)�'��7yE���H���&��w�%)��,�N���2��!\w��P�]Kv�����%���͍%NK��l#vQV�Q-�N��0����p�\�T~���z뇦��{X�iF���[�n�Na�]#JH��tw��1P����F7_�����/�p�s�s���3�"�� N�{.���nP��G D|��I��4MX��k��~�F�vo�<ϧ$y_���Ud�ԦX��V�М���4���5�>eE��Q�u=�H�f�Ņy��k@��f���I��T)Ѱ��{��X���ё�M|u�Y���M��	ay�è�/�˙#���=[���X�.�h�K���j�U"V_��.?��;jE|�X�,�0c�!�Ph̑��t�Z����#�B����<��Ӓ��>x!@�ae ��ý��%6�È����t�\��4'�7c��d�}���_����q�+A�jUU-�Vs��8G��T&���7�(j������h�|������χɹ��Zvx��ɺ�O�t��Z���� \tZ؂7�D��ᲁ/�-�����p��I겳�lJ�u{(�n}?�z��K��=��'�DbUٌ�XE
��&���p;I���P	�;$���>�R���޻��V��Ǹ��Ʀ.9
i+֌�����l&
��C���-a�u�xD�Ԣp��J9�u8�J�p���˴��W���ᷧ-Nˑ��ǣ[V=e������&`� �IkT9�yBC��*s'*j�ĝ�^�-,��*�P�I]qss�:�gu^��s���G����G���.�(ށʴ�����;�*tm�p�#o��w��P�N�ԋ�bG�)� S.e���MI;���CT�oqor���uj�15&�ɚ�]'��a𴆜&�`����`J���#4���v����������a�j���Id$W���(��"	/��½hg��>���������=zdS2��̨D��O��BBy�_|��FZ�&O�T-�x�E���=�����Df��L�&e6qStf}]��"�2�ʎ[��%�j�v\#�[�/.4�G	���TGG	{���V���FP���ӭ��1>+h�)d�e�۽���S��pt�=�`�k��&����*y��7��E��r�}����ӥX̦⅟����F���˦Di���&){ևlO�hO�QY��v��i�HP��ti}GA���	�HnM�T%� 1�9oE��0U��u%WjjZS���O���c��]M�ȳx�ߌ�����ᴌh�	c���#�v�}��/�?R��.�(I7��RQ�����2�5��*a�t�P�lL���ш�lQ��i~.�Y�c�N�l�j�U*k�ekwD����.�sc���O�:���" �[�g+�XU��沞}[���B+�י��F�p�����g���Q�;�D.��&��~i�1�����~�%����i�z�"�C(�]�[/�[>q�������	�my���)�G�<C+�:QݞYgI���y�}r� �z��3齥J���0�x��=2�u��x�wH5�8��F�><P2���w�����Q���a���!�?6�.i���b�5Ϊ�+��#�nM����`T�4�e-ί�����E^_����II8%C�E/�no�
Wj|�E#y{9{�J;�C����]��/��ݹ�21>@��tV�����8{W�/\�:÷e_��c��
? \yz��)"Q���ۣZ^I�1�7A�TO�=:��\�2��E�^���O����6�Z#',?�=4�L<�C��w?h�m�/���+���?3�f�Z�D����?/y��`;(Ҷ��w�\p��Ti �w9=M˶J��Ѽ
hȴ��U��S��L�)�'ҁ5MQ۸ah�^���Aoې��I���\dY����o�s� �W�5�!3��#�U�E�5���π��cEɜy��1_�'�m�ތ���P�����YU(`%��/�$vn�d�>���{�����[B���m��Up���������]�LϽ��/�Z�����:������B9g
�������aa9�l�U�a�+����v�)�ܲf�{�*�@����Kbާ��Y�S�4���V�EY�[�
��$^�'������36GP����n/q�7+����<J�R3�?Jҭ����v��/�}z�a�k��GV���1��|��n����Rv�^���D���a��7��lRҰ�6��z�z7�a&��q!��,��qd�N��k�2�j�//��d���*��$�������j���9���cY�z�5 �M0�f�cRE�����s�2~���t�Ƃ�X�`- Q���?��w�z�.;?��v~��v0�*6�!Z,/{&c���E,�&�c�*���F
wClT̿�²�x�n(*�,�a���F�(XC��l�nK~}�+P+�筨S�Kb^k����	h�#@�W���Ϗ��Qŵ���Y�r���SN6&�/I�S��J����h��/qT^���_��BH�����̋?�	�;k)����'zߧn��jN�x7��6�����3�]�M�v��V�X��Xݤj�l}nt�"�PN}�u4k��ELj��Cg�	�����j�#���/>(K�v��ɥOX�;<����u�j���N�cƦݪc+Y#��Y>5ya��>.隣;!���#�j̦E��H�/���v��&S
i/�����CG��<�K��L^� l�l䣞�lb&�͍狳^�~ֳ��/�̬�
\�Ȟs.:]O��G�Vn�(��ݤg��P���;��N���pj9�-ь2>�h���[׷���07=n8��@ƭ'�)Q�]D��������XOM�S�X>�q�L�M�:ڞ
��JS%����Ex����^���!���{.,���ф:ٟm��X�ퟍ�Vͺ$��-ϥ ��<s���mD�T���T r:d�_�U�Ԫ�T���+7C9d<>U
bCĞ����(���\�R��h*|z"g_��d����O���,��^O_�g�d�<1�bE�S7xL4q�U�;�׵_n�M�-^�m�lUH.L[�Oư�����O^�'P�'(���Q5��%��ίA���'ޕU���yb�s��3�Y��F~,�֓V�ew�P���n�ef��s#�>�m��m�~��tƫ��L�--6�K>nj߯��Q�܁�p�h�z{��O	B·�,q����#�?��73�+&s�n咓�]���i#F�܁dR6��t�\{��Hb>���viw���a��J�^�i��A���?-����;�/�Q(�0xs.���Z�ME��j�Ir�s ��d�Qv����~d"O�CYce/9�f(�GH���d�S�C���V�>>8^��[��n�'�b�ύl�Nz��)�n��=4�K�h�	l�~k�
�-��&�/j`�B1V��`�hn�IH��Ȯ�TvPw �
y�T�M������'Y���jw������ɷ��O�<�����]�-��r�v�9����rJB4'a�`M�����p����k�Y/�M��S�|�[=<��Fp�8�ɪ���	5�A��f��

ݢ�N�[�S�,�/V��~&�a��H$Q4�P)�7�H��4[wǬƤR�Rߵ�w�ິ�s�����xi};��VN^���K��.�eJ����~�`hl�����>�烵6��ù{����i�~�4&eX��Nl�ǂ����m��'���Z��磢a]T�ĝ�����Lə ���6��!�`h}�r����7�?JުG�Co�<���������/����J��p2�#�t}m��_0"?�-M!�;_hz~gˣ'z�Lj������E6����&�,��F9 =�*��O_��c��l~�K�N�A�J�6�1�-�V���78T�%/�ڍ4+A~��Ga�t��s�O���aFYY�z��憘ם��E:`�k�K��>:�[Ll�
#l������������i�C��{�sk����c����)��TF���0\������C�^�#�loRɛ� �xy3Yg�����ES�uÒ���^���-գ�WG��{�^���τ-`��%������f��L�Q����
���8�yK���2Lm�e��`�朾'Q�1�ֺ)�ɇ��{����95B)5�͕����;����iw�Q��Y����� `�B8��[?���Ft'�w��s��K{����[\ҕ}��D>��!�"�����S�i�}Sx�M����e�3��9�
�Ҿ��<�=�Q�;0�<Vߡ� ܚ���sa�6���m=H����n%ڄ?��a7��BS�(�
� �7MS�b��;Ӻ�i��d6��>7��̪&	9��O)}���8�zE+%},P-��\:�W,�P"Z �:�#�'M���t.�Gf�)�9�Sy� )ׇMK4c�6�����q﷟1�Y?.��lP�|"�m�\P��d��y����m�Szf{P�U���L�4����C~KF��3�(և���zH�u#0�\�{�7�v���3������2UW�)�A	��?��)V�\^������T -����f~�'���Z?5���l�|:�x�9��r��}$8f[�����G G|g��xW�BfJͯa'�޲Pd�m,+�אꖳ���u� �瘬k�W�� ���{�YF���[���!g��6�ȋҀ��]o��ω��|��:�wx������v���d�~.�O#2Yt����;�	����TU�}���r9��&�1�h�z*��M�y�n��(6k�Ղ�L��"er�iM�?8����{�S�lT��r����g?n�(���*�i�䗅%T}���e=���~.eS#[?RB�w�!�L��*G��Ӏ�S7}��d���"���e̽ ��s�)X��u΄�u��r+3�Eji-~ދr�Z ��^Bb�A�}^����B��)2�D����Y�^S**�ܒ�X���4������yT������8�Ph���+j���X;���_���L>��oc�qW������Kr�+�c_J��"5[o�j�db��7b�q��ug�6m��x�n@p

�Rv�a��ס;&�<�:n������~�xN�I	?)$�I�8޸�N�:)�'����E�úz�|m�uI�),G�ܗ�J�i�=��`�,��V��6z-;Iv��ANj�Fh�(���J��@�y(B�?f�h���p	�H��&�
P,�N>�_�ݏ��h�k��u�-=����9�7�Ϝ��5�^�x��Z��Pˇ?v/!��9�C'�s���o�d���"���y*��v&� ���i�^/V}����^��\P�k<��j�"~tC}�7&�v0�RQ2���J��t�Ni�x��K�7��[	�����ד=��8C���:�}���vKҪ� ӯG'x�Gk���# ��o��1�̸��TE.�>�:NYo�3>WN��'@�����G4���d��:��}.�>d����
������� "����1��2
���k*g�li��_C�:�� ��`��5"��c�<�%�A'���k���DI��jҥ�؇D���%�c�v��t.�c��-J�N)�e�i"�*6G\�T)�y���Yj��ѡ�HQ5�{�CϝIm-�l�sQvι��`k�Pk�P�]�b�ޡ}c���������(����)-d�$xj�����u�W��8/��&���/�ҜC��g�:�F�n�~�뎣�Ѷ������H2I����!�6��� ���`C#*0~*gq>��0ʨ�?�hg�m<N�x[��<~�eOOE�k�����?sOfϷ�K�H���E�SJbe^��m����d/�`U!���6�{ gZM���~�0��Ȉ�js����=�����'r\�i$�M����Mst+��b��"�!�WR���5l�ٻ`���3]E���PR�#�����:nD֩�O�MQ�HL]�1E���,Lk:�m{��N{Zm;�7#[7�����S*��>RDǦaeZ�}��vRrl��Sb�'7�Ah �Б�u ��%��4�ca��kD�i����6̖��g������*�`.���v6�i��غ���!5���W�<L��̏�{���s7N�&ӯ���wA5�d�`QTW��.���
����4���M�o-)��3&N~bm�{�&:��x%�'q�Bwq���);ƫh����_(M�a������Y�ȧ�3��_�?�����ԵFI��{�W���#�2]ƹ�����e֎��i���*&�-�ءFʸ�(�a꣄b�͠�_���"��[^ i��}uwƴ�鬻�'����eRo�|�O�o7tq�6�$����Ø"�j�cL�T�Ŏ�T�_��;mؙ�WA�����-!� �����N�����ǛO��5ǜ7ַ�+?����#����W��g��D�^<����uzV1�
��؍E�F>��:�&bRĖ��A���^ܟ����}/�n�@R����[��X���U�IQv�jX�I!��~���Z-��Laۚ9֗|O�෼?�E+�NM�>xpA�3�:������{ϨV��c��;�	n���-��9 V�.���wD�Vn\�.�P[I`~����ڼ\��L�j-LE�P��`z��c=;����W���X�������&���q��v��ֈ�5�jS�(c�`+�)�{�䒺�����c�����[����┝��-�͢wr ���Jȩ�4��	��. �COj�Q��P�dL��UuP��DW!R"^��8\�lŨo�Mϥ9�$����_ITCg2)�����9�ʴ��K�S�Lj�"�Oo�9�0�o�G�8�tw���B�9���y�^!?c-��b�s���"	;��l8YыF��ĢLn �a)��O�:�s!�t��!|�p��mr|�Rx&n��2��R��(	�z�<&H0~m��b$�$u��x��j�����'%�B��'{>n�������R5t^o���I	؁���{�QK��n�ϬVz{�9V*	iL����c��G!����e���t��᧍D�1/�����P3�k��k��ws���O#�4�<^���(�A��.�a�\��g���:�m��"�
9�Yh-]�=��0���pԦ�烨�6[���5���x :6s����k��o]�F��H n�6y����z&���-[`0qe��+y�S�3sO6R���������)R��H�<��-��yk��sGp��٠�֋쵘ssy�O�ή���d��^DƢ'u���ig���-�շ���Nj��уtn|o�e׿~F�j*t}1Wi/��؈a㛴��t��!�a3��>ݗ��@Xu5�*|���m/Fps���!��ٗ����E�Vf"ݯ��dgI1�6����+<Z6��Ao�̵��6oN��r��IFw���e&����t�T����W�KN���^�Ī�lX�RFDY�'�u`�lq��ܐg�*�Ų��������o��0���}M���'��l��ct%<�����a�e�uȘc]Ĺ�m�R�*u^��7�j&_�ꕎ.��5RU7+��`�<�ײ�D8��L2~P|���tw�,w����r�5Qҙ�8�pq��½|d��{[}��z���zAR�5�xTWr�R�ۉ�6��+.�f����{(���,�,6>:V����v��ԝ}k�Af���v�U�t���9'iΒ�>��ue�tN\xJ
e��`���6�ng&��s��w�CJ<Y��rZ���3�\�YZIx��A1ˉ�n�qO��R�m�_k�p��)�&�{p�������Ւ�.�|�����q9��V�ttlVx��Ma�����R;;���R�����l�;4�㎣�	�'�b�t��NSn�=�@��`i�^�7�0No�
mD�%֍ ~�x�L&�g�}�I=��{��(�� ��L�CXPL!���iw �;5W�b'������B?���N������Q�j	𖱵T��I�6��{œk�Np��/ׯ:1i�40�Ϥx�%$�x,�E��g��&��1Yy�'�Ӫ�O�g��7B^7B�Ŧ]���7=�D�:�5��w�f=<E�Pĕ�k��Dٷ��$�5E��\y����[e�65ktW@ŀ��#B�w"Ap�O�����n{~wی܅ŗh��[���D�{�Zwb���Ix_y�cpWJ2�G�"���Y��|#$�'o����;�L�\�!�<��Iൖ����w����Xs�-i���2����庫����Fƴ!���˚+�.O2�ڼ3�o�����E��P�]k$T����*����n�
�G<z�ώ��ٝ!�cWR��즧hfZ���&���6���[�Z�
�*����.��%o���ihK�b�����'?�����v(��ڳ|�uf�Gq�F]�ϝ@7�{m�����vL����<(���H�i��gJ�0f1�3�l62�X)=t�Ƙ�e��g-햡���B!�v�@?'���-�������H�>���w���V�[�[��Ŭ�J6^b.t��M�X�B;��Vuڜ�,��<;��1�c�+˯�b�%j��kC~�Tx��0D޹;�|�:%����d�\�0uP^L�MV�.�8=���l������5�.:[^y㠻J'=�aջ�y����rRŌ��SI�ւP�������fzA"3e_�'k̈5Om��]�j�h/�V��)P\Ȅe�:�/������ᙔ��hG`�1ﭸcۑAu~R|��90Nt��p1w��y�n�5�R]�mZj�z�����P�1��F�\�Gab��/���Z.��Yf��� I��
�{X���n޴(�I��[|A��>v�9��1v��
ˢ�mA����첤�M��)�2�2nχ7\7��]�����P%�fI�-���t>��м����@�CE�"~t�r�0��,Y{��v�d�yN^�6��f��V5mG�z�&�Q�'E�����v�Ā�]ҋ�%�����m_��rj|<�7W:d��>;F�}���9����1-*�[L�O�*"��a�����s�Us����JVz�Y�d���H��&��m��Ơ����k �m X���:������:K�In+�߬�>9���I@�{p�3s>_�_i��"4:RoW�VfV�L��h�4���7�)X%}��W�c�����-��3��i�kG��]E秧?DFL�����g��獐� �U����X�L�.�jp'/�
)s��;� 8|�Ѹ8
�J���2槹%bcnL�
p���U5V6�kra�}�W����/d���i����]�����%a[B���W՟��ߓZN#�4-4�!�Y�~����G�c�f�,x� ?
��F`��[�gqb���K�O�vD)��-��yS��f�^U:��ڽ��4���K+��݁om18��XӒ�"�:��.fЌ\bׄ\⇸�W��n�	h5�3Z֞�������b2�Qg��E����"b@)9Q{���f�C7���ּ��KiI&�3
�����Iu��u͊�%���<�M|t�Ա��� ��H.`|,�����b������e�˻�2��olB�����+b7�<���YĖ�[�	j��z6֜C����U=E5`���|�mmTjN��.���4W�0$������j�ܔ�Y;b\!�z��H*@1�p�*J��l�ʌY�^�m�J���J�u&��������߉$Z�rz�Q�B}�����)��i���Vn���te<�h���+��~���
���t^O�#���7��kH�����~̍�_'��3;�ڄ�?N��ʹ8��CeJ�^Ϲ߬=j��i&׵0��
3�+�+@`�63�����NyHw�k���nmk&-��D"t�ђ�� �@����0!C:�^��~��J�KP���w��1�k}�[.��10��PX#ǉ�=z&����Q�L���'o�T��a0����:�i��\Vʆϸ��0s�Z<�u�S���|6���_���I�pWk�$+`�ͯ1�#1?]~��BA@�F9O	�q s����࿬8?����Ӱ.��T�:$��NL3�w��e������� �Ǚߺ������1��l�ؑz�ws��N3�<Mhw~��{Q��LSI���B���j�d$xd�_�̉{�>�$�5�3-���uK2/zQޠ�z��(��ϏC��B�	�� ��*KhT�Z���mf&��}�����x%		c�C�F� N�O��*��#{Gќ��uTecpfb��_v|��fpK�����.u�Ht���M�ī>�q��a���6	��jA��~�-?���A�,�]Yt73����K-Jz`��{�c�rJԚ!�m;K3wD�<*�z�&ޔ��[g��&�Imc�yٝ��qw�ʟ�����J ��Φ��p�U݌^���U�v�Z[o�g�I
�����k�����X�1�v�/~�K��n���l�t���`��Y
ث �p BN���%�P���ߵ?�U+ ��������ȅ�߶_�X������$��\
Z��~0��A�Z�s�"�0^jߓ��L���])�GV�P�;b�\�c�~�^^P���u����q��Z�D����3&���=v`}.�i��B�&�U\P�3V�~�i�QU�*r����hV}c~#��Zw��k%i��k�.�#�t�[�^2�p6n�S|zr%��;����rA�f�`�+`�Lz. (.�Hfr��~�6Iy����jAVǒ�Li�CN��.ߛr@w�
�Uϴ���9>@�-����׆nVO� +;���LwP�0d{���ܡ;}�]�zb-�$�^ۡƊ�����-�?J=�YB8�BЁltF�Et�G��j�v��^�I��%lĉR�-6��K��󛑸q�z!��!ֈ��t�	X@>E�i8��kGg�Ɵ_G�Z�].`�q�M�1���F��>�~�jކ�6��=ܟ�f'�޶�WN�&��2�� Rޒv&��u�L]NB���e]p�J7�_J�`��]o�.vB5^�W=,�w'�z�Ten�Z�Cȧm=[��o뙟�}q6�n���E�Xԛ����Wcz���5�÷|3�qj��G�R�K��k�^�	�|�.Nk�K'	�Q=v�t�42�X�*~մ��gz?ߞ�q����TH\E�R6�DH�h[�ϧ.o����(�&�|���b��ǡ�t��P#�{�1�5ް�\���K�� z>�+����K�h���] S#v�Q4�I��bv��"��Ɇ�O�ë�_H�::� �q+$�!�Mh�WW�c��mh�TD�J��|PG���u�~N��w��Z����ڜ��S��"�y<�'��y=SSdrUʅs�1�4��5����8;����-u��HSAt�eU��՝��j���Zk�>\\�X�Qؤх�����Av��-@�!糳�Y���+N���S$1�e\W�W�%��"/�^�����+Q��Ҙ.P�Z��#�e�iUv�B���I�V�
�#�(鸃���.r����{�Ws�ɗ"��ݡ3� ���43��t!��֦S�z㮵���/`�9�&>���C�;��@o/�!��n�[�6)Wm*+�,̷488a�[e����O������|�XD��mw�s�VI�ʜ�e�����m��#�U�֒0��1@����`)�vW��s�i{�n'� �s�Z�����oR�W2k���J�,̐9��x��^�N7�͆�o�@���oug���m�����I�}kռt������>�֬��[��A�R���K����0��{ȏ�w��UK9D�&�+Ҏ.�*o��c��u˶�zT������0Plz�"l�C\�|��Zb��U�z�p�qIR���ŵ��i i����@՜���n��8~���닰��N�y1wW�r��P��9��Z#�U#y�L�Y���޻������V)�����G�L>q℗K�_���Q��gHF��,��Џ�ԭ�=ϦE�����`�����������_�
����:|��r�sw+/�\�l�+��9��7�3okp
|+L_�t'�����]�Q�����ɾ5TK*L�
�]U V�:F�^7�CV��a���$V�6��s�g`��q.ě+0
ś��*R�\������z�Qj^���;'��+v)�8򵐼�s(��E��������'���ʕ~Wa�����]#7s�t�me�4D@�����WY�6��2������>��CB�S�/�e����B��ۑ��;&����n��x�ݏg�/]I�	�#;�ӡ�JO@6�Xi\0��:@�N�7�Cyzc�1��n4�8友�J��O	��-Ox[C0��=!��cj����e|s}v-��M�`I)W&R���p���gחr��g���v��y4}o��T�GP���HQX8�FK��^�~��Obk�J>#�aM�y!���Z�A�,!�N�F>�Dg�;�8��e���=]��J�-���ϊ��<#�Ꮎ��r~:�������2n�e"��x}%2ʶ(%�-�?����V�����9�׳�s��\3.�po�u7��s�v�Y���8��fN	�n:�=s����4��l��F�!p|�J/���7f�y���h5Т���p(���{j<ͫ����PNRvt���@
7W~Q����2���$b���J����k 퍕���вd���_Y��V����x�X�Ulڍ(e�w͗?�3�&(�3�%9��?�}�|�E�2S��K�X�nX�C�`� 	~�'}d�N7օxz�~�n���b鄹]�S��*��e���'=�����u�-��.o6�fx՗F( �Fz��(FC�'��Oq3?�����} �Ӡ�6��"�+�/���ç��ѧ.YLLR�^hxD��D}��Ԙ��@9x_?���7�p|�ȋ����fUJ%.X���]N@O�F�.-y�E��Z�2��ʞ�-��N���Z��xh�����(vx-�7�9V�FM�>�!O�|�^�� :;o�S��-��A�O�L�~/Y﴿_�XO��YL;�^G�� ������LuJ T`K�3	P��C���OSL(˫��Mq� �0���>��4�2f����Y�)@�}-��g�+�X�(6q�u���8�*�z�
�"��n�0χM��*`��6�z1���>����ƿ��q���)s��U�2�f1���pO�d$�����<�3�2%���A쌑GX� �_X���4wk��@_�홐?H%�hfu�!�v��p�l6T���[ �z�_��}'�R/���@�[�ݹ�{�����?B�� 5�.����Kے��`��㋣׏!����24�wr#�~J^t5��R��_+}[l��]u�,����c�L�G|�޽$kB�vg�|>�K�2�G�Ӝ�+b9^U��nk:��T���C+��.����Y�O?OZt���2��v[������ ݷ^߸K��['�)ֺ�*&�����)6M�Y=#� /2��Z#}M��GU�.��F�>Y�l��-]�y"�1�y������.3�Ȱ�^@�<�>���P�r��(���V�j60���a�{:Lu�'h�~r~/�$]3���M�m+0��ڂb�M�*]�����e��bQq�8o�� �z��q�޼jy1+�Y��/��S1�N����+,T(�Nki����~��n��uIx~�q�����>�**��f�ވ�d~S7��ï�#���n���%]�۔3mAya��#�33��,��P�%,WId��E)���	���S�a�6k��=�E+~���Іgyٶئ3x�ئ��'���n�1��d��"p����v.0���x���`�����(����FYF`s)^i�P���F�(I{!%`b�W��7`�"e���L#�>�S9DI���e�,��o����p�.�*|�+a�9q��:itSd>Aϥ�Γ�2�Y|��M��<����ݥ�\*ڧ�cl_��?	�����Y.�������^o?6�M�W�"A��>��v�+�W\>#vV���=aY����^�xy&:�:s��F�wDE�Kӡ1���wl���U�9j��GaG���_H����2�p�F�q��ۅ���|N�1;+��o*��#]6��A��B���^3������M1�<��%{���f�^��������ٛG��M����(���6�=;��'�;t��9H�c�o���K�w��\���.K����d��j��jU3����v �"�4AF��;:�;�\�s�1��� ��O4�T4�`��F�V�\�և�ZUz2��o��l�	��0u���ei��I���b�;�Wgk��n�3%ϷW����ߌ9܂%�ދ�d�+���no��r� ���K����^O��=�ɲ&�؜ry�`�o���I��w_)��u6���}z{7�Q�s�1�����������n�ă|���0��D�+d]Z���A��er�Cg�����lֺ�Eb��˙�ms
�.�:���g.z�<պhG�����eG7hxv������I�+݇���O��Aj���$\��'O�3��"|��S�3_�vk��۝7m���Q�r x�o@����k���ޞ�x��s�����,�2��NzF�~�t�~t��j���M,�}���X�ӜX;�|t������~�(�^�`lA�
+�����"^�\��5"���F���E:j��X�s]]�띥���؉暑��7"F���!7~��L�;�m�K�1�)�K�\�T��*Y{��\��G�(>�Th*�#={���`t�j�=s�ڋ�%��4�d)�h���u9�o�Y<�3<F �1u)���1����>�;֕66 �	�V;�H#9�ڸq�v��Z[զC��JL�%�Ua{lI��w�20~��NOO;��̖���.}T�T`�>s�Ve�+��ɳ�.4IǗ��ߘ��mй�M�Ð�"j2"�[�jHȁ���9,υT���iE�7v�X�}EC�V,����B�.=��������#p�0�)��4��k;�vi�C@����|���o��}}o�%HY�0���xLp�n��̰���Έ���ȭ��CmF��q"�R*pp��p��`�r�Ή���*@K�?��[�����fk��r�����1Y�^�.�+�)�A���g��J����܀�+{�!��r[�?O"���mg�cL�Z�d{EW_�`�{�Y�͝�z��,-��wgd�D�!�o��9�I�9kOV���?��C�h�G��}�Az��QDK���]O�h0 }�S�Jc�V~;�!I�]�y  ��_��ʼ����@�����7���(`�Q��ɭ��PDa	c���Q�"��c-Wi����k�s�b�ؘ7�Ŧ�W^U/���qM�	�2$���9/��v%}7�����<��N���)#5��;��,��o���-�����~2#��I��c���"-�MNp{9���k�ZG&�3瘩�Up��؊�F �.�o��U�ŵ8º�,�*�|�ڱ���a-_��t|3_�ð�J%���%�����7_�J%�ta|[3~�h+;O�9YmVl�w��|������H�P!�oF��9J ]ٷ?��vU8?��'����Z��N!I�e*,�e4 B���ʤ��|��g!�6�t��=�RO'E���z�w�:6�B�b����@�Fg��tmR������u7����P��[t"W	q�u%݄PCNd�8O~.���d�I�Qb4û��b7^��&��t<4��24��Id�]I���<�;�&�l~5<�G�Xj��{�f��QLV�(�C�me�_�۩�و�ȯ_p�[X�Y����y�K��A�P�;�����%وhwu�Ne%:�[n�����A|�B��`���{�?���y�T�`[@*�j5�]�w��������`��Q猹�����ob�,jEW�hL��ĠoԨj/��Őj硎���j�4]�T��Ydv�z�E*CLaZan�Z��<;I�*]�%hL���;F��|�"l�����BK{{�Ո�8�hȟt�iQ���\��k�'}����R������̏1�R��5c�#3����C�{�GZNX߫A��y�Yĝ��*�µ��҇\)��{F'S;��Ck�GE\�e)ӵM����!IT�Ӆ1��̺c���3�m�y��
�<xk��P�~��?
�̜aV?�'f���Z
�1��7�Eg��('dr�g�&�p���`���/%�J���C.�	�5���D-L޵�op�?�EC�͕E��[��t��m'�7�T4�u���)����'�d&�Wv�ں�ԮP�zĕ.R`X��V��-~�d�C����3EbWi$C8(:O�5~��O�K-�p͏�J���f��]/{�
ʶ�h`�(����"~V<C�]A�cre��Te��"-���
�G,��̸H�2�m�z��P�<���DLT��W�nZ+�%�(�IP�%�FA�aH� ��V(�T�:�#QS-9����B��s��5����z<����4�@j���lL����-��8N��L҃*jȎ�$ *��3I�ɃW�ޠ>'u_;<�!�K�I�j�.�>E{"����Wp��u�ցR�Kqw� ��;w���R܋C�(�N��� ����\z����1���kMYk?9<�G��i��)i�3�m%_�l�������g༈*Q�[��³�O)��R/B�&���3;��`|?W`�>��>~���ō��L���oܞ�+��N1�D��[i������8�S��x[f�Xc�i���W�͗��`�G>���Rj�QJ����.�^�<`'�����Kj�r�|'&������5m$DA y^�x+2�J�ʚ�(�5�r#�� s��P��R�b�WGܽ�a�����ߪB��Bu�R+��o��
TZm|�eC2���l�T<�r�b�xlU��-�����&�b�����R�b�ҔF���}�~�k0���`���0����l�-�}�>��l{4�*M	D�i������nUx\
߲�\�=I'e��A2}�{�a���@وlˏH���f��e�$*1����A���܃�[��zi��,��3�Hލ$��X�ܯ"�鿯�)�/a�|��rH���,Ɓ�?��K�k��יO:�?r�-���L+�NGݚ���W���,"��1&�	ω�O�q�ZPM�`g�R����3yV�E�la�O�T���I�a��6�ҟ��e�ߦ4�>�	~�/O���l>T~j��D*�C��T�5�4��V�Z��;��|�>IY�;�q���Ç|î��ϜC���WI�i���x����J�}���i|�{�V�T]��'C���s���l��+�<�Wd
��<��=�%Τ6>b�酁)���g�C��Ul�JC!n�$([	x|sh:!��j!}	v��"g�T�΅�i�B̍O�2ظ��]�M铘��EX�'dڂ��!�ʣ���l�g�m�1&����^p�M��#���v5;јfڠ�tR��a�'��u�ģ--5�U��_�]�,m��<SZ��"�vx
��uj5�qWM[�f�c�zt��\ۭR���/�c�3wN�_4 �u��ōo��_S^`/{^�4mUb�y��.��Y���d��ڙv�<���e�e+��f�M���
�2O$j��/�_,�����q�N3�N6�?��/o��+RO�d)Er�y����2���_���3���gv�+;��y�����]y��	ח���6f|��j6�$�o��K�Dt̜,=��Y[�+��K�IG���J�rJ�w�(z�c�b�\���Sۍul�J���R,����ns�ӻr\#���jP�6"��|��}���&���veYY �6�!B��I���ڻ	��f��3[��kR�W������ɖ��D�㘈<2f�1�c~�6֩%�ݺ̜_N�ƻ�s�lE_���Y������:�T���m���.s�ki�m��U��� ��v�*��3�r��>c�D|:��� հ³)Kuѷ,�4h�5�/�L>{
wC�����ޣe���D<�ށCG�S��9������o]���:�ƙ��MPS�%�ca�{z
�x��*����3o����
���[&��!��	K
�MCH��rK���@iu?=������ۿ�-t��L�+��F��Աz�՛�����A�wG�ʳ����k�E��ޔX��R�����Tx"O�s�����O�6T���8���vaOU���0t{��I8N�	�g��6셔�����y��|P�ۢ�j�zQ��f4O��rlh�v��ʃ-�����嫧魊�{Ζ��b�K�����/e��&��v*���;�6S�Y��7jk.ϸ]2�x�I�?7)~�I;#!y	rx@�|*�?~���Tc��
,��F9���/	�c,+T�uW���B��l��U�����k�Z&��TtN �^Ó���E;'ص�z�r68��,4�	�R�x��x&&x�0|;h1���/���w��1��bH�P��o�x����̋#"�db�Y����>�V;��c��>���W�ţk�Ä9}����ƣulC�}����Փy�$��Y����^wVFc�bHt��F��󦂌����f����^�\�$e��G/P�Oid�H�9Z��ڙ�'H `����"e7`���'�
��
/}����e���8�^f���br��e�?�������2y]c��x�PS�7>�Pi(�W%,�PG����R��.�lq����D�	�}5.K�� C��=c��>��ll �t)ܙ�`�k�`���	�U�B����I�y���)v�G���v�ǝ:vV�M��H�ú��!  xU�������
˙����Ej�"&���n=�RR�zLMmѷ9�<�P�PV��
*�8��B#c�\Z^�>o�Uޗ�J<g%x*|��P.&��:��=n�V�v���S��%o��o�7��٧*��С����!n99�a�t�,76-�&�o0�R��l���&d���|�T���������N�Xﱭ�{c��9���A��؃�k��ʙ���X�j�Izoc�^s5$�V0f�׋���:�+��sޢ��X�e�[#w�m(Lv��Z�|�}�/�Da�'9�a���ѭ�ˀˌ�Kd�H@�ޡk
��,)�t�J;�O�#$��%�<�8DJTk��Y�����#�:���Պ`���5Cս9��V�稔])l.�����=x�6��%v�Kְ�8��۟q�7�b6EX�p�|s�� K���ߣd�qOJ��_�Bd��_�����C�u�X�/2V�|�V?n�r��;P�]�Q�TVI3��-���)�o�+����o`� �.�����f3�y!��3�XBқ�W]�]���i�����_���/эB�qY�~����[�dڠҎ�A�9���tK��hls�������������?�ō������!���*��y\�C����q���=,�����66B����M��$��7��:��9MOf��JV^n5�R����æ���MX�A�v�#ں��k6�z�/�f�bZ#���AU���)L�j��s~b�)����v�z��x�Y�h�������&�ٱ�;u�����$�'	;�-�-�n��Ɖ����
Y�Z��׍#�u���}ɇ��Ly��ɱ�@���M���̋��YCk�qca��������qQ��
r��D�x�CY�%�V�_.��[5
�Z��<eB!����O4�g�����Ű�� ���
]�x�Fs~��u~��)��B�-f��Ձ�ƿ
q�?0��7��MW�����'�x�'�کň�.���Z^=�d@�_�>#1ԉq���%+�� o�1���n�S��`&^4��A���G��w�J
�>s�CWn��ԁ���σ��b���(��a�uNf��R�s�[�-��،Mѥ^0%�%�8Ǔ�\��ϻ�<Zˁj�~�c{��Nes�N��ϲ6�n٘���ZV��&����E�Qnb�N�&�ao[�ӂ�+@����*�l��E f;���Fz�	���@>ĲI��Wؔե5��f�3����	����1�ê���ʛL:L�2"��r���
\�K�3י^�^$XU�,���Ef�z�'�Ҩ�A��~&g�5Z���i��QI,�ߩJB�O������1F-�Y���}��w�l5[
����p$�M@{�p�&(-���[_�Z�:##\�SV.َr�?اfӴ5C#,�磴��ԛ0��ͱ?v���D$<��nost��RO% jSA������dy���>ȝv�*+)�(®��.r4|�2I�󧘈z���	����2���Ջ���A�U"l'���"���~ǐ���,�d��SA�:
���\sl�Q�`�D�����)��Lv9|W�p/���>���h6o�����,P^������4O5;���l�{�߰%��bm�sW/W�ה����y������]ZU8S��	�g;��) �=���[���1�df���XI��A�X�y��[������>����2ݛ��S�6	�pB������D>�Z�I,�5�~��L�F�#�xш{�^��"�k���z��.6�a�������!�1Tռ�(��y�b:�-k���E�4e_#r��;��-�r"jM8�Hۑ~?)�@����}=F��g�p�y])�-��ɼ���''8$=��W�cDC�Ѕ�2�۽�m�&&��w��-LPC�a�d���O�&���1W���ʝ2P�VoK�Z.�\��"���!�Co0D(�Q�o��� �)~��H�b-,��U���9؃lK�V��}�/I�b�4j`�jL:��Gnt�E	��Mߊ��mA�K�K�+�2����&����CJ�s��w[����[Q-ȂB�.Qi;?��Z�(���sJ�F��KR�̏{d�}V�����#�y٥#x��n�q�,�hzC���xn=Jc|1a�AR}�Nߴȍ�zv�O�6���>���.�7J�@c'��N��>w&x���[�7�\��GQÒ��|�zĂ�/�c��\N������Xu���7�����T����!� �}�N�'�r�g�W�z�.=��d��D�(}m�Zh�x�k��>e<=0�5��U�uIZ,������:������Ki��S���I�Ȋ`Y��p�~��%�.^?����T��]�,�����[�G�Fw&���j�5Dng��S��J���V�����+�5�i.��!̂Ѡ��V Z�yO����j�Q��pZV��(+1�g�|�+�OϑM�N&�5�/�w�;/�s�c )�t�6��'���O��ח
��ٮ�%O�?�τ$��J"�㦅�BQ��;�`q� �0oEU_��YM�z%�#�s�o�-^�@f���v�6?;���IަGJ�iG���Mo��Tu���r	��ݝ�v��ְNK�O��,�Cm	^n=��D
~�<����w�W���\Dtp�6¨��r�i[�{9�*��z�eaf9�=:�c���t�WR岞��[P��z��
WIzqi��#���C�̥I
����|6Œ1�(��!�ޭ۵������W�C�����Կ�tm�?��j����Nĩ�]�x:9��mO�<>��jS��V����2�T\�nC�TG�`�}+�7ʉ�,�^(��nI����H+�/�	I�����%��0�cȿ�h&�M�`'����wLUS�ő���ڂ����R�5�]�mk����<�OA{��'�f��e"N���v�(���ͮdT+2+@~���
�k�ժH����;�}��C�;3�_����2����Pa���/DI�N��!��f���43���������DaZ����[��F ���
�?8[��/��q�|j�V�^���X(��r�S����K�$��r�`�dVL#�!�0���2�DFKO_��0��/�a�x�X���R�f�m�/�_.��f*�-���oԳ@1φ�I.53;=3����y���-7\|�pr��+�=+���l���|S.lcƠGa� ��@16V�0C�6	g{���c�8���1��~{d�L�[8����T�fl��O�̈́A2]�Kz�{%$,JMz�p�PW䉴<�5님������;ZO��	�p��rx�/21�F�=�9��t�e�yr�h���yO���}��V��>c仞�-,;�7NhEO<+�fUyU����i�͢�ߙ�6^��jΦB�~�z�O5�:�k�m��̴�e��5"��ѐH0n�4�Z������[��σ'`��(1�ɟLR�Q��aW��g��g^�F���B�*>��ŦW�
�a�G�z��$Mٝ8v��Z�^�8��6"l<|���Y-ەb<�`�[��\���u6�ny,��TA�W1�Y,�o�w1��>�w�y���"<YL��T������ �J�#�kC��O�n�>!`lqf2m�z�Pb�r�mf��ݒ�x+��5�`PJ����Z����gh�X)ڌuye��ȣ��c���.
�Q���u2�RHV��k�2;ү�lr�A���ɷ�n%��䋿tt*!Ie�6���ws�e������v��j�O!��9�L���"V��K��1~��H��	o�������?�_��2�V��hƛʘF%���J�W��D�1�Y�Y��$��F���x�DP��,[&x&k���׳����_�cօ���H���.��a

@�S)�h゜�A�~範I	Le��� ��a��S���"8������S�Bo␅�@?�����s�:�w?�.*V<����i�6��s{9T��b��wqU���5o�h���q$�v��Х;mV�S���N��:�E�۾�?�x2�=	���Ebڗ ���W7����B��4��n���t� '��(a<�Fz��Z�%�D�z��o�x��@O��ZU����gļ�tw�E��v�^�>2����	ARcU�G0�n�p-dcPz��M)��g�c����	�wG.j��f���.F�o�Fb.$11l�$-��f�$12�H�:�f0�	K����ޝY?8��P�X��ԌZٶ#�U����;l�mC�z��I�݉[��|��J�d��qK��p��%(J���p�S���/'��#�3)7����֥������v�^o�TqhD�����wJ|l|�6����qUS�Cݦ�3a���>��J��|hm��c���Da��u�/�<�zk��Sf�]�I�պ,����;B�욌�R��E�1�-�� ������h�}��Ej�����H+8dmow��-�$rs����!� �mA$:�`�0+Z؋[�|��� �H[�ئƚD�Kg:�>�
O��-�n��(�Ѓ;d�7��*�����~��r�^�"9Ɵ �w��G�4�� �G��&�:w�:="��c�<@s�5�/�o�ot"��7��c:�r���X�oW�����hf)�?�P������yJ�L�@�q<Y��m��R�����6,�r��1Շ����?�Q��6�4�f[(��u�lhR�����`y�h��(;�=��b,
�.v�u>]�a��t��ٝò�|�hN��s��n��Ds��%�ێ�(�\B{f~��wP�;O]�q�e:��|:��ñaX�<�jfJ�!�ߪʝ�&�#�~q�QA���nT͝�ݻt�7$���(��3��꥖��GM?
��@QR�_�2��g17�͑aR�SB��0�"S�r��_��oP8-�p�u�{K���^�_��䕄M~MCCH�$8f�]c���n�;yɑB��{���.�����b\�Y{c��`h���	���<['��t������V[h�����Fhpu�AҾ�O,��������Xt��K��O���1D
*���6@q��^9{W��xd�`�B��5�fݬ����D�N)�$:�,,j:�����C���w-2|K�J	�(��yA!���WS��NV+l�5 �$H��'�(�c���_L�~��~�JF~�����m"x�vw�������(2qW���F�U��8b�+80^e̼�Z��c�c��J{�$҃o���[82�y6�8��\�f)�ѝ�恎�wK���=������^�형�ƚ���}8z{Qw�阀��A�|��nj��O^�b��[��l����i����#�@uAS��v�lk܍ƌ��RY�iS%�@����7�:�nH�jxO�q"3	�h�-r��h� �H'گ��=�C��o�H���^57cb��p��(��Fٻ`꿃G����_W�(M��~�U����2ic�ǖҖ�}|�+��E�~��[7�?��Ǻ�����a������!�)���w��}�����m�����!G֯�>�v%}�|�H���A���Ͽ�+�S�X�M�/���H,7;�p��.D�G���=��q�W|u_�L �r=1
?�b�-s��8?�;�k"Ra��D�)~�F�F��N26+���=�K�6Y��E�w��+����k�D\9���N���`?|l�k����)�����O����S�:RUO�=�N�]K�0�����@Y��y!�J쵱��������%�ٍ�9WA�*x���R�����R��[6νmϨ�K�� ���m>��w��˧p0��t��4t����tۭ*(�͢����O��� վjs� \���lP8]�!]�c	/4���j��X�6V�7�YYPOC�b6�M���b��h��. $}B^@!�Kv�g�d�X~���`�}q��!���z�NE&紦�ad Ҍ�z�Rd�Щ�������3�%�Y��\�>�4�z��NP��D�-�x���$���ͿZ5*� k$����b^Tբݔ�P^�x+�nt�߄>$��g�k��0.��q^�.�Xi����)��VQ��3ܩmV��"�)�D;���3�O�/z T�ن9�5{Ĩ0�V�M��C7�ZA4x���T���Gh���2feb�or
�p����G��|�Y��j[&8K���_1��	�RG����\*7�+b����e~4yqud�HZ4������a��$���=R��֧���l��*�6٤Q�#���e��Y��~�-��Emn�I��'!摾%*V��w���	�4F�Ҹn��r���	D�o1~��PeB�?.H� �<3����h��?�Gy���K~�����u��'�U�n����'+�[���c^�k[7U����Ǜ�>�BH�Q��b(�~ +����k��y�t�[=�.�Coˣ�t]�"��F}@NF=����T�� d�9f7������4���ףb��'9�Qt�8:RgE���KEUn����lϫ���=JkH L��7��d���>��)�t�y�<~����e��R���曾ֆ�3��&�,�_]W����	m��%=/}!�aZ_�s�~�xs�
I���gj!�5�+���<��Y�<i1���=�Q9K��"gD�6�mS�%Rh��q�ӧV�@�-�^�w�"Z����G?��<�j� Y_71^�1� lM��]R��I�+��/V�#Q�١�YB�����_�ں����<k���ũ�11=��� �*pO�t�ů��N�?�+Kl��j�>��x��#�qm8�_YQ3�ӻ?�m�,%v�0JN�����B����(����^㆒�>ip6��+o%u����֣��3�]���|j�������&�1]�F0�UϞ�|��I�[刦^�]鑢�fEt�W���e���Rq�^�T�w ���P6�z`�e��N=&��/��5�z�?Y	��j�_~ ��2�W�r�⏱��鵔���G"��a�|���B(��G�})�Vъ�!k�B�M��/�'%i�[tޱ��ݵ��T��;u�/|�y���\��Y��{��0d�%���fL������Vd���m�;H�E������$�q��W�'%�ua����ĥ͎W�Ǚ��~\��o��U�Ͻ�2Г[᪞���~��s�S{�2G#��WGǷ�;��|UY���&D�S�g"���&:/Z`!�(ף�Cn<��{S�J�b�w~�����!�4��:ʱ��!Z�[�ِ�m>����ͫ�A����QL��X�����R��m�^g�s��;��3c�v�C��{O��$�X�H�Ť�f^y-�ϦV�;�E���Z5�2����"��Ī��f뚢|�r���W ��L����6υC�l�"�?��6CN��Hl��[��e�����ٿ�<��xMeR�C�����Fѿ�n�C�:p�����Q�+
��eT,�?�f�&�������O/>.۫��Sc�����a6=s+Z�o;׶�p�b��Ѽ��Mv��`~S�=@*��-�bͷ"� �~m=[sW�g�n|4O�B�����h�1fmQ�P�U�á�L� ���F�]�l��yt����I��yQ�qk!�j�7�Gf�S�]���B��V� 9�b`��x��QH�[�^9�1��gw���%6H�z"���Sf�w�q����o˙>��H���Z�i���<�0��w��<	9���+���,L=����N=>3���2�!���+Mչ1�3� �F����L�~��^:g7YWS[�S�{S��_��oߎ]��^B$v ={����Y�gz®���ql"?vz�	U��"��.��K�2D�E'�'~+.�Z9���gט�wI��D{�v�L�QM� G�viŅoh�����k�S��֝]�8	OAWܖ_7��Ki����6i��5��Cb��-Ò����s��Y"}�pT�6O_ U�.`E�K*/y��^8���/0��y�L؍�)E����~gI����T�ޝ|=�mM?��X �<�]�����+>����Σ�8�mDMs��$�n^�����"t����o�6�v0��9�o���r_�17�����گ�QwG9��-
�:M����a���chGM�m�Φa ����⺃r,3���^zH��?ߠF�]��ax�j�s�2^C`d��u݆~A#}�{��V�Di��}@ �D����s��uފV��@����,~���r�l��*)��������T!ƅK�7:�o��nq��i�����,�P����}�!��\\X����R"��Wg�R#!1}X��������@6|A��d�ݬ�����{�b�M;Ь�h�n�tϤm�=��ӛ���Q/�5۾P�0��_T��P����5�.��J����b���xt>MM���6�-	��i����?����qT�(���3�渊.7�:�5���eo|��f\vMq�i�:�3��vz���Q��Tz5ch�/�0�t��7$��Q��������g�+r>"Y��8��Te.%;�7�
��߉���ڮ����؊��׼��쯺`R2�U_�3��O]�:?����*����/��HS�h�'6luf�P�	�@�Md�I�t��\��WZ/Z1#<0�]�_�6�P�j�J�Br�����كP#����is�#�I%��sD��1\���U����� ��SS={�_C�3�J�7���	0>�L�e)�U�j�b9�?���]��"4�顃Kv#'�4а�wl	�aO�J�L,�<�E�u�n���޽-�����Yq�&"(a��t�8��n]�'h�����0	��٣*�Me�j��]�(kEP�/o�F�6�t�(��<Y:���EWv�ޤ����t��$;pӦW���x\�'\	r�&���nN���w%�{wG�S��v\)f����x?;p�e瀲;�.%�f����t:�@x�q�r�:�a=6���2x��v�%*���ʎ!e�]�tM׼yn��.y��)�M\"7�rC4�-
�v��筥�C�V@�ge����X�m~�D��;�m��bG���`6��A����Ҫ�zO��̛��P��.^h��<�Y�_c�Ux�d��3�?��j����b�Mf�h�)��W�v���>4f�S�z�6M���֢��i�̔�7�vj�#_��կ�_
}�4 ������\�~���#����5��ýz��p�!��u��Vo|����[�h��Kb���^�̡.l(�`f���t���O�x9]K�^}��h�B8{���95��nߛ�߇���\��Ů_����A�'s}Ju����X{�qtF�����jUh�r�;6�o�	E�ڤD��#[/7�\��r6��ϻ��<�9�(��i��-'�!�x��L��S�h�!.���6u���N��3*-�X�O�]Hz�������KX��Rb	g���i������z��#�Wm�k�;��-��0 �L�������z"�|�}�ɀx4��Fu�5'��ʋ���MҤ�Y��љ������6f���|YF��A�[7�щ�#ӑ���^�����9o^�6E��zA"�D�U3�;�f���ؚ�T#�c.Uמ%K����VʀAH�J��^D�X�!�����mK��d��G��ݜ��`�$���\T�ǅ�N�o?��j57]z\{������j�8�$�� ײV9��Ѫj���@z�ht�����ݬ�Ӄ���һ�n�-{)�w����������5��Vܧ���0�&�f��Ԥ:�I�Z�Ë�3b��8x<E9+E!Q�[=���1فl�+�20Ə��7�Z����[�tϛ/n�8���X���Пl�S���6��Ӳ M	�H/:���z|��PB�aMb&���
��v�δMK_�h�nkJZ����6��� )���]hד�Ǝv y�K�*Bq�l��mRT�!s$i)�M����e��Y}~[�H*ߠÏ��d ��ޏr�7y�6
rO�"�F����2���,�����C�n�v�� X�U�ڞ%V����A(�*�=z��"����(%�rx�_)�������lNU2�f����WBd�'�r5�x����@�b�6��4q����o�4�R���������>]o����+$H�r��?oH���ϡvPK�5o/�S�=��u�[�Mf[�R�/p��)�v�@"�|7�**�#�B��8ţ�wh���ՙ��]�G�����(��]t)�I���ln��+�;mS ]6a����5��]Ҧ��ͣT,E�et~ɇ{�/�drW�6�����|hymR��G�\�B?�x4�B�>�2�'L���&~�KҴ��tV��<�J6i��b:��'O�����m8ylA%��<;����J$�����&1��PD�P|��}�&F��F0�E�\w������b�Ae�:��o!Ӥ��-��h�$F����a��I�����K�^p��� �b�\�r�O��6z���g�&�K6���<����q�m�ǽ4�Y�ލ��M�]�.��\gQ��yֆ�%5�^k�"u��)aS-鵳K��*�ϟ	���r�{�e�>BL��k����E9���6�^o����Ҟ���yb���Qe��A]���*'���i�0=�@���R��	{���G݃�����j8*�^��������{&��%�6_�\��n+�Y���9�򺯒g������eo�>�*����f(��`i�<k�AΜ����Q~o[�0��=���ۧ�<u�n��m��~��#Y�PWL�nD��7�}p%����j���ȇ������s�_�"i�fr<��[��Zty<^��~Pd6�ߴ�h��2{�ȏ����Q
!����GO���E�h:m��S��V\�d�n�i9Ϙ�������맘�~�z ��Օ��A&@�`J�	UϘ{�B;U7�ڬ����K"ot�m�rtm�&m �g)�3si�[ep{��%��:���6�ݠ��'Ꭰ\8d����;�������6��df�V�섩�c59Y(��,�8�Z�н#��ӧ�2�1� ��l���gl2�����A�s2����嚤kX�Y����0�:=?Kc5��2��T<��{!f���{�'��ޕ�����}BtR�{\a�w^����&��W����%B���^u�͓���8��i�;
�U�	���8�p0�`�d�Ɇ�}c��$v��"��I�p�:�]��<RE��j�u%�f�%h���Q�]t�l{;8��q�݉^D�R	��Gw�mB��]�L����jpЛm�O8���K�"���+cp�e-~���ag��W�=��_��	HިȒג2#w8'<����}&�m�連<`�ED:����&sg�">����^���.{�㚚�i��5"V$=B��"����N{����6�W������l����0�H�	��>(��W��b�Ju~6P4N�(,t���w5���w��+!p�cB�L��W��H����nw���=:8���t8˱a��@�l?>ἔ[��zڹɀ�n�L�G�����p�<BNƃ�"ۼ���8~����i���~D,66R��è
�B*��9K$�V}ّ�,�&鯗 :�kK~Q.3f�ӆ%��yK<���e����D�����Ň�\�?�b@;Z����.�[Fw�,�]�^bP6���Cj�,uI�$��o�;1Wv��4�3�S���|�k�5z�A�>U�Uiē7&�a<�����#v?/�q�G����7��xwO�n�[�M��ٴ��>�=o����2�ل�E2��u��W�U;��U�.G%��� ����i0��	IWVK2��Q�Ń�/��N�op��EPVŕ�̻�1�D��x	�lyg�$"yC�&u�K����������p_=�l|�@kA��!���p�D�t)]�)�Kv���̆Y��R���a��NZ2�Ê;��G���G{��k1���<ˉޓ";�� \J�߬�=�7�Nx�����2H���<)���=^����ϖ������O�S\�fU�:��L	G�e���#���{���\a��8W&�g���L������U�e|]7|�8 �$����[ڲ���D(&Rw��t��FN��f����v�ʗ�}����M�6��.�?�.��1���'��^�O�$N�"\�v����(�dpCO�ԯ���6�{�L�X$��W=@
G6��oRw/W�~���`�y;2�>h�h&+��0�l���RWJ;�R��X��`�04p}O�? 0l��S��Dߔ]K��n�k�b�\,ŝ�m�N����w���6�"�0#�$ٖY��1D�
Ǚ�V�0�?2R��04�����S�O�>��.�n�FsT B��33���.W�t{�[N^]�d�RF�|��\�:n_�]i�L7�Z�ٶ�Sl�*�w��hvPʇ�<��|7��s�\�?d�0������{��@�{aYsp�ba��.b�tr�C�+��"��~C3ÞnK3L�eo�b��pd�1��l�2;���T�����CI��/E�_�	tsF��8+�j�e%�}��ƃ�>��M_Q�y%�Ǿ�l2U���Rw��*rpjӻ��4�b�B$LS� &\�՟����N���}����f�jr�%��-Y-�{�c�Ę֮+��L�XCTi~ګ��+��_��9va��W\��G�A1�l�
N*�2_N&�:��#���w�����/�_���]��*W�E�h5�K�`��:���j�m�����dc�s̗�0+c�[�����]��ʥ��B@��|��m5��bp��A�F�K������~[�� ��N�K�d*�Ae:��ڠ�Z��l*��}�v����R5Zs�\a��]�v�K2����|�³!1���L�!���F]-7e��0��1-;�./���I��׉�T ?��]틕�7,>�d��4������9����Hv/m�h�%.x8oct |Z�%/�H(�-Oށ��D�:֝����.ZW��
.Mo��=�n�M�,d$��nwb_X"|
��:��=�����X`BhQy8	m��.�D*l��ˠ6Uc��I����uQ�m��+��M�|]x��!�cj�/E������AHR��6��������ແA�(s�NŐ T�s��U�]����^�i��4����m'��w��OV���A#���K�f�'T`���m�!��1��5-�<CY狤���)���W毿%����R7h�ViH�Hd�������L)Ju�D{���R MI`g5]��\A7�?����o�s���v��<�~_�[<��qи���_Nr+��;w ��߶u	%����ѴTZ�_�p�n`�Y�-�N�ն�{���dz��н,�d͐V��D�O�4��R�eU_� �����1�b���U�Eۤ	�!9�% }�������a��o��]��i�i^Z������Ǆ�yK�����P	�g�Y"C�{9d��^�GG8E!E��]�|,��Θ�$���ܒ@(A�N��y��X����QX8l2�?Qӿ���%bܳ�_9xqK��$������q�~��,���VʃU:���vnޱ�2�����Ӎ�y�q�g�*$ӽG���.�${F"nsO�"�D�_��$.A�/\w8p��!�\��A��
�1T J��m��	i�zτ��_�jG�}ݗ�|���-��Y������w-�;�.�g
y��S����a��HE�4~���_x�Y:e,_�"�د�c����Yf�ļ�m��inY�|T�m�����"�S\�;.��uŮ���zy�g��$���n��%���ʱ�}�z�-9����� ���Vk�kܔ��Gr=�?�)��-�pP�e$�����R�O�%j��(|��ޣY�@E�F�Ry;�Z]5�5p1�y�-����j�4n�v�?o��[�Xf�t;>������]��=u(���!�] ��ޮf�"��?��ծH�2kI-6[(�t�urNӺ)D�����v9�b0vLU��X��N9�T�;�@/��5Ț��G�����f7���29˿BD�ՀГ��6����I��n�U8l�x�6��Ye�ƬَE��w�G���\�>�%I�ߕ|�����e���5
;�<�����^j�ﳒr�៙�pڼ��.?ZB\H��5�,�I���)�u�J��l��6���ɽfR���r�Zb�� ��2V�)�΢�ͤj�Z濦�V�|�Ii�����y�2H�am~9ГT��j����:*�FJ�n6�9���P��[���O����
����� �#]�H)H	�-͐*��1�9 54#���9t� ~x�����9`����}��*SO���gYcU�w�$ݗí����gՆF�$K�)�eO��=�ϳ�+4TNPF��e�;�h�v�<'��(̳��|���e/�H�yJ�=?�牄Ξ͊s����fp[��(�\}�gWXK�y.�+UC����u���P��q�=b�ߣϴfH-�>#kni/o��"�!��$��g�+C�])��E�*��չ�T�R�K�������|�������h���[���r���b^��;��H�3+�e�a5K	���M�]�����K�'l�Nl�E�L�6>����.���֐����ШǾ@�C��'g�;F��u�^�i��+��
T 
m�WQ��SR��v��lB�2�=ШoP{�]5�]s�V��V�FW&mz;�<�Jް�կk�wG�p�ˑ�������α1�^���� cĩ_g'���l|�!��/�k���I�{K��Zv0�[��|Ǿ�;�FYV�|�E�� �⮒��N/s�2�]��6r�173e�b�̭&%6��:�
~r��b{T����ݢP����y��52Oڭ"�ʆSz�t�R�V u�w�yS\���*����nT�C�B��Dς��ԃ�L�k�Ȋ*���0/�䱧��]��>��_-�������?�u��"䐤%h�r��L雷r��;s�$E�ݍI�)P���,u���������o��M�)	��*NÆ[�)�/ַv�r����]�[�/�$x߇�N����<���h�hS�Ǘ"���41�|R�7������&P�/�a�g�z����7��_VF:����j�ƥ�i/�W`�+�r9���?�����_l<� �dR���Y��ȕ�`�v=U��=��/��:�S����9��Qbrja�ݠ����<ǢX�e���Z{o�Jo%�G�I�ͯ�Ԥ�ά�x�j��b&ƻ���|�a�y�Q�5 �_N�S��>w��L?9� �K�;�$���h����pI���?C����:�QA��N�ǿ����]�y�7�M���O-ɜ�w�&d�
��%5�x	�+��.b_�ZC�.�u����ʕ��
���gG{ڗGY�=����g-t���'���������+Eͺ/7)��/�MHt���c;*�!��t�ˮ�zmO?�f�����13?q%��Q�X��`��,�rY\��)h�}2���F�}:Y�Rݥ�gg��g�ۨ#`Peτ(brD.S,����w���1��܏��ؤ��ہdM�NGk��l�P9�Խ���-�ja���Y7s��6��e��V�G�v�����x�Uc�nDc���;���+j�E�U+Ͻ^�ˍ��7����'���L�qX�.��|r��1@�e��o(~���	�ߓQq@�ʈ.�L�5�p�~��,�3o��´�.���T��ଭ�X(C�Ң��[�¯�.�ݴ�;j3U&	�q
H�|���ڧH������veЭ���"��
�_7��̲&_^
 eK��F�OW}H0�[����2ۦ�%���!}�A\u3Z���Lb���B��-�z7���Iu�WJR�	���ax�
q��z�8q�~7TO�)��3s�84�X�ҫ�8�\y-^c��˯*n���l5Hn�&Ȗ\;Q���G%kl-�tG�&,���1�1����ͼĘE �`�ڼ &�4��M��)����Pk&�E�󜃦��=p����rϼNh�����9���!#���dE����$����V����X��;��_�]Јx(�\_O~I֋�qZ�]�L��*���X�R�~l\�(R�H�B!�d�)Q/�����cJŮ��k��q�z*�fN�IM�*�Ӣ����8\�l�lbz���X�����0��?J��u�&����E��=�L6
�|Q��'$9A�:P<�,1���/���7!��OZ&�-�΂�`�Z����<��ɚC�|�`�=/v��M޵�JHc�Y%9�Y� ������3Y�1��!)�#�h9���
�{�*,H:g�A���u	���ZY�g`��Ok�\��c�>�N��g5�Ѳ �0�.��s[��rW���"]��W�3����e���X񙮺"��CrIL{8�>q���[�P����k�߿l���K��+D����]T]	�eSm��g��J�u���`�1��I8��,y���T&Up���I�	�hm�G�^��Wfĝ`�JIe%��ð��X�}RBC5�x�D���=ӻ��}��<P�Y^����p-�W�f���3�����jJnv  ��f��h{���y���מ����<n����,(;���G���ۥ�O��ݩqIw)�=�NY%��c;�؋L{���Ky���f�� �5El=�9dR�B�&�A5rŀ�3غ^�۽~@a�ݻ��`�"s������xԌ;*��~�4@�)�G4�`�{�nC��M����'�2��0 XX��i����/4��c*�ڳi:A�,��f�ޖ����:��=\���D�ގ�w�kN^�x=��qq�1(���W��ѓ�V�4���y�s0�e�W�a�S���Xx+�y0uK�uu��w%�v�wӉ�Q߈�l�2׃;�?��+�8St��-����|��GTf�_�.�B}}y8E�طEm�U=�D8��2k��|/%6�{N�FM,ڱ�<a?&�24w�ٴ�������&��|4���8<��掕���
8|����K�8�;�.������!_wMm�&��c]0(3�(��y{�Ҵ�PPJ�.���Ş�F&�ր��<\X�R���Lbd��L�C*��/��\?������k$���Y�VHϿ�4Y�o$u�F��a��Dr�z]�2���*$�6+�UU[���_�B��U��9Lo��D'���_n9���[1Ðg1�� ���W�{e.m�+�����W�J���4c����O*0� 4�y�=���!�Xz����9��'Q��#�Z]W�ʏ�|�% (�Z=O�&f5k�����vO�_v�tZi(x뤫�_i�����9E=W��r8$���\ďg�ب�u�h���8��\�bS;��������&z_�����������l����ԯ�L�v�L?
�FUu]v�P���͒S�Q���(ǿQ!K�<�����g:|�ܓ(��F������ &��}꾘�	YD������X1�����p?�R��y�9��&�����'P����A����lۯܡZĚ$6%H�ƾ�<�nrn�Wӯ��la/�u��ݜQӄ����6��3ҎG֜�n��mԟ������ݣv+e�BvV��!��6�ė&)о��D'�S��AŌ��(�V�b�U�1P�(~p(IG:]�Qc��v����Y9���b���?�
e�﹯�
��	X#IQH����nVpx3��L�ԉ㺊��w���$�Z|* ���򭥒+4��d���I�ؙ�ȥ��M�Ji M�r����.��Gk=�q�ȕ�MN@�5��Tu~�I�+�e�SK�"���)6�*�P��Y���3�;J_�/$ A���j�H
s��Re���eV��F��F8A�q���yغ��ȵ,�#ŉ&Z���V�������h3�4��R'�v�Ϥ1zVޅ�0A����~�<$Ic�y�[���f�@��x6�8�|n�#�(�$`�f����\t��w�{/,�(���mE��bUXL�:W 򸴻J�+Sg�YH9Ʋdw�N���]M}������2L0E�^�;�
Y};�}�`d��Fl0�9K�x��,��L�gz�m,���nJb�F��]��)��{�B&��7
��+��k��.�x_��,���$^�5����@�����_m���/�t�)�?�U��iہ��U�L����$%�����
0)�
匹�=�؉��țٗ�su�)�˥ֹP���?*G���[���fzaԄ�4�BN���q��cp����=���|��%�e�Y(��"��M���s�ˊ�&.�#\�}ܻ � (�6�-z��;$2��������i�%���'�Y����|��f����n7��v3�����Vx��e��3��pӵ��_0��3,|��}?lg�z�>n�5��~z(~�����N�Z�q)��\r�\?vim��a�lN��E�H��Vn�܄;��:s���Y�֗{b?�\��z�q��<,KĭC�-��p�9{i�f�%y�<��ǡ;��]q.�1�[�M�q8\+-��7�p����ܴ�z�����(�`{�*,gx�
b}��|H�^�s�h�����I�z4<�}��f�8�ޞu���_6�Z8 ~�/DWY�W�[�Z/�ʥOJv�w���,$R|�K� �C����fe%EK^ָ%��؊5F�b �����qA�cARIH��eR >���-V�樏������</c�����u>��J
�>�v[C�_c�y��m�����L���Lo�;96�U�ҝ�@
���ϵ�!�hy�ÑϹv��gK>�>ы���vi3�*fX�m�Ng�А���xmj'�z�t�?_�ΞQt��7�w�������m=C^7��o�M:�@h!��^�བ�L-7�'��J딫����~K�
��*3�F%!Jٟ+<b_�$�ₐ�C��N n�i�����If��{���|��8T�&` ��k���M��er�U�;T���$��v��U-���c�Ǌ`��Y��|�ǦС��{��x�?���,��Q�MP��2�'?-�܏S�7nڶӨy����N�u�quoxe���XF;��!��������3,���W٢pܩT�tj9�E����gc(����QX-Fe��dm#D�#pҦC��,��>�l{EN=ն�P�ym۟�/�I\��Zzd�è�:Pw�U�{�ST*O����B@s��)�%+��CG��hy?~Y�-�K�v��~P��S�yϻ� ��y����M���y����빅�G���o^h��J�^ fn>�҈wh�.�}k�2����rQ�w9Cd.�=��e
i��#:�Τ���Y�'�Ӟ��>~2=սt��y�l�QWt��R@p��#��=_5�_O�F����^]�p�S��t�d�]���D������]��g���K�˝v���7�zx����X�w�.���U�L?)%�\|L����l�Y(�79��ž�սSq貄��6�F N���c��&��h&UD��r�s���W��6���ݾ�%�Л"�o���(�(�}�e=,U|r����b<�Q7 _�u���>l���B�	�;j3l�|"��@I��������l8r��<���_��E.����H����E�57u	<䀃.xe�*8IaG��G��߹�IR�u7�E��Nq�K��m�d(����P�b���滋�U -�9})�Ϯw��+w���z-��zQv���"0�U�]����*O�/���������9�Bb�^�h29���6׀^3&cD�tZ��?����NA.�%j=��&8�f�՞��̀8Fx8��n�$����o��{c��<e$Io���\+��-R_F��7���R��R��Ey�mR,��2�:]a�9^D��<T	~"��ƻ�Q���Vύ6��1������ڊ�S��z��e�]�N�D�usS�{�mz~����fҗ�-Q�d��7�-��&8�^��wB����$gI��5�[֧�&7��K��RnΑ�G���#�y���Ɂ8��D����Y�/z*���5� ����
�x�7�r��L���Z��r��"vXj�NЙ�Ij�*�'V0p�=7B��:������k�wg�����x�M=?�{���굆��H,Q��E/�F�W���@��N�SvjLGߥiʶ9���8���Z��(���c7��T�zU��gk�u�</�O�����&�(�k4���:i�IR��MM��xy����q#Jk�:����ɟRr㹁��*<Wb�b��@���M�j*��*~q���}�}��se�dY5��k銍<Q�םwr4���}��(�,��@ܓ�=�K�H9-`Ok��@T_������IUۦ�%����N�e��(���{��~{�_x b����p��f�P���F W�%��	�q�U' �UI/'��}�Y�ѓ�&���&qB�ii�����0`2
��% YDocc"ܭ���h�c=��6���#���å��4������W�Y�K����1"R� �M��֐��<���s��	.��?؟�:?4�����o�p%69�^yo3�4i���,�����s�m���e�Z�#<5Lv���^/�M����8TF�(��0�!�5WM�����aױ�D��D�׹���`�"4u���>:�v����oI=/�X'�J�D�h��]*�Ρ����g�	c�f�8����-�_�����G�o�-I_s(im`��y\��U�ə^q,�'�p�|{�n>�"
�(8~4��m��<�yd�sp�r��(�6A�ueb��!����U����Ў~��'	�!�T���a%3�����0a^u9��$ҥ�B�ܟ=� Mv�ȷR;�S?�� �JFC*N��6�B����:�-��9�#�	�X���5�()ť$McA��&�Z�b��|�K@��3{1}_^n�s�;��S8�$�/�ܙ��K����!i�>���1ڢ��Bt����&���x
hR �zˉ�����~_]�c�򽾠�ڼكݔ�]���G��4S���vs�����H�-3o��(5�H�c(*�'����8+�^x� ��O��~7�U��:�����n2�:�d��^��GM�=��>��3|g��_ܺ�bp����[s=�Xdr�t��zOZ�P֬�:�R֋����Q,����uW���������Q���#�]���h�T"���Q�_Yb����:��J�p{fQa��@�.����0�����@Y#��n���������y�N����o���kgM{����c]/Z=I�ydO4�R����/5��q 6�L�b���4r��A���t�J�Z]��3����o��f��v�����  �>U�ʆT��� ?�</����|��}s��2'G#_��x���|�ݚ�gd?�^��#Th�2��W[2�d���1��f�c�]hb^?��[M�� �����v��}��E'O�������ǩ'Iu������.�0/�6EL�팝��7���.7(dzY+��.�O����-טzrif*�o�ҍ�C��P��O@��}0��;Eй�w�.e�>���͵�1����>�7�:���ӗ?n?������9����.��D���c��,<���^����X�
J�˿��J�4c�Iг�+�$h,V����/+F#��5�j�%T/r^K���â��@��r���B��t1 4�,0dw��$�.VGؽW"�ksQ#���j���~��sn�_�Nd�4�f~$��r? ��O�m�#����=�b$�W��5<wٮc�I���Vq�R|� GƯ&5�X�X�;B�L�Š�w;W���P���G����0If���� =��n�D<�d����G�/����տ�:!�� 83�M�olx<w�֯�2Հ���y��=rt@��y�_�^u�H��Jm����a����زCR�Jț��z����J���~�ez��ΆH�k(���X�4P�;�/��:�͓	�*�;����Y�(Te��K}���Қ8
�@�8����ea�[`Re9$�D-�VLr�����+Z���Ѝ�?�Q/�b�%w��0�,�^mg.�J'g�O�0�a����e���ة��ϭ)pF��S�&&���T�Σ��sY3��1g��J��g���?Eu��B��3_���3�j�؅��54ׂ�P�t:���.n���E��t�6�;�c��G*��װ/��Yc �87���CM��Y"���}���Mu���<Sf΂��o�0Q�l�*��Ֆ��d�������%�ۀ�!���j\�=1�䗋��U��[�`�IfM��VVD�⡰xv"�v�8��zi���^�!mB��mtqj��W��r����/����%ޕAxZ���f:�p"���Xz�M8��Ld�xz2�:ņ�v��
"|{�3��q��|����(��d���2Q��Dh޸5ڿ�	=04�,�Rj��/�s�Y+MU3z����~=z�$���Ȑ|�<Q�j06%A���U�b�Nm�lS�t�(ea�����)2k�$�A�HM�ͫ�1�{�$��A�����t���� �0{��9�h^����e\��SG[;��9�2Z[��X}�"�,6���>9�Ͷ9<Ј�m��bYL���*��C+��;�>{�;�L�nikC[�+_K����M����U w��1��gQ@�`J�����:�����z�dMW��G.vq���,��COaX+�Gg���vt��b'R��rd? �ܺ�����S�w�s.�T�Ki�~�,���\g𖥲"Λ���	�'�Yֺpi����iBR˽
���
ə�c���_W�d3��&Hxy���"]�2R�@�G�4K��*���mM7����p�S���H��a�Q�����wh��kB���B;�]^E����Jc,�8Cy����PVi��F��?��O���jm˯XAd���{t}� ��E��{��m�u�/ ��K\6�uo}K��3(^m�FF��~&��@�K#g}G����F����;kQN�V�k�0F>�2����2M�x������q��g����?��R���fV<"�X`R�C�%��x�x�XQ�xN�c��hu�6�Z���}=	��6�צ��+��)��G��ɇ4(t��A�,�Q�q�8���Ԏ�6����g�7޴�NG�ƞx��������ăQ{$�L�y(�S�;Nc�r�e�+��ix��[:Ys����Q@��%�{b��DWeʴs�G����-�ϙ�͹MX)� ���x|=w��ʴ��'��;�q�B�9��v6�������I��1Z�������&��܀�Q�
��VS�H9�#�:8�*���H&ګxdRP��`�ĆJ���ܹuevE`MH^p����a�����ɇT�~J��c��6�4v��Z�"��d�n�[���E�<�3� �=7�zr��䵏IH�� K}��R����R� U!L'6i��'e�ʬ_Ub��HdbY�����[ϸ���J}_��vw4��r�@��^L��!L�]bV�y��;�[f�5�_C��OX)\�%K�Tg5��Ʃ5؀;�j�/;����Ǉ��\�5���l$��\��(�mY�}q��@���yf��k�9����Ԯ�[q�/H��g�	p�@;}o���I�'}��)1��>_�Uڄ)�$�W*�^)<�^��J�P�$d%'�������(Pȇ1��K��"�P�p�R�	P4	t��n��nT��O'f �H4��B��SF�z��G��Gm��T��Bd��pt�N'�C�8m��0� �;���zG�'��cJ��J���N'��H�`��S�\VX�o�C4�6E+��L�
?,7KdֆV�N�v^�b~	��'�iق�<�E4��~�%dVN�qx�[�b�i�[�Z�zY�n��[�X��#`��׭����-��p��O!��n/Q�_�P��u��&��(�;r�_��w�U-_V��f�n���X�^�8#���ݪ$�l�*�l�=�;S�U��C�SUWM+���)�z�L��_�cAK�ba�ڋ �^�	?��87}��h���w��f��G�"�:e{��zY=��un���kv����	�����9ˬ���؂��2����>!��A'�Ͱ���gѳ僻�Ľ��{ͤ|�[�Ξ P#M�$��{,?�af�G�F��:��+��3)p���,c�R�B��>&r\�)ׁK�J`)��7���]l��Q����h7��Ua��r�O���:-�Hn����:��e'�R�PH_: dP�QI%LU-�vTQQ���SCl�I��H
���(ۋB�;��=�2��v\:]�o�������^��Q��hX��@]/�S��ryl������8�>Q?� _��@����!c�ӳ���A	�������S�2߻��w�����>p��S���,T����p~��6y�;Tx�ԇ�[���c"��Ù[�w�PU0��N�(/½x���Hz��:io��$����&|���M`�|ec]Z�I��5�����L�ǚ�Wy`<LQ"�_8h%=ݪ��%�X�и�hsS�ƻϖd�F� 9U-�3xh�no>_�y�%� ͬ���(L�r���VH�L�����)���{5�.`�7xè��j���H��[>��~��n��u��D:��O9~ct#���yU��V;/�~�~�b����$õHi�;�&�	�H^9�n�v���Ean"�k7Dn�[�+���ơ#J?�鶥9{V t$�&�r���{�?_}��1��1�J�t?5�m�s<�ɍ� ��_�u?O��&�/�8f��9�O�P�G�|������[w-�>�M*S��D��T�7'������%'X͚��2�F/z��w~����m�|a�n���?�����>���,Dk�uJ5�qO*�gz߹�ѹ��W��#��ɇi,k�:��[D�Kj<�)OLEx�"�㤤F4��Bc��1�0[Q5��4L��e�^7���_����?mg�REbER>�w�bDz�Ė[�Wr�Z��C�$���>��J�+���٬?�oIq^��v:%�7?(#��lh���|PU�2,m�����c��T��G����Ѣ�C�akD�Y�p��ܾ��8af�hH&� �7c�u��$�޾��迗��z�j!�!��^�`����:�и�tC$�mY�d��CqT5�$�u1�_d%Y n�䝎IdN���&�ex�M߱�rk~��A�lŜ~Ts��&�GgFd=I�&E�'HBg�����(r�-�[���K̔�=���65��JR��;�k5yAϝ�=]�A$�f�X��rk�z`ͼ�R�I�ME�)~�l�<�I��d�.�LV��#3_D���Jy�&V�[�m|� �y�����C�����"F���C��;�N+u�Z��Q�H�ᄷ18
� =���hk�  �3X�^���f-LǷ��L��p�E+���H��l�p9>ǡ7|՛P�ȁ���ਢ�:���}
���o��WW4�.Jp���ߕe�i���xO�8	*�n�./k��jH�1lt�������D�CG%��Bn�C�ꅉ����/�=f:�<$]��Q�2;.�|.��] �i���z�de{A���X��4�E�}������y�T/H��p�P�I���4/��q�Iݭq�%m$T�GT��^)s��{�:����L���#Y�0��Y>�(�ON�<�ۺWU�ĥק	��90m+�]̚�}-}�=��������!����O:�V��k�鄼�&Ȍ�o!��Kl�4IF�0�,��y�+�ZȖ��Y]U�������!����o�.��g������.=��b�%-R�B����n����͡���*A �� ��@��Ѥ+\Ƕ��+q��M�RB�0Rl�W������n` ���'�?��mݪ�@�+m���i���P�bf������TQn�ͯ0��֯w����*Q�,h����_�}`|�ۼ�7�H��i�	���Q��wj��F&����g?g���2��]~�.�p����z8��y{Y�VEH���H�P�����s�Ǘ-��w�Ӭ���vV���`��d� ��.�Eby��n8jeZ�~JX�M�	��UU��QQ���N�i��C��!����*hWA����$S��ʲ���G�BJ:P#c�Xaj��[%2Ux\�Aɝ��l)8���bO�
4�� �DY/4O����=��I*���F��f�+�����Ī�#м�θ���]���*}���[+t�R^
��Q�(�a��b��o{ �璽��J�	��57��	�2݀�$M� �:��[=u%�����Ý!�����(j��9�6��X�R�/�D#CDǗOr�),Q�WnN����*|\�zK����qlڡ�Oş2d�S<]������B_��'��	�AM��?�� ,J�w�0�p�B�{3����|�jt��B-WG1�s��ys����K>!�!+ݒ�' QQ,���Z^�:�c*A5�g�����s�k;d��Þ��n�?9�����.L��2��ܱ!2�l��ǹ5�ҚX��.�S:fD���1`੮<����
EZ�_-�hF�j��Z�z���yO,�M�o�4�d@/<@��-:�磬��W�MA_�SӚ��מB��Gb��<���<���3��սj��r熫��L�d�y���ɬe2T=�W웲���ސO=F�����m�(u1?�i�U��:����	h{�YN�.R�lS�K�^��9�{[4�?�qHѦʔ��2�LYl��l2#���u��~�]��|����m;}�nyߘ��0��OQ�Gq׃{C�dmN��;HGW�]g�w������|�9��=5te��[�Ht66R�O⓶4��/��D�ۤM�����Q�5~�V��4 1�'t����57�R���_�fo*H�<��Kf2����h_ȇ�h@j��$	��j�*�r0�f��z�Ki��2��:ʍy��7��!j��nT�KpP�[��N)����tV4!�-+��l ?�e�M�Xl�;�ܣQ��K�f��#9��?��I�q���F[��7FB*���h��w�h�l|�gO5[��c9������WQ������n�?�iD!����u��'v��A�v�G܊�����S*ߎ�WիU@=�;*�)JJZ���'sς�"�z4'��G��:�^xz��7��D�n� "��t	/�!Q8SBCf���D�o�L<΁�m���=�\��.}5�\l{��n��J�Ʊ����ľ�㇍L@!V�S�:���bI���Lfx2M��)�"B�#�@i��# ���i"��PO�3 �0^0~���u���&��"����'��[���mu��?�x�u.�z�m�vE�N�K�_�<ƵL�uj+�Q~��#(��"������#?��p�8_�[^L挆�{HJ���J�p5��d�hri�{ͯ'���~�Z����S����4T�P*S�AIJ���?�;�,����4=fvԮ3�.�LS�����{�"�1Y,{�&m�M��N�j��1o~���U�Ӎw�k�Uag���l�0S ���)8�Q���o�>��!��v��UvZ��$��{�U���u{��{c�;�	�oά˫*��v�UU/�9�qP$͋HpZ*f���/��W�|�F?;��ZM��z������*]�K��Ft��5�U:'Hc{m~��O���T��e�^�}��c�2/�������֌�He�o��
k&�A�]yʔ��R4����Bd�:��Nm�U:O_ҙ`��E��7lE&�>�}�"�(�V �g璆��m����5g<�2
���>/]�B "���aE�#%xqq��>�U�t��(�92:7>�;3ه�`�)i��ﰬ'�T��^ż0쯯�Yw�d�U�r\�M����g���aqKdb{3ܪ�31��Zk���	��O�o������@Ҷ����æ��҃��T�m����#���?��c�Ne�������C9�:|09fG9�Cx��Ή�d�bL��x��ɘ��h��劒�������RN\Ö���M�5�B��ek�����f�E���h��ƻ���=T���&pQ�O���^��E`�ڒ�Dhb�6���;!�L��]㩟�;�:c�n�H�����rc-z�O����R5��X����d)�E���UY��!MT�~���~�����
�O�	62���%��T�[!���t�c�$�21�w-^nl�=�]-�y�`� 	ȩ�%��8L��s�����������q^9\�(�<l�]VH��ĝbc�7�����V�Z0ϙZf"�s����&�����������5���D"r�����@�˯�FO�Q;�%� ��|����\n�����`�{~�h�y�_	C-ĺ�D��掠�>���.�Q���3��4����!/��]N9ɡMB�]�����M��N����e���پfQty����� �]j@pk��k�ջj���%��)�m��{I�����	v��U���S%�޸��`�?��_��
�4ˉ5�	)���t.R�U��\l��zp�0��d�o7,������ ��[�u���/ ���u�-���X��o'w���^db������OЬg�G®L/�D��T��N���J�,-��4m��}�pYȭX+A�$pb��[S�t)i��]�UV�^?D�"�\��]}��*��ChV�Rh�M��eo����_��Omڐ��ꅈ�B%����:�<[oߝ�?GF(��X�U��9\���M�%.�.=$�3�����4Z�j�H^���}z��>i�����sJ7.
}\�gJTi&��V�
4�ڑ}�P��G'D�9��f���7#c����|�3a����0J�I����A����esO�"��H��g�Õ�<��OV�0>�3��5�����#țҚ}��(;�3^B[�Vsb`Io%a�Y`�.|��X�4��j,��5�h4t3<t��ݲJ�2��
._4��i6�ȴ"�?<oJ�|%��p��s�hzl8Hտ�9��o%��aRC/�'*�a��L{�I�~������8��o+����4��D��b�3��2�[����N_�̣�('����#kO��w$�Qi}���Pt�@�6
8�EN@��ۮ�2D��n�����2�EH��V�f�r��՛�D0O��1�5��0�W�1�ڌ﷨|Q��y���^����R[�L�o����t���a�=fVP}@CT��Q����}���n��h��y��$�	�b�Z�ٸ�p���k��3�j�=�%$�2�^�~�_�r��۝��8����i��A08���k'��M,c�����R�G�`�~�b����Źq��~,nO�?���)s�;Y���*�L=k�K��s0�bD:�d���g�-^|x拤?��)k�s�<3X[V�^��Z?[eչ+��fo#�pE���eb=���im�,j ����*�o��r�i���E-��>Sߘϼ��SZ�ƪd��9aVg�Mc��М�\�h��GvWg��.x���O��螚ޟFJ>r��4��o���'�۰}��r���!�͋p[�#�t��KIS+��=��8&�ٲa��ϻ)Bx��u&m�d�\�/u��=;!>��Ρ��iO�_��a	PW����9��G��/��/6���������~�9lM��B#�&o5�b�ϻ���j�,ɍ
`y�kub���f-g�x�JX��=6�7"�Ԋ�yk�/4��H�8��^t�ׂ?H�5������G��<�d���f-'������1�$7	�l��P�/ĎxܟRM���A_*�5��.'��Gջu����t���8a�	����q�C��4�x�"m�;�i���u39	�=S��2L*ʷ�E��j�WB�̱Ӌ�"�PI��o4����wG�IsqG��?Ma;����u�8~x�+�Q���*�/S�Ž���`�CcOʦ�ʍ����`Y	�Sm��ۘ�۟޺���WD:���1vJ�)�E�^ ݶ$�	w�������������j��ɟp���� �Q�v�Q�J؂8;����2#�
�s3�G"2Ű�`|x���F��kx9xe�����ޛ����#��r�{�K�Q9�}_D��Q�`Y<A��J��"�+Ê�;3���ts7�.gT�'�Ҏ�q>-����fW���䕻��ѷ����Rۅ��t����n7_r�~��>p~�>"�'^�rO��{���oB`�:*+�9v8�m�e�k0�gk�0�t
F��J�����!�v;�<ԩ��(e�؎���z5z�y��Hߤ���멩%�����	y==�N��e�a���c���31�0Ƴ]խT�A~d�f���KR\W�[�����-��lӂ��_^'aa `�-	��X�oW��ah2�R���`9������E���������We�_�O�^���M�x蝹���\SB�a��ހ���O���Gϣ�W���g	�������Y�N�W&@ϹZo'@�����s������#lr�|��fpB�� 0FZ�q�p���V��`d�'KX TI� �ztu]E�"�_D��է�|�[J#��!����<�c�f�=�W5<z}T�fK�j>��C"L�7^Ōʫ@�k�gN5����`�y�V�(�B+���
Ԍ���uT
�>�o�j��0�z`"�9>�OP��9��d��8�?&��!����(�HI�t��t���tJww��%� ݃tww73�0����~z�_��Y߷�����@g.0��z����@L^i��r1�p5�,�F�a(�[:
�E��U�´P�Ie3h����Ͷt��8yKbS34�w[7������S���R�j6�ay�^[�����ۄ�:��2J?(�$b��������t����em�й����8sm/l��Kf�l�\[�1���0x+��������.ئN�+�b����jO#"3�$���e��[}gU�4@Wi��Cx��)R#�W�
h?��I8E��xJH��Ă�X>�;������!3��?bX,w�Z�.-y���������!�[LW������i8�A�	��C���;-��B�n�#���X��&]�f��|�*G����9�Qi`!C���C��|���ROϕ�L��c_�7�?�>��}�PR�{,g���z�}^�F��X��x­�qn��^.5��)��ӽ�Ī
��$��eI4.�[E��a�	�rA���
{�D6��E�p���������.�iH������ޗ{ |��s�C�b��P�v�9 M錅w�3��;�x�T�ti�r�\tj�*����j	�����h/(G�D,�Gi����R�v`�XrZ�Z��˚˃�z�\�{-��-v����$����>�֞/a���C�M��/���ærl�8n�}�08oM^b�ꝥ�ּ'�#���d�R�'���}%���؏%`To��LƋ/�w�Q��&��4󶣯v��0����ks��Y�o�&��*~��,h���� ����$��lg�*�)�{RD��mU�S���r�ޛ,a�R����??�w�Z��)�GPy���$��-3��lV���X���w?�%M�bi�7�Sl|/�-��X�����	��K�2�B�,�꺆���vzl�p)`	mD�r��nG�L,r�?��g�y�Q_��N���R\w�EVP@�Wm��"� ��Xߦ�)��Qg��/�o.*|�z����6��g�'^�\��_��8G��\n���O	A��Y�E�ȯb���l0��R޻��R*4��22|t�s��Aq{�&1/L$r�:i��g����L��]�j�cYjU1�A�0��7L�(���!K�s�l&��f�sY�t(\'g�M�B4�_�"�6]Up7»��&��\�s��e�lK3����S�N*�R)m��Q����ǧ���B߫�ʵH5��������ܾK=DJ
�O��`b��͌:}Q<��zm ������ߴ���`z����ۏ���8�:y�'�H���N5��G�'{9�Tg@亀��3��R�����hD�37/]��N��MM�/����S�.��*��X/t�#~ɣ���3����y����0oEO�[fx=�C	�ޓ/����"g9��M)���7)G��*���>,���"`8������<ym��I�������e=�����eF0v�ҙѻ��wt�Z]�Q��=$#v��s����`\�r��ۿ"LOz��s;;�ޭ٬_.�� �HW�E4�zE k��m1��4��!8U���7����J�����Ao煗;
�nv'�<�tJՕ�$�0C�ԃ�;��^y��w��Xi[�2]�!ю�/ƭɍ7�C��x����̸��B)0����z%}h�:T!z�m�L�ƒ��g�/�����u� %_��0�K���[Gыw�4:���0WN����G����h�j��k:��7Mn������ee=���ֵ򪭟��v:]�{P�P�Y�gi(�w���v-Ckr�3h�{���}��^w�n�9�����SRTY/��/rCq�J�mE��Q"?;Q<L�d���$��GzUۛq�r�Jۤw,��K{ד3sF�G!��x�E��øuu�B����gvo�u�f�"���Ӳ
п�>{vETt��*"%�դ�;��0��M���t�a�D�<�_�Sr��zGoڃ��ЋF9���Ani�����q5�,qQ��m���igV�h׭��[�/6O߇��.G-� �=�8c�;i�U"B{���R�1mq�r1wнIp<��8��z��̇MhD�$�E{��M�T=�$n�r�K}����mI2u�DM��;��n�����ĉ��1�BY0�\{Ǉ�:���^7'���hG۷��3��~۰�X����M�(���<_�d�ό��V�ilK�W��	�a�z�<ob;�_䂟P#H�s�`��m��j�u�v]�K:R�qj�E}�.�D��U>b�QG�&�xI��4�c���Z���|!�Ȭm�ٳ��$�lA3.�̎��ig]�3kGܾ2F`vO�Bi�Ϸ�K�H�墡e���i��I<���'^���O�.sr�sJ�"�#s;��g�%3��g���5~�8x�@7ý���3�Ł��=mi�T���i��7����V��OT�A�fږ�L�������K�D��䎩�e�$��Gp�AtcT}�(���c�Ÿ���җ�ѯ��ufSh�&=�Y�aOx.q:ɘ�.�m�˿��v]("�Hs�Kh��&���q��[��ۇm|h�t[�pn9j/V8�7U7�>~螵8����������I�y���WX�L����7�3�k��g��B�>_��)��YU���W���W.�y��4낼.��l����
�����vQH����<,ꌿˉ����Y�y������"��w�e��ٶ�x<����F�_M �јh�g����xKN����^J�ӥ��u"=�\�[ �8B�þU�[+|������x����:�b!����d�Lo)r���N��*	�km��B�G,��sU$�쒐~��]IB��[72}�E��Hp�}��+�c`agpv��H姭�0�a���Q��������-��ӧ�Z��%�M~�.���������؄W�.���m_;+�/keWV�Z1_��y}c������	�c߳=�Pv����-���l/Hβn�o9)<yRB��M̧?�@,��������x���R�4���==�4�=���ys,�����Ĭ���1�A���k,��wr�(G4͟jjۛ�J.>��jX�On��o 	ew)�2�l�����(] H*H1tk�}�*����.�2Z6�ğ74� f���������ط�w���3Uo�!lS�8r��	�T5��w������w��lI����k)Q����KB�3�0����U�º`��q�z>E�夷o=��@���F�9k�Ϣ��]X65���J�~�$�-�3~n4����b����XY>���֩�O��@����d�6=s�;Y�8ߓ�q��|%�	��H~��C#WȮ"'̆ZY��1�x}��,�I�=b�P��^Y��$z�O
��ү1냪�et�����fD��������P5����<�S�~���V����0�}N�S���~�$�_UQ�P�MXl�0��&?/D��7���'�E��L��jyQw�~��]�޳�&<8����r�fG�<�P�9ц9�GgOj�}&����L�8����V�%�Dg�%��/��̹!7��H	��+W'j�9��吠�RO�省/�o/C��_��9����v���9:���\��[��l�nx���f�Km�Ұ��θ�J�윽�Zps6���~�0�z/.mX���B-��P��K8��w�����J����{�@"�e��k�D���'±��۵�V�<c?�W���t����-?��|a/'f0�)��>�F3SxAf'����4zzC#�U~�r���������&��[��d��\bnU��:�N�0y�Z'ᘓ�?�M��|�|�a��È7ݧɞi*:����>odE0������y:�~��L=a��<�a��4 eC(;:O�k-
�_��L?�Z��[X���W���j1��ʝ�|�]͡Q��h�
�߂p���` ������/�J��!��C��u�������9&����kJ�>�s��X��:��+��T�-�3W�&�0���7ǥ�K-`��7���R�y�����|j����f�V݁��'���;]��͐����
w�� �#��������GWh�m"�u$xŜ �<(��>ҎGM���\����]#*�vQ>���J%ƌ�r�Q��d�^	U��� ����H�un�{�^�$��yE���gE�o�m�7A~^˶ߵ"�;����ON���%M��_��\=T	=�R(�i��x�����N���f���,����IX}�@�s���y�"�͑��X���vS�h�q�}}�ɼi2�}$�#��y7� �}8���������6��5�o6����+b�RF%�7�GE�uَ̅�?b=�:8Ē4B)`�[`�z�������-�3[(�*V��z���b�������ͦr#�!<�����L�<�`�K_���f�V7̙۬Gg��/s�o2��TȲ��-P���_�&^u����=��P�!��Q��D���Ʃ��K�N7��0N`���k���E���숉����Pr���w����.5����Ұ2�:�#��ʳ_d0�1-�����ph�S,^�ԉ�s�M���"R]B���3t�e��<��V�Z��U���R�cmj�Y=~<5b��B�xl81�N	��G	8d[>}N�ݮ;���6f?ա\.e�~��&N6�&v���54��%�j���,{_ɿE8�b_q>�pb�8Bh�k�j������u��F�d����P��������/K嚱aJq��3]�m��݆�=�bu�6oyn~I�Yt�J1g��pr#͏�)]b�3w��Q��X����0C,�^H3�gN.��ؓ�6s@��J�h�<��OO�=
��)�v��B֏���ּ������X��-��z��}͓p\(�g]E�;��$��L�u�|3��P��穲�SR���i��C�K $�׼�3��h���u$�E�s1�{�����q��0�dF�Z���1��Ѝ��5�Cǻᦒ�ض��ű�/�-!^���M�S4Ţ	I�H|�ƛ5{O��C5W��yg6R!M���]k�%B�N����)z/{����C�w��)�*m�Yc��w�g��hv�io�����A��g1�����$�o��
�5��=��-��Z��!�|���7}������-µ��M,����lG�n2�r�.����S)GxW����g8�B�Au�:w&N*C�=j�3�Ju�;�uZTx���4��%���t�M��4}��xÞ�ܷ�( ��M �����%�ݖ�~Y���|�+�)�ꓫ7�Q��G�a�Iy��5�����5���}+eR�x3��Y>R�D�p?�M-�^��YNUO���z6�%+��''#6�[�WW>�4�4Y�,Y�e�)sYC��3�ظ�K��i��X/�Ev�f��c@�P�������O�{Ϸ���'�Y�4����qsd~N6Oܘ�|ˣ]@�{U���\����e�]*��745�?���K��n�.�ѡ�|"��������rH�I
��?�z���	��O�Tv��Kx��hO���0���nI�,�Sj~���m��bd�'{�sx��i����5���0�9e�3d��L�%,�>ug�Ӥ��β	�<��@h����^���$<d�{!H﫭Vq�����ل��Ek���}N�"/#����{�Λ��P�7�F�X��_��&�QV2�������'�z�܃x/=�{�#�7d��x�gaΉ��7+j�C4љ��|��~[�u�a����F	#9~�4���ul�{Yguf���#l3q�X�x����K؋�5��id����#/u�H(⟯�V��7RW�$q>m��
|��`�E�c5�W����ջ�6�}��`�����z�W�=>k�1���p.H�R��y>3�IO�VՋ#!�s0=ش�j�}Ӻϖ���r[��&�z���[�Z�+���k���v2��왳o�l�� \Wi{��i�y��D\7�:G���'��d�:Ud�|"�	���SQ�ýoӬطx5�%aZ�M��q�I*c�?��!�e}ڹnHӱ��n�פ Hp�N����v;Z�]+2����Q�Z� Ȟ*�x)��`λ���)j,�q�hj���Id%q�-���_5��\�'���^�(Sԕ�?��^Z�m�Zq��_A=8Z3�J�����kH���[ʥ�~�yF�j�o	"���N1����r}F��;��-S�Q��d^>yu3�	io��[x���9h��������r1�s�z��eMOO���Y�VI�aj�b�!�6�jkJ��@��'0y��H��3zZz�|2pM������$}�k��~OPh�u9K��J!���˘�ߦ�B?~\�b l�YEJ�N���|xo�W����"\����82U�[�[*2�Q�΃^�F5A�Y�U䠵�"��~_g���������S����Kt^�ٗ�N��d�w�#?+����@}�����8:4�h�ѕ �������o"H�$�h����.,��5;���,֒�q#�����>��E�멑}�$��������gg�_���ࢄo9��ަIsp�\��]�[��UT�qx�KAb*
�8>F| ���:�4�l�J�}Y�TgB|��8j�����Zu~�r:��s-0۾\K��������ۜ�㫫m.N�C�!�Z$�����~�}*�{j�෍��|ͳ��V��9;l� *GMW�y��=H"_UC50�tl%nK���{0{�^��sOƼʥet�nɕLr4p�?�: �c5��+�Aۜ d��*˓vh��VNI.n`�jae�����5�Xc��.�nO�c�">D�G=���e�\�i�>����������a�\�g��Gk��Ⱄ�}EA*��p[Q�=]u#�.j˧+���5�2�\�@F�F��՜M{���v��"_;�K���$���n�N ˎUQ��!�l����Se�����D�����P� �!����ye/n��S诣��7cK�a���#c�- I�_��{�ر�cnf���VCI�]��F����K������tB�;��[�/=�H��VW.��ܫR_�yxu� �V[�]X���5��_�>��'�MU�??G�nd�-����~�8d{R�_�����S1���:cph	�W�G2���Ԭ��A��g;Tѫz|��l����Ys�I�O��|������?"+�j�}����-\�5����{�����s�n���A�%��VT���-J;��F�A|;Q�,x�X��|7%�8h����^[G�LZΞ�p�EZ��Ȉ�<�H &)9z/�{����f� �#+�'%ʃ}l3����}�JK ������(-�tOi}哏�Q��+�ő9�@>ވ)Uś9�ĿW���`�����<� `�Xgi��x��?Wn6�X��3&�}zN�+xr	��^�׵(�sσ{\t鉳ʞV��hkz;�)��d�.-&��:�N|�*�>�K�=B2��lj���N�uTֶ֙@�+���|﷢�c�O&����Ȼt�F㑑����SZ��/tVY�~8_�BSj��Ν�5�w�L��J�G�;�u۴<��3���:ϳ��֮x�z����>�OzQ��=U�����1�����F[�N���{�?	�|ׅ�J�"��(cϚ�I�&?���xᡠ[ue�x��������$��:���C���b+s`��R8T��u���"�*��n��@�T�ˀ�+mgֶ?�xp̥�j"3Ŗ��+��w�b�ˍ>�Kce�V��,&�f���C�l)lx�V٫���l'!7B�����5��	Y�F��"b��K}/"&0�|b�`:�KVj��"(��J�]��k[��D(�R�$���'����I+�P��߳��Y���`�M�P/�l��H�2����y��)�����Kz���B��:�6�L mݵ6��2m~}��oJ��0y޿�+����r4!M,�`�u�q�XB�V.��u�e�u�l>+��z~�\B�����qMc�3{���h��E�����
��p���'f9�ʅw���q�A4���-x��^n;�,�y{��@aQ�#�h[�%�O�pn�iP�T�և����x�����sF�������'�W]݊�^�z]�J	b�&xE� Ѧgʳ��[�8���5��4Z��$�G��ק�99����Z7����}@ΐ�)%"�Sa�+��>��N��0�d���0�(���s��CϬ4��e�B�����4�+�$M'u9�x%~�R�i>�=�U~,��鋐��Yn������,CN�����{I�rX
�y�&^�X���~Bo����FPl�D)������}cm�sS���t|GS�����p��M};&�����R��s����I�#��)���qn���s� .쉤�v��4$^T�����+�Z�^z�0 w�j:5�gk�sd��<��{�!l�(E�m�p�Hv����Y_�l����Snjog^�^<�z�c���%��D�\f~��"�@�ֆZ���P(�_a!����9�U9'��&��${FFU 8��\7]ז�p�t¡*=���1Zg��ko��jK�s�\�u�Poz!ۢ�ǍO�c_�z�5���n�	z�*~���,G�֎H}�>ť�3b|��{'�M/�xo`������f9xRe��N�����qt�+�b�*7*�2�$}�T$�b�k�	 ��=�YE���e���[Y�e���+}3�=��'�8�ٌ�ѧ��E��>�9������X{[�d�5����z���U���'���T'魟W�4l�ږ�dZ,�\	X*I��Aj�����3�G*ޟ�NXXT�_��*&
���X�ca�P/��(�}m��ڥKS�5�>�jY�م�f%bo���ܽQ����+ 7��i�hM?x�V$�`r��Cq|�p���h���Q�m*�����]A8�����Q�dz,p�n��k���@�#ă6}�_i����ZXKGxgF$'�mɠ(Ϸ�Z�2��A�f���]�{!u*"͙�`
�*��G+�������ic���WW"�G�o�L�L�|؆��M924��TKY���3�����(���+�a�\S�r��Xhi� }���a����<��*������;�Ǯ�b����?<E���f���z:7њ�߿e�ƍ�<@��O47�r�A	�"�>ș�`�����Q%Q�u��֍'Pj0-�4�]�m�iC�����r���'�J�!m�,ȁ=1trM�ʯ��K���xop�TR�x.#�m�Z͘	���vn��gY�}����zw���} ��z�\i�f�QU����0�b�\��w�5�1�����O�]��0�kA<s�&i��щ+��P>��#�s��#�m�Pdr�;�.�-��5k_>K=ܩ��f�p�ds�z���A<!5��_�?E�(�,�4_�:)���LE��8�6^v�P�Hh���H-KR'q��%����ha�&�pOj����rf˱Y�hr6�줿�7��}��R���J!6Ŋ_�_�?�qGO�S����� ]'z��X-��	�Y�<ċ�#��p\�a�o6���)�m��e��K�Z3{"�}RB����Đ3
�seH�fe��gY��կ�E������5��0=�bX��I��@/�����,��!�����C�5Z+6�4}8�� 	�{�������N��䁑&�z�I�"�K5#�eS*1��d7��z�2.��8���\��/Hb��3h��f�"��d��{�Q��=�ũy��&T�vx3Ǒ�]_�`�����;h �g_
�
I���cU��rª�oZ_��0��yŢu�&vm�k ��n�]q ���a@?Q.\s���Y�W�+���+��{_�w��:&��x�-:nEs�"����f!OI�����ʆ�S���zRd��R�������+�Ʃ��Ɔ��׼�[/7�rg}�'�(�f�n����(C�4�,��Ϣ=1߆�V�Vt�-�΂�u�Qi��V�T(��w*��ͯ���@K�����Bx��sv�t'����aN�ݤG3f=��bv^�!>}��[*����o3��Yd�(�K��WS�睷'��`����
!��r/N^��s�DU��!� �1�����u�sJ}�����'_o2*r�ͺS,\
�j��f%wGQ���3�'(F8Xd����&M��M�AK��}(�ᛩ����]��z�ɺ$s~�k_H+���ly'�#3\�r�*y�.�:�T�ԕf��+T�㉅�瑘��h��c�m�24s\4�<~s�5F��T��S��`Jl%�2ZI���gR��x�����x����Nmu=3����0���~<�X#���,ph��XX5�T%�m��f!̚����C�}f������
����~qOe��zdݒW?�|�N���s��;SUe�r���D�ٛ)���;Ko)�h9�e�DD��0��lޖ����2�mQ��1~�'�s��[}�Ň�����pm��>��+sWCp�w�'b)�#TQ%��w���DM~⯂r�8�X���6���ơ��D�J��w�>�H��� wI�����ϟ����R���Y�ܮ=��L>p���:���xGWdudT�dl�E����u�itHBb�qX?��<�GRs��Sv��	����9�Yx7F{�G�F�9X��3=rH�zk$���;�����\X ��k�jܴB�f��ɶ�X|�#�w��p�'�p�y�G�.�GC�9X�u3��_Ge��Wk	�lֳ"�=T���c�2�)s#[�ݎ,�z�ξH��e�V�4�2��#�"��$���_�Ԙ�@��U�!�j�8I�p;хi��7v`����&����n�-��[���7g'$6���!o�Z�D�M?�$�y�<}ivI�+:#�[kklÄ#v�g���[M�1?����s�y�{�����hWt
�
��Y<�v7�r�������.���-	�,Gmnjs����|�6`>DHUhJ�5��&@����[T��0�8(�W�Y7����g	�IR!Hv�.m��]�;s)�W�6�.��g�\[dD�D,w���b�N!�,oPe�V�j�'�\m�;�l^�=��������^�޸t��!��Ɠi�~�g]�M*$�x3��Ñ1X~A�LPF�kO^^~|5CO�B�AFv��G첦qTL��
�>���:��U;�T�e��
 ���'�DA�s�7媪�.<��	]�4\N��m쭒��82
ګ^OW����S
��,0%M~HHd��x��[K�,����S�1�Vy�̌��-����Uw��E`S��|m��U��S�J�Tn�d��7>b�Ga1���5��/��Zt�û���m��]�M\$�Z٨o�<�LK�;������T�cR�嘊�z�����]�L(��!UW�l���(-��?`��4�=ۜ|yuumQB^pi �v
��j�Δ�\Ս�3)\>4��^��������v�����,������t��hQ��N(�OG�#e3�r���z"�D��� ��J�q�n����h�x� �pl�z���i5�vZ�qt?uHEO��U�].�-�LZ�U�숄%/�K���D�]�����JmN���I�:��E���6��,��/�w���M3 �F|�ytT氄~IV*hX�\HJ��u�N�̃i���}�]��T����y�Z��?����9w�D���Ќ���w̌�@'/O��\�7e��ŀ��V�$S.JU4W��S  ���'/���Q(���)#�j��3d#l��%��1�tu9�j5X��ȍV�o��8��y�.��A47Hh��J&#�"Q9�!^Yf��MV�$��oj	�]�3|��>���C�0����Y�.�D8p�n���}���Nq���;?~0�!�H��2�[���ǧ��\`Sr��U�������̏q����zerR�.-+�8sZ�2^�i�����X )~��>n�<���]�=[O�
1?�H�ԍW���L��,DM5M�ǒ�.%���]�%�:�o�_|��۱�ɚ[^nk�W�U~	�G$��^�2���q���(�5Dg��t	s��l��ӎ�&s��1�?����965κw���̨��yY�e)$�=t���_z�
��P&\9J$X)W �K�]Dƅ���`��)���������|�a��=�;�kRwiKi"�om���$F�&z�ݩ�Nic ��Z����'�E
E)l�S��Pr�e�Q����?#�S����2�~�o�9"�G;u��Z�/h��azB%aEe?V�k�m�I�̳ȁ9ú9U�E�K�a�rh?�b Y��F/>����U}����]dH�=ҮU����&��7���	O�6\� 4����^w�1���J-x�fp�4����/3�(2j�o�݊C���4DFh�� TI+����K�]9J*Y�3�qw9���ƫ�2M�B���o5Zu��8�Ց���<7U�Qo�h�Ñ��d[@�r�*�[R�5��*���ȼ�O������E[�r���`!�䋫Cv92�]�YK7a�:��
����~�������{�BJ ŰU0DB�]���t��h��b�����+փ��!�?�?�bR����u,���K�v����0��#˲8J����V��e���@>�����F�^�|����:F�r���~�S������͌㨇�ڧl���V
�mV{H���M�5�,�tpq�:�74�t�s>�|�b�P�Jk��y]/&�?�������9h�J���O����������W?���n�/�~�ܘ��T9�厊w&3�=�n�(;/+k�V��(�<��.G��]%.>Ĕ�
;Sp�mw�/���sV�r�ӗ�(��tM�'��Ya�9�b�#!!�]�o��Wc>���,3�YOJí�����*X��Φ|���sm��͈�}���ы髄��/�
Ķ�b��"�m�������
���n���oӡ�y�=-��F�"�g�����/d���%6�����(�z���hU�Yr���K�\�,]v5I�܅%/�+�~���0Լ�8L�|���}�E���F}C���s������y�-֗���9�$��<͂5�<�/X���+-��t��߱u[��z�ͅ����_6f�����w�5>�m��r�����X^��i7˥qc��r3���81l{w�.B������w����8B���/�qց��\k�d�'�k2����*--��^���bv�Ȗ�KM�F���������p�}PU��m�Zcl8�Ѐ��Hl�d2~e�"��$z���[�J��/��buL�{{�p%Y%(0�O��5-��}�?$����8��u�<M
��_$��T=u�×}�I�@pNؔ�_N�#b[�d�i��3q���4�O�=1�+�f�#��N���x ����~�I����ܟώQ�E�4��u�����?���<j�䘧B�2�!BB\Ы����9�-$�6z"�f1�����g�,�ym�'�t�bVC$M�=��
J5|��5��K8��X8�wm���7���1=�<kv����9G4� 1�W��м�f��ȳx��9P��^�^Q�"qk;�\�{���)�r��E�eԌ�]޸��3#���S.ӱ�(U{��S��-4��)�C|]
k&|S���ˍ}��lo�h�$�^�Nm삘GXx(�E-���.�Г?S�,7Qn+�A��r����ȴ43�#g���a�(%��!SO}�����x+}��xx��&AC���l�PPe��}h(�y��UX����F9+$��a�h���U��`����
7��NT@��)��r����Xж��'���'k�s.�)7��^-����������3�+{���dB�����Q����"���H�h��8m�{����\������ɕ�+mc1��;��mng%�g2�}:��8�'L�[��Sa��B���R'�W*Ů�J���|o�4�PX'�����.|k*,)Qӯ	���)�15���I�jdr&ڌiW�6:u��%.,ݭN�W曨获y��f���ĕ+9R���[���q�C�4�
�'�+�(�7hƆx�n�:'�$����׌�F�m"4��C��;�{�Y�n���-���ϋg�Kn���۪X�fQ��԰������f���f�ӷ�)���{*u��鲰.�h��kk|�5���"]�F�Y�^�y>�-˥mzM�F��� ��_�g{�1�&'1��旾sA��7�N�"ɀ�o��iz/L\���M�y�Go.u��ʻ#%�G���Z��z�*}�vp��&~xe�.�b~��;m�M�C3�x�C-�Pu۝�W�"��'\S\�z��&F/�nՓ�x�TYN�jG64롦s/Bf��iB�����q��Ƕ�� `���Y�x��z�2#�{<��qNzt�2��c�`T��s���g�>m½B�Mf�+�꣊O�h��.۝��v��!I�%־&��7��e,�\���V�������p?�N[��$��\�"���v��h4�~�`�q��=����N�P�Y��/!�v�5٣���z�ez}��M�(��-^��my�]�wc��[!ޚ$�{S��<�o���/	��/���3���1 ��C��[�a$G�#��knw�r&�7��)j*�q������Ť�� '�����}55Cf5̳/7bZ�9��Ě��U/J9 ;��B� ���� ��Cz˳�_��5�N����+)[dYC7-�nnc�:wv�;Dnb�k:i#ШM�Yl��| 3��4/)V��)�5!��|�KV
�Ȳ����������pR��r"����Z��C!�΄�(З�͢���7?��F���z���Ug(71ǜ�&�r0b��i��:rYGC�W�ɻ��O<��?�[[ !��j��D�y"�BS���+]���ZE/�L�DK������|]���O^LO�t�'�q�^�l&S�-��sV�X)X�f���pu���k&U����=�o׃>*"���/W�c��8֖����"��� 1vl��z.w���W��G���pF�T;�t�\+�H*u�������[���l�3rP5 89���bm��� Xp�[���Y;�gKlr��M�r	��d��W]���3ͧ�����[Y�mn^�Uί��`�+/n!~d�'X(�O1�Su����T`fP��x�<�4N����mA/VW�h�x�&�Bb��3�~�N6�jB��ƌno��6[��E��\�!���/ɝe_���h,�ƈI��x��i�߈�b�mHh��DYPP��K������sK��чľ�P������A�P҅��rV!��K�ioNG=5�gs�Qhh���'㬒�ͳb���m_�(����J��i�%*͔F�f	i����"wr����Y���ڎ��ԡL��m���e|hH�񶶾���[�b���0��Uv/�d��ΗW� �����+:��n���=��};�N��YG˧D�����S�b�Uϳ����'��B+�����7��{p�,:W0��7�������9��T��6�y�2ֵ�b4g��G| EG�M\�\G�������/�!U�h&�cMy����#S���;�|Q�҈�iv���&�&_K��{'��d$�}:��}Ǡ_N��8��GS6�c��ʑ4�%�EӠ(iM|��kX}��yM�r�4�qVF����[�Az�}'jy
��4%C��AY�,��O�o����O�v˧+�z�	�J�����u8
Aed���a���1 �+��᥇��M�ށ�c��/��R�m��!-��b��uN�lc;k�7#����8i�e�m�JA�����h\�oӴڦ�P���-?K	5I�d�f���@���-���@�t�qnw�G%�|գד������-ݧ�����
�%0]�+[%1�����εv��n|�ގ��U�^�U �	B;3eR7:*?g>�}�u�<��˺�����	ā_�J�U����k�$�4l��6ն6gԴ���1+�y������ǂ�=y��k�\G �pǆ�f�˼ſZ����n�g��x#ȟcW��x���p�p��ɇz\r�N��K�;�F�y| y���4����TVH�TW�8�؂�,��f�ț�>X�,���������r"��[�S��	���%.m���%/ϧ��K�pj&�#_Xu��u�â�"�R�}-�Y QX(Mݿ�تm�����`CQç����p�"s�9<������Ib�jޓ^��IsIڬ�,J���6�K���M5�c�ω���3�_"���d`s��&��/�ʟx��E'��<�5WZ�s|�>a�ʮt���]���k�,����I+���VP�4B:����1R���XJ��r�.,�b�x�
�5�˖��6ꂌ��.�G��q�<�?5�H�Ev8`d�+-�B�<��H��8`v��|e*�s,Q�p��1�3=��!���}vz(.���`���$;�Lx�hL	I~MbH[����+��^߰==%)(J
H�Q	i�fJ���c����ь��3`�FH��QcCb0���>�{�����~�羯�z���VW7�:rU�+x��:��b�b�Ɖ��5{!vP�'K��Q>.�e����%�Ek�S�A�ÊW%�_�CLT
t�_��E턡M�o����	��F���Uw_�&�|m����6����4��ܠ�us���v��5P8��{X��?L ��&0�uxԚO�U�C�nY�Q~X�����~[�V����/��;o����=wpT� :k;7���6} A� �*4��[����D9)(��La����7i�B�n@q����\��0>�"���Q�j��Tg�_q,���;ͪ)F�r�Eٌ�>��p����m�E�P�kT�E;�v���6tY%�N��N��GǮ����ue�,OZT�%U��x���=!ϧ�x'2���^�?>Q������	�b�(j:J��a���@zلW1�U�SX����N������]��i׽�Zvz.$��rJ�e�i�� �l*�1޻=I�R?Ϋ'ζ���R� EQ�Y���� Y}PS��bd�NNN-zq����-)q?�r�G�?��\A ���!O����)&z�].�z�_?�H�%
*�=r��>�"U��}���u7"ɗ��� ���na=E8����<I3��ǲ"j��0z���N�q�?���-|��/��(UuO�I� ә����C��`��P��$G�ʕ�~^L���?�_��Ljd���S���aa�C}��ʠ f����vv������	�=�?�S��d���,C��O�� ��xaX^zV�R>"��7���efT	��RL����o��?��}��o
Z��u<������L��6�Q������o+2�Sf�cSW��ӎ6�3Sk+�>��a�[�2�͔��v�y�S�!�����c	���p�����`�WCeq[������a^ �j��8Y�9"��#��s�=�(m�C�*��;/V���1�>Y��it����RN+�E溻2a��h�S�5���׳w�D���gZn���ތ���L�i%������'ps�{1�<�� �ء�il�B�8�"ۃ�z�������c��ΐ�Q��|MB&�u�}����r�dm���v="�U]���,C�g�R�����qs�G?�ɒ*�^P'�x	t'S������'д;|��{U��?��z����F����{���$��I��V�Y+�Q�:�������O)%�\�n��[�.�@�v����i���8ό���ƾ	�{���騵u�C1hO�ԋ��c�(����TFZBC�5�'zϭ(�[A�xP����|?�Q ��畟�sr���_�y?#g˗F��L\���V"����y���[z�E��=-��d�!�e����� ��PLo"3�e��>/zǀ�Á-ŗ=V���6�Y�#�נ���!��m�S�S���9@�Am�Y������|W�C�yײ�.������|
�YNx ��s���l1���J����J�Z,n��U
�gG�t��f�O-촕��J�I%g�����
����d�1gnJ�g��ۉR�F�9>�E�����U_NY��%k�2�:�%}�H��43�Q� �}���s��i`�c�W�dP!�-s%�sP�}vbK�ה�(��� R33�a�k��pHz������G�O��M8�-Kɞ:����pD�oK�]->�,��� ¾@�5��y(���/1�����.���K�d�Tغ�6�>`�
�sy����cC�����#|%t_���I��Q���ƾܘ0�W��M�
<G�w]����
�_����i�Hx��G���hQD�62*�ef�\k��{ވ��q %�R;ٛ���H�Nv��1��KQ�� v
W��_Y��;#���+G��+��9M�Y'8�x0�H�@B�[��+舃;c��l�[��(x��޻��NѨ��޷2c�����[���g����H~�rhu���w> ���rM��O�����g[����@�z�x�A{���N���kC�FS2(�0FD����ߚ�ۅm9b��+�����RyQݓ	���ó/�*9�ꐌY;W�`�������ڪ�J�$�Ҏ��pt�2hJgWQNP�"�n3}��?[����=z�����M��%ԁ�x�ֻ��r�����!G�����5��E~�^B�8_���0'������ྪ��>�������I6����Ш��0�������Q	&�?��'bCF�a.I�.����"����>��|>�6�2�{�����4���X�M�*JȂ��0��U���^S��VU�2Oe�cA�u_��i
q;r�����3%��<U\��ܼD�R9?p���2��'��\�����W��4��%b�zG�B�a��Fpgnj�����[�JF~�����H�U[]��������t�	�c��[���G�!��`c��t�pi�Olu.�	�|#��%����P����pL=k�T=��$�(茴=)D��\��;
��S��z��z���3%"��9��,似]-��.��ZP]�}IT�ճ�#��4�/�q��k9s���#�9�B��A]������Y��B��GJ��Y��)�๎�c�smbn�Kx����,j�0(b>�ڼ�x��z-mՠ�_&������n��;����M�DQj�g�5��$��h~5�����U���w�YZ�?��1,;��u�Ik6{��5~�Q����+%�eW�:�y'�6��v3�`O�V�6oz��@W���?������p�ކ�T��1�I}�c�_9�Vg,�=V���K�L��oA��lk{�c��F��e����L���q�Q������;�'$��7 _d��T~�@8>p��\��R��ދ�	YvM��Ə��C���&	�@|v�s7z	rneB��9J��#��>`�z��w㴐tg��c�Vu���$�[t��Ϝz���f��MW9�:�	�R4�涱�Э�"̲چ	w��Ӱ]��y����)��^��zX�(Fg�`7�EN�����әl�)�4qL����k�J�s�I��,oQKM����/��f�y��:h�~�y"��l����쟩�v�Q���%��{c]7�o9We��Gu�	�������#�'�+��O7��$
����T����m��6P�Sn)�e�t\Y���a�R��<�O�}f����u1w�}1��J�%�'ٵP��AqԘ�����A�z���`)`R��$�j=eS�ytm��t��7\#�g����y�YfӬ2���9h�5���I�gU0c��tvb��)���$�T|����wu�ؓ��;��L&�%��乃̢i!�R��!��?�)F��8�6j^���M�Telp����ie"����\�c�y��q����D+P��7�����/Wp������ͣ8	I�=�� ����ke�*�~?������	��쳺:��o�����7H�RJ�)� ���/���8�Ɖ��kg�[$Zl��LI�ȧ�>D �d%ʗ��6��:~ N�=�'�o�<X�R;�N��;־�'-�b�A������O����4)��Y��E�w;w�u������߇��q�N��x2>������(�򟆶O7$<�it+�N��1~���I��2��2o�X����[�%� `�a����(�-1D�W�;�Kɴ/����ƯY���������J�@��2��$�ï�G*�(q��=��ٯ��g��?�׳iK�:'��`L�3d�Gn��v�6e����rmh�� -��i|9嶼͜�Ω�qu�F̺$ꮖ�"o����������hZw��tlV�D���{Ͽ�?��ͻNZR���_��!cq�5B�G�-2'�y: /��r묹���w�>C�W����LW����ˢ_	�e3\*n�����g?
im�/2A©g^����8N��iK�ծ�_��ćU�H 6d��#ݞ�T3NZ�b�C�_c$�X����toMRC�Q��{�����&h�Y~F9m�jw�]���Ͳ_�'_%bR��l:�Ӥ�M�8�.��N��ꮯ>i3up�C�����lӳ��J�}J%�9$c������?�@�Xk�㶓B3\�S<�OU���t
��������4�4l��w��I��X��Ĝ��6�-C<p<�8C��0��C�����P���y������&��#�j���jԼ�����:�QĆ�x�jn����^�]�� }�f���y�(v�N�D�K7t�~GO�����o��ԯ'�WO��e�,+}�53����nc��w�G�.Y8��yk������3���>3���Be����ظ���8A����R�?rH�za�E1����#g!�H#��q��|�D̫۠2�͵�C��oj��S�Y�,Թ��@8�nŜOS9�M!QWJ��(O��i(��7��;�_t�*1��S	�o���\j_���R�3Q`g��VT}�ў=��fޅ��Yp��:ب�7K&�B��!�h��ʯ�)[Q��C�i<��W��_)	1��ߝ�K��|܆��m���H���,��Gk�J�瞢��<Q�{	�L{M�>}VB}C38	��F��]q6'�El�En�3��?�S�a��=!�?%��_��4В�l��ض���Q y͡jK�h��n  Zcq6li۾Pk�K���^>��ᙧ��1kq�;�Z���8��aSwIc��OZ��N�ކg�W4���|������Ž�?@e�VL��'#�1����/��dU���g�)q�-jCOl�Q�nh;Uo�q�F��T"����s��n
����ٴ�晬Fj�$ݎ.P����"g7����6�+^̨2{<����s��I :��f�$A�d�*\>�/�[�T�d���4�^�'��v�����r�_�d�V�R�T!�]��{wO����4����?���-�L*$i�f��4�N�>A�j�*U#�Ȍ�D�@
2]�tv��e�\�ũ��亘P�EJQn��/ճ�K����)2���J�pA�έb��vZ�ɱO�`���fJa�=H��4�/��ָ�7V^4��P�]G�&�M�
U%����#��G����=N\#����N��*`�Č��_$��1Z�@V�R��;!���@lAQ�R�ٵ�tW����z�M�P����C��W�}�eK	�8ɫxW�@`E���2p�4��m�6T�j�f�%���X���䬲2��FɁK�/�G��̖L������?8���[ӰY���hwƺT��Rń��R�[˼z��C��?^�^�R�P��j�O�	����x���*y�,Sz�l�KW����j��"��yE��������rP�kD����Y���z���k��:/!�"�U�Ze�[�w=������:M��Lfm2���`:�3� i�q4ӎ�¹���a�>B��B��g< �(�y5��E��$M�o����/A_�����Ļ�$6��J�����z%^��v����e���\&��Jތ܃3������l�Yy?:}յ��08�w�U�݋�ɫ��f�o�o���w�5]��,�_M�D���5�:7�r�"������4��}��.);&�V���x��"����㴑�| !C�_�>�ո�����?�/��`��~��j�"���y+����9�U>�D���Oe��O�_�/�;kP�2�f��Y1j�R�4��{��*A�"6���A��NST�U�_z��o�60�^��L[7c��ϲ}D���k��s#��R�$���Yg�ꋮL��\�?�xx��᫱�V�}��I鈈������F6�7y�^�J��kM�,�t���O�l�M��~v˒�Y���m�^�a2�砰Vݩ�����V�h�X���o�+�8��@�|c�Cc�O��ý�u
�ǗI�˟V�������XlPJU%6&�NC�SԜ#L`�CM'�䫫�e�^v�o�lE�K�U����7�����������'7���\o�L\��0�xT�X��	Emk=�>o��aF� K�Wf%��0?���@I�Q�Ԏ��ui��K�'[zRV�><Y$�Y-	��y��F�~�+#���C)���z.�UO��ۢG�u�D-��C��y�N9G����'������N�&��"Y˸�
��X3N��������TP�:�E�]�4fa��w.z�'�}7�;|���(���z0j�t�'�����Q�57ۿ�1Q�(��=��ף�Ұ_j��ʿ'#A�#�E�M��(�=�	��X-d[yB��u�̀�.c�Yn�����}����G�'��*�����C)�Ib�	�~�w��,�C'��;99W�%7����� 5� ���vO�o.%�!k�gT��m�iV����-U#�g���fԟ�ݟHZ����=2#[�l��Ì�k���d�����Rw]��R�"z�{�	�ǣ���h����b�kKζt��(����2���p�F^�H�v��=iA[5c�y1�Z\W���J}�ii4$(bSBGU��!MN�`�;�ݘ�(�8�ߤ��Y�G<��T�V��^�(��v��7k�\�s(m�H��횉���}.3�DV��M&'\G��DAA�J�a����#�ߝj��������(����6+�M���Dݧ9`6�Z�G��k'@!������]��Lѕ�������Sb[j��P1zJ��p�Ry�,>;�^����u* ���ҭșJ��Vv��(B�̚�J�����^����mHq�S���I�S�\1�.<������oW�D��T�/`bN^Y_�_�����AFB�뤐�:�N�Ý��l�X*�et�&s���_����NDPDtX�Ҫrze}���V%|d�F�����F�� ���]Ґ��lLvA1��]���h�F8@�
��%g��PX�,Rps���kw��\�M*�f�na|A�9�6Q1��`��������W��H<�/G�ႃvIb��;?�}�!e�vI�B��Hu��[��Y.���r�?L[�)K �W&H�J��5������h)c���n����>�����+���=V�UQ�7x&�n���P;p����ͩD9||��%YL�a�JS�@vLq�Z��<�5nj��EXZ�?3 #�L?̛W�~S�6�Z7y/.;��n9aqe���m�� ��|nF���;q�T@.o�("� Ըy8��R�a.󖯡͍ț+u?���xG�x=�A��f��͞i��ڋ����y`���1{%��&���@־��U�;Ly��z)q(����D��Ŏ=�_=�L�<w��J�ֿ�Y�`{c�=O�T���+�4���g�;u���Z����ʢ3��o%�z���\�ҿ�*5![�t�a�Gx'j��E��C>^E�M:S��/��5+�b�c��>�th.J�?Z8����tǺrUlK��}�U��/Ϧ�҈�\r���(�Y���m�罇_��*�Бsv^B%��~���E��J!p�D��y7H䓝����Rv�B=+!5e��E�~I���=�.w��Pw��RoV���w�XσxYPw0�n��Ҁ�\�=�ǐmێ�]ꐤX@P�͟��1dx�1�;�o���>(^��ޤZM���l��K�?H��L��Ծk�^x������	�����֟�^�	џR
���ҧ]XwO(L�oK=���f@2�|n��8Tx���h���@y*3Ko�����<|5*���qK���!��xpVH������M]3�sB͖:~��4C��.�M<�0�����m�J}-���� ϲ��Ƕ��]V�-&lΚ���J}��jr�6:�Pd#<[,��Nw�$,�ٮt4�������"�'o�?���5N7���_���F�V���ddf�$���#���"XWި��KQM����>ħ�X��<g���å�zo95��䎢�k�����
'L�J�6Տ4#
�ܷ%L�	���aU����}]��"Qe�\���x�$�>����,$A�?�0,B6g���+�v���q6�rVPCK��4OK5̺ە���o�FH�n'���
Ri�.f*��E2�i�߱t�p��}w̳�ޡ��Tǿ�d\��,�s0{��*���Av�w�Sx�=��ڻ�	S�����e}��U5Az��%Cg9�|T+��'�6�!�6�"��n���8�h��sR�G�ɫ=�αa)eԛ/�4�|��!?�m���S��~�J�Z_
���T;�
���Z\�Ѣ]�&ס3	�k�4KS:6��ZZ��n��� w���*�M��E��i�W�_�i��p�+f�eG�x�:�7~��Ս�L��F�_���;�`zE� v-�H�O����Z%6A
�e�N>��x�XPdU�D�W$۞�t$��ţ]B��ol�D��M�!}�R�WD����!�1�>�	@���W�����	��pY�u+�>!@��;�YH���d�s��"�C���c:�	 �Z(��I`~�o�L��p�Y�t���y���<auƚ�LkQ'�$���K�H���q�̝��NNEq��i�7�s�7�y�
罴/[�.<5�~����p{(�ْ3�AEQXm+��h�0t��p�%��&���g�Ɯ�n��z:����A�n��,���ND���s�U1��2%�ë�"��ʱ�縴��xw|���@�#e6�c��Ξ=ݻ�3�ځ�/\[?֧��|�kL�ZZ�t�8�>Z�
mu�?�ǌ����s
�1�ɰk�<$�$��L*o�@㻫J~B8�ε	?�/G��ȟ|`���3�7�9Y͹�{�{H~7�)S��E��H���4��HB�-����o�_4���U%*d��}B#´\��i�FQG�j;�뀹$�͛�f���ze���[���0o��Fw^�ٝ��M���)���ۉm&��2bee��%�Wu�}��O�B+1��>{�z�7#�XŻb�4���&w�B��Dy͜��(�6���ew�u^��<e)%�u"���iK�k嗩�[k�3�k�u��*�������"�W.�=��t�lL��Ƌ�(��%�BQ�'��1��l�2J���x����7�Γ�֝�fv��%��OGm�>��}��m��	OYk�}=��]	�gs�:B:���q^����x��T���:�M���Ç�[��&�����x1��y��7��K' 5�@�!�u'5��u� `S�����r�!Q4�ٮ�z���g��D�G޷],ѷ�����+�h�+W�:��ɩo������Ͻ%99XU�YҖ�x���5`�i���ϩ"���*b���Q�vǤs��t�L��@���'�w.l/�a��C�����MbX���x��g���� }kK�-H����0C��D{Վ9��������5�JtfCp~���vo��'j/K���t00�H�F�=DuR�U��\�*R��R���?��E��N��5o�[e���a�Q-�4�EW�(b�b�fՙF���8b��%��9�k8 �$�������N1���k(4bq#˪��=Z�W�m�1a�)������l�+��tUM�l.7���k/_�#⟽F���'�[�K�6�2"M��P�;۳n���8�~�bM �j�8���)���T�
��w���a��A.���b���������?�vw�{I��g�|��k%-8/#�ni���s�uH�ҁ��XX���Ե_���>2w�A��n2�>p�D��ǜy"A~�vX���w��Ч�d=���m{��w��C;A䵕�߂ǯ�����wx��GA�Q���g�u����s�@F�qy��!����.	���_+�|�	ը�������:
k!���
Lf�Ḝ�޷����`�ə*�ϡu!���@�`�P��ᆻ�p��B���u��"]��\A��0���盉��o���?�|Q{d45e�ǅ�_޿U�*^ӽ�р�W]kc@��pCg:f0W����#�NH��A�\�G����>�h��y��L�� ��<m̌���4�eM��sC�m�%���y,�M�OU	x�M���]��G�ez�`��8W��%��3�G��e�^�+sN&qR�7[�P0?,�.T|�����m��G�mr��v���q�m3�j�~�-��ѿ��P�y#�W�=*��[6�g�}��i`��L�E�kYV����X������<�[bd�.�-�ۼ3ѷӒ���8�������ԊlZp
�$1c�_���4!���Й�6�S߼�j�sR���A�BnA���l�W�dS����`Q$7�"���l�e�qy"�,��C�-���zs��x~���B}z�I��"j�'k[}�.Pp{Mx��I�s�ʫw�'߬v'�\����a"�2,�-:<���=-'��T@=h��%��8�s��l����ŋ�=A�Uv�}u����ەx��:���3����	/�D?[3��&1��Zt��Q�;4��F�i�E���.
v�' ��pR�k�9)/���5�c�,�t�i��∟E
�5�*xZ�f��Ԩ$��E=���$�Gع{ǿ�
�cB�U��u�� ���� ��B�ZC"��%����m���K���<�� ғ���ٝ
6f���W ���ܢ�W��^���>�َe�>�PK_Q��Z^
 4���ʭ7��p����'�j�m�CVb�N(ʼ�Թ��<�c���3,��g�Q{%�T�Ϫ�z٨���Q���h�{�=���[�И�b}�����U�#7^���ѐ��R�����ZCWsXA"ٓ���6������Q2�rO9v��e��l$����Ǚ�ɰYe���{luο��2WP�o]��F��<,�+�mĕ�s^_�Đ_b-(�m�a�����`9��z�-kM���Q��C;�{
{�	v+��VF��VS*'����(L)�60~���q�Ex�B���L+��OXΈ�y�?�+�F��_��
�������,`��y �a���(���Ulj�I��a*u4��eV���-�$t�y��ej|�f��L�n�2�eG?��K�pt+/�'�f&���/i�`
�Ȧ�V�0xr�휭��J��Ð���wFQ/�[��#ɣ�9߈���,�)(��yqE���I���t	���9�[�IVJ�Y[U������*�x���7�fϕ����描���_o��o{)5��h8wԓ�I���*��WF���)ߊ\��٪}�
6t���?�?�?��g�_V�lz��ݲ��--./:�ܯ�\����"�A�c��`-��ֻ��#��k��N�V=0>�6��2d�<w�CH-���b�"-EU�N�*�*n����U�67lSSV����/*~EKYL���e��u�͡�,�Q�|���~����/1�C};��,����M��v�����$���=�������aV����T��BV��S+G�HG�b�z��� TJ���?���[�X�3����76��l������~����o�]�'HC[�G�C���7l���^b�g\Ժ�c���k\7��� �&�á���01�~x��#uхȈ��H��!���t�q�h=����DJ�0����!�� t�p]�E lͿ���l����=�պ��"���@���i��/�H�[ޛ�xa�B�?�F�&U���s�9�a����ƲW9�`݇*9�*�IBʹ�W��O˙ͻ������ވ��t��5��Rq/m^";-]m�|���Xe1>Z}Tp2	�h�;�O+g9r̼1��Z���j�ZfK�� ��t�X��`&ܘ����a�d��?�)&L93)�h���̬�&�X5����#�Dq{'7�Wg��S��6H�ǰ*
;��/��!����[E'ܵ�*�|{0����p�ӥ��a�>�x�{��9�P�0��,L�uA"�|���T��t�=�V_5���� o�({!E9��~sj>jYԚ6�h�J�W�g���D9�"ߵ�������ڙ,�*ǶM��	�g8bܱujL�*9�P�� .�9�fs���R��.d���N�fi��`nl��)}ǟ!Ƕ������i���g�l�!V�,���:#�P����Ȯ�ڱ���Ɣ;!_�կ�p�ɶ��k�CONw���[�.:��œ�EV��]��ب���!����l�@, B������������	s5���"�L�w`,V�i�a�gg_ˣf�RzD���$�Qh.�]�����my��q�g؅����
��H��_Ɋ)��Zvg3��	N)��ο]�=�0a�[�~K��=&\�o{PWɺګ2�d�y��;&�������c����½}��VWxG��U$ެ�)\6'�>��j�6c.���i�n*˷�Yh��J/�٦B5��Ϟ(;|�mǁw�(Q^-t��6�]MdC8��Dx8I�w�[`���?�5G�*�k�'����iq��������$v�2u��I��[�n^��^��?Z\6��v3]:�#ފ���lU7�O��9�>�a\	��3�UK� �{RӔn���������l�N>6؎����.)�R�[��5�G��ni�`��rH��z�i�\`5��g8~�E�u����y�#2�R��5��9��6���8�z�u��u�>Rz7����.hV<����W�M�%�{���B4=Aۺ��ւm�Z(��=�^�>��"D奎׎���1Ҫ�@�P�X�y�g?F�ŨRh��k%����>Sv0#�I�37=�r�������݌��2��նȼ"�4\G]Ϲ���z:C|��W�Vc��U,O������%��N�j"�6�((���r�7X^|������
G��O,�_�<,q3�2iC�c��߀��<���ٲ��ƽ�-Y����mC���G"3r���a��2c��#Zus�h2����|�:��L(�j�'�M��)���Τ{���a�4'�� D��C��l��.Q���a i� 3Gr_�Q����Zd���^b������9�q%ah'��ʙ�B�^.���N��Hf*ԍť���:Cz���G���>ɯB�[cQ��Py���?���P)ѓ���'u��oK:���0~���)E��
�:'�=[��hd��@u4���}������5���g�}����^�a��TA-HX�%t�ƻh���56?�-2J�J����x4���T��_�F
��4��� c�q�_��.��*d�.��b�/L��2t��u˛̱h���D�p�qd�D&ϛ��f�&}b�o�Ą��| $����
�U�K�|��d�v��ٹd������;���׆�'o�:�Q�#��4Rc2H� ��z�%�Iŷ�YY�R����G��Ã�#x�Pk���C�����0{�/>���9�������5]�$�$_W��{;~�Ggqﾸ���hI�j�hD�̿�A���E�I����(�7�L�:}|�L�e�8Ѭ�3g�UY+������-����b�uz�_sb��;����γ� �X� ;Ҳ�/�M�W�_�*\2���ކ���~:n�����]Q�HY6?���O��>�����߉�v��-�7Q�x��¨�Z��Fՠ=�@=0�V
Z'Q%s7Օ��M��y�s�iI��x֭�Ev
+�3%8��ojKٹ6�xc,��K��cä����0����_rE_J처���h����L�Ir�i��z�V��j4k}�D��I��;��wbq��>�"�Ά��٨��4l�lb��M��9\Z�ɠ�l���Fh-�o��N6� �%��O�`Do���~�<�J-\?����(����ʉ��n��$��8�\��uK$�<��!c/�X<7)�/�<"^�y5k��g9�kgph�
����Gu*�8��j�ڶ�͹Y��T�H�5^j�K���*b�w�uf{o>�;��oN�jG�G��T�C\\f0�nxn�}�Ɏw)��o	Ox��M�I��u�r��>��k��6�N݊����&8?
�*8���<�C2J`�
{铰$,����]���H�ӡ�� �2-��o�!�?���H��;�I����ͨ�̴�'�;^��k���V��+��mZ�t3���/����t�� �E�R�K3f�j���_�I����c�7��եo"&�W���dx�A����۝��?���Qjrv�|��V[y�neW$6/�ˡ$5�?q٧rK?l$�����;��g�Vu�x����nd*�Mo��&��50�V`���l�jd�pHֱ��b�l�o��]&�����Lz��EEgPf�e�#/�t4DTAB��x
B��-�o@�7`ֳ'�B�Y!��7A��R��,9r�q�H��!���\�@�|D~���9v�Y]��t�]}.d�®z)/J�7��[�?%�>R�-�x�F87�}�X�k���~�0�����\���b���:A���|��2`X�hRh�N_q�BH"R�؇�0�,<r�wIr�kB���_��0��Z�]��d�6���=���	��|��2��p��rQ�-$��HS�	��� ��o��c�1`А9Q�4YH+�)Jr�ge$t�"��q���Z�y-�HUe�'�%��O�	�À6�1�tG���'u�V����>��\����ڰ���	�+���K��B��������EY����X����ZAQ����cТ%�Y���w֡ ���W�C��7�8%y��%�V�����MU�{��N�	��������$2�7����ޯ�,~�dC�歭��\�St(�Ҽ@umn��7�'t��_���|ˋ<B]���t������D�����&YF;��%����v��t����ш!I;��WNZ�������2E��9"mTkqf��R��2�'�'�����Z߹�����tp�\>��2�=��:��Z=�/��F���u��Q�k�GOQ��0�7�X֮)���F��܆�J��B��Ν-̎�sLY��Ug�W�$����X����c��Q���>�A��a6�����
�@m\�&�P/v*f`$y��"�
����5�_�lay=x�4�����1_o�����mư��9�1 �+m� ���[{Or��t����W2vX�g�jy��%�y�:�:���'-��p?14N[���*�F_�2����o���FZBJvӶ����<�	m����,��E�k=RBi��>Ү�6u�t���Y�1��a�ş~��M3��ID}�Ŝ���I>��U���%A��?�"���+5k�W81q[�����"_����nׁR{�H㻹`:	�@�Ѭ���o���W�j|�"eI>d'c��o}b���J��֨?���y�-���@g��t�3b�	z���ԡ-�/)I��QP������]�����`6�!9�����y�W7MG��r���"lZ��R�R��l�iVwbV�;炥���P�o��U;�&{>��cTtx�8JW��F�Cp_��& ���]����Ux�������Λ�	���b
қ��@����.>�m��y��8HJ_1%��/�k6l�2m�Ѧ�R︵��a�9�|�e�2f�G6�"b��������_�9�=��[�$K�zj��^9�M�T	l߿���K��9�b"��}[����|Y���#�pA"�A��9����|��@�T}�K��#"���Z);J�?JVT7�ػڢv��Ѐ��m��q��-Π'P��}�@K�Fŷ�rt�o�ļ�	��e{6�뷮�z�zշ[�ϳ�s�8��c�w6���q�Q���$��<�G�u��c�ѫ��!�>�.����O�|Ҙ��ә��{V���S,s��::˵�g7q�)`J_��Ħ�uO}�3��iyڜŇ)zde�%5�Y�A��u��M�j]$\ñ�4�����p}�Z/���7�w�x��)r�[����t>R������w2)_����W��� n:h4~��rV��=Aq����P�sz΁�~3����o�vCXu����v؄0�fjoKl׿w[�xm�"��EVJ�o�a`�	t!΅P��D�_Ώ{�*�B�=<s8�W�����7S���]�!S.�����S��f�BO�N���I�,Yaj��0wy���)g-@H���Wb��k��p�ˠ��#|*���ׯ-A�Tq�&�>�9����11C�i�ͨ�����Ϸ�)#Z��)D���v�y ���Z���~�J��K8��R�6��� ��f���s�FW@OB��9�T|P� P�1�Y��&]���e��̡�-?��5��Y�������E�}���<̍6$-��E��C�����<m���_@��t*���vB��qH�%:$���X���%���i�Ʈ��?!��c�~r��c�W!\H�2��#�mu4d^��L�=��wjXRùrJ�b��7I80�����"�]��S0�w��@����پ��>������3�Oг��8w�'b��;�j3�:��Z�9�A��4�Nх<zˈ�x<��)���Ue���p�!�����]I�� �p���x�(��Xo^����	ɴ�?T}w\�KЮ���#�DQDAAz�QzB�R�7�$�(�4B�&��^B	$�ޤ�J萄	I���w���ewg��y���}��䢛��[t�.N�I�Wx�gP�f��n@@�"�z�Ů.�wo�0����$�u+]��򛚣�Y��8Gbz������2������u�����kG��%}��m9w蚓��OЮ�E�w�������EG�-6�a�N�%�1�\)��q&˲ɕ�K��@�����Q�h����+���XǭL�H����`��뭔������cHO����e�%5�,��-}��1�i¢s�͉�;^o��L�Ӣ��׀e���\�#H�7'�z����ނ?�,����FMak�ҺD��~4iG9"M�A0aP�A�4{��]��i�X���Tg���.?����s���
*�X\��%ԎR�$s���U-��B���Ǳ���/���"7'�z�0��+��RL>�׹�s��.�)p��x��9-�h7FȑBZ��k�[�d5�MRG\������ˁ%. /m�0�Ï-�,ΠEN�wZ�oH5<����6͓T:?�:lé�Rc ��4�����7�}=�g��SV+��K^�L�n/��ϵ��{����=+G�������WR,ys��c�TuO�E,�r-e�����������q(";R��w{*�C��׽g���+	UQ&=�eĈ��fŦ��ύ�����_�������V�l���Q�-�p�̀d�pr�4�q͚�k<�N͗�2=h�t�g�~U����-eo���y_����fJ�q��	ǗU�������EM��ɼG5��I��dc����=�R3��Z�Jc��J�����u��%M@O�8��f�U@#γ�>�c6�ok��v�k�������x#�u�Aڨ�>�W\���FR\c:p��ä�W��"�s�ӝ�Q�Qd����HL f��@aw��"�1@��Ua���ʦ��&5�|�)~����"\�7�YC!�w}x������������w��9�v����I�[5C�җ8�|�T��K\tb ��}��cqhK��-\�dbF�Z�2$�&&}�u� 6Qw����'Ԅ�_h�
X#�>�٢��]�O�"ҸLM���O�����<���g��b����_�r��TI�.Ǡw��V�/U��<\�[#��T�Z��(��e����K�������ĵ8'©�g�ա�U*\�\m$�2%��`��0\��9�}��S�!���3F>�ss���sZ�@��Y�|�X@���A�����,@��e��g�������_mt��\5���2��'�ȏRof��fq4����4�������)֯�C������殹�{<�{�<6��N����y���ہML���>˷�cQ��0W���AY��|��O���m���>�!����d�#���x��E��d��|���ާ0e@�V[:�J�Y�P\��)�tg��?�՜�r�$��}p����.�)����L�J��K�!3e�lV�.�17D���:'�LJ������A[�t�r��s�b__��G$YǷ6�R�x�pݩ�<�7��V�Ռ�$%�R.q��*��X�_鴥m�;���#�ss�X�X�W���1u�o����A��r~{f!�Y�0]�����>7�,�#��c��(�o6�J�C�Zh�]��Ɍ~ڽ�~{ y�tR2{a�U��]{$�����[�I����Ľ�2.���:|���<�)7cb덀��ID��o���7߄W=*�B��6����6�jk����@�P�s?b��/��"�]e8���V�@��.�fb���W~%��3K�=��ɥ�I<���'w���l����O9īӆ�D�/��8�A+?��ҽ��h������3�'��-�|Q���q$��CEI�݅���l��&���f�@�O�9�}��_1�\c>_w=p��2�����4a����Uh���ެ�ƁNG Y�k]�^��rm��SA�_5�Q�actfdK53����A@t�6��</PC)�v4�,\`,=P�����hF�(R�3R���,�.|��X�<׽K:(4���)�K,H	��h�w�FB�V=����(��wVW�E��Ǣ ���U�X��L�����U5n�A�}D���俫h �����%���f��4�ݞ�o�M�l�*i�4c���5f ���aYK�iD���`���g�����*3y����KJ ���E�j��crײ��8��� tWA��*��;T�R9�yO�o��[�g��;�n������7T�b(o�{�p�,��n{׍����o	�R2���M�=���2���e M����2��y��Ƞ�7h7ˊMr�JҢwWO��j�vd���>� ]�L�i�N�|�]XYZ����8�J�)	7}�$a۞������\��p5����A��`��ӂ�\��^[ANv��	��0 � ��HM����?�`xz˞�_DB�H��u�
�{�'��+z+�c׵�H�O�4�2�;R{8.�5���~���}oy��kt}���$���uh�:i+��V�(�vxUQ��
���]Pbؿ
����H.M�5���D��4u���̴?u"-�M�C�1��7��OB�\B�a�21,�T��sb���U�y��d�7aҿB���ּ'.;�a����|��%&���\8YqD�/e���Kjl}�@~��^��>�h�p��D]n�;����#NdC�'9ޘ�l�w��J�.K/Z�1W����?����7�%R��Vۙ}]�����fs�sx�lLۣX�X�/-ߩ���֍J�-H��_��` <>D!2�3�v7�M����'�$v^Dn�g��iuA�h�e��8��Q��.8�u��`�~fo�ܿޅ�N�v��VN�;-�&�>pG��|�n�S�ʣ��8��#�遗��������f�֣s��яR��y�X�#-� �"a��@?��I>�?�_�XG��L�5��++/����y�n�����������ݷ��l��`�7����t?�l����J<���*���S:�.˫�=8���TԠ�}g�5��}�E���	^/BUT�N{�3rF�q�j��g����/��K]����Q]K��������歩Ƌ?y�b����ɥi��{VG�#�������P���;x�\��#`q���Ѻ�XLĹ����Ļ)�ӟ�;������}.�����~ ��G�-���$���芳�~�~�PD����2�ݩ/y	��9�Mh\_n���B:�T�f�8�P�]]�Ѭ��j����耕�i�.��7Ic��V����L�4�+}����Z����fR�L�z�Tۚ�q-�S��2w�"=j�`�y���zm`�aZ�ИF{(��`T��W�%�RK.I���9��]��Vóu{2��m>�n��\-ĥ13�R*ҿ�[�
��xY��O���ޭ�Em��If���	���*�i���y�� r��^�[`8�ʣf"�Z�~�}�[�"������w�����{��\x��ܖی����oFSK�����%q dQDAIH4����6�Ney��ӣnQ,"�l�罻z�Zfv�nMh1Y�Y�����E��/5p��>�+-<M BHk�_:�Qf�:��N����c�����7�7e�Fq���-Nƒ���w\��� �.�.�{D�, ���$�����˒�S=U~�#k�T\p+�M�["]��
�����+{��/��e)��R��\8]��J��C�QL�=l���U���#`x5�4�-���ҭ�fs~K�k��7h{�,f��bǡ��W�><ё���n��9,*W�)�7�`�W��X72�p��4�=�.-@`�I�&�J4�l��	9��k(\\5Il�^3�B�[)Z=襗.�����i	+��-�uJ����w%~(08�yq)���Ki����ѿ� �ɉ�����"g6�m,ID2>���7�|�6RYk"8%�Ĩ��X�y��n�oR��}�!����im����ǌ,��:�t��ٜ��3�W�ݒ;����S��s�4J�ٛ�L- ���]�v>��P��H��t*�.z+h�M�NG�Ub; �(Ƌ�xR��vl��rdZ�7RH��/ۏ%N~��($6wjT��@o���	��>�!�1���h!�Y��������A�:o��g���["�/�Kg�nM%v���fڵ�������׭	^�,+-:~�����{�ۃ�݌��	�i߇n0�7�8IN�G��OHG�z�4�aW�����1��i�;�y� �e�s��ۍ5��䠧z������`d���Ë`۵��_���s\얒J�V��2��U�J=0��OT;���ħa�~�Hx�_����7NA-������xN5zQ��+B�Y��OT��t�✵`̈���ߐuuVU��j�1�g�(>n�~�MP�n���]�K�L��aVz��]��%�/�q�޻'�G��5�� �e�6��rc�7��0X�Fmhl�%���I���������b���~������ɑ�9�U��^�v��q�N�O��*���(�]c�l����w��̬��6�,��T��lN��J�LM.���M3�ʕz��a\\]��Ъ?,#��[s<~D/����O��$�P`��6���I��`�?o�N�\��^���5�%m��[���bC�� 	��˫��w�:d�?��k�v�lv������@���J�R�lG_dQɑ����i�,F��%�2Bʏ�K���z������fd?@�'F�v��wB��-Y��q�SeK-E�r.KET��}H+3���'~_�X����!�~�i���yq��.�����I�F�G�V��狟{:ГU\��&�ν
#դ8�*�{��t���L&=�&	y��z<���e#�;���諾�o��8)���Xu�����$�m"t���A�Z�&�-/r5񥩽��S���"�5��tACG��Y������R�.��Bz��/�":μDPp�qH��c��1H��tؕ',��(M��l���}��rv������
�Ss�����^�O�u~�i��	u	���eD�i����r��wL䱰K��+^>s���������m����*�)�|��9��n&{zv���(���;���2���OF�@/��i|>��NP��-��4���C�ov�+&|
������u��ɲa��v���je0�F0������c6�{����5rr�Zv�z���[�.A+�ή��U�o�k������|�i$ {��!��Wջ"�	��b��M1��xl������떙!
�wõ�Kq(�؊>�S���e�A��K{sb]�d�����Wu�j�����B��#5 ���hr���9���v������x:%���{�>��i��Ƅ΄���h!�u��+�5�n�ć�b�;3"(�"z�k�[��6.l�Y�N�ąF67j���֤b�t:�6m;
qܦ����wY�v<.�#j*=�v>a*娣������+z����|��I�����uӏ�sEpћ�xl��وhȫ��CpP���K��fe�ɔ�k{�
�`b~��ܔ���V$��LfU.��*���bs���47�~cH�?�M�$(�-9��"t��W�Q!�ﴍ�-�����#�%,��\��������QTԴ0
	�f8Ua����8�:��R1[���o�&�gk� ��0bN��d�)�:�YvCsCJ�X�ٶ܆��	��.�����7t��A@,��k��d�.�I�&�t����e��/���$K�a0x���J�� �X8�Z�L�}��X�i$&MVb���Yg]�@��|V�TR^�k�[��j�Y��p��z�g�H�*	���_�h���RF�MvVm���%�~R0e7�0B�S�>^��3撧�Fx��i̛v���frw��Cl�&�y�{��N-�'��Ey<�X�G���%��㰺{R���f�`$�v���F�2#6e�|�6< C}�(ױDx����\�)�#�9Z*�E:d��>�o�:�B���P%2�3�%~�}u�o�K�N����3���iV`��U���	7�-��L�t5����04��w١pU����M8�-v�7���?��H��ڷ������D2�3�ҭ	��Z6>�ݼ�"\�N����=�/\�"���Y��@~��������lgsw��&h�7~�(�;���kp�{h�O��Ӎ�RDT����&�i���k1`ʷ����A��(�NNs��/�ٰ��N���e��#0ZS#[׀�6����Zh��my���7\�(��(�M�i�QP[Oq�2��GPs0�-rY(�C�o �5jd43Q��oǌ��";�%G��"��<�L���o��q�pŋ�w������̈'�����u#��iY��G�}�S��91㋱c)G�{qP~�%��T)E�e0�%���y�4pʢk�d��F�.��ڽ����&Y&%��B�2/,���N&çj��a2��h�c�P�ڙ\�a�E�}�X�<^��ۛ�L�a�b_ �8��b�;{�G/��/�i
��%���oE�.k�R�uiTNo9D�\�s2i|�B\kD��v�Df"K�~u��CĊ���Ы��*b=��v�iB�:���iv��kT�쬑��[�6"����Й����%�zٰřn�@��?M<�_��#9%~�*N��}���Bxzit�I��z+kM��h�7l��8���r�\�ȳo>$�J��L|�k9�(�A|[��>�f����VT�#�[��i#�/d�!F�2�b�|s:���מ�[5�Q���x���pt�1�ko�5�����K�O;睜8�5�
^�������U6>{����Q���0���,-��	R�5.�Kw���5��\�뫧'�u8��qq���vJ(_��xK��=�����G�q�t�����<6m"�%� ߟ��ǺT�2��9����w�;q�?�b�2`�!��{��8j���Gp��XsD�7�Guu�}�}7��A�y޲���ZA
2P�6p��1�X�)Z�-�~�޺���0�#H00���YI�V<�*�L75�\�����*W��"L��������v#��c�����@)x����䒟;(d�ڄ���K���S�[�mX7S�W�W��Z�s\Z}G�w������R�\ ԭ'>&ܘ�G�ď��'t䑳+7�Ւ��I�A�2 =g�z�꩚D���{۾~M�h�G�{���+�����Z\61��V�}?!G#��b��oh�gx�����a����UL�yE�R�{��9�\L���%`XW'����lR׎@��E���EQ����sPǌ�MQ�XGb��������L������'��+�4�6��r����uV:V�{;�s�6�в�	���fJe��1�޾�9?l�o�w�\d����e� �ʌI��u5io��8~���~^o���m�� �80�[�S�66�d�{�Q�bV�ublO�z��S`3�6�2gxS�6��0xP�u��V~����(/8'M	2�N2���?��^��g��]t�
� -��9�L�N�6�9��Pw�Y�+�!��~*�3Z�p:���Y��^��Y:��;:�ƴZo^�[)�`0�.�Y�����:(�>���I�������<g����]r�7ݴfF �FZlb
�μm�J��h�5�wt{�V�BQ��ݍ4�v����e����h��>{�q��>���DTPC^��U����n-�ɻ����4\�<gN��u�	ܩ�f�:q� ��c)��7��1/�r�����e�v�h�"W�+}�~�fh��1�Q��b�gt�r�m40'���9���Pw���O"�O��Z���"$���o�$tq掆�j<a���6����ۖ��_�eX�U�J�����p�����3泇Wl�����eڦ1����Y٨����x�M��\�a:��ƨ�:ܐ��;Ca:'�.���l)J�j?rI1.q�F��6�"=z��@�ٯ��	�hٖ16EZ�St��M�_ e�6�'b�4p�-%�,aR/�{�J>R�߲�5"�7\���I��̬w'>��nEJ�c#��8x�(S֊8�c�0B5=\NLl'9N�ת���
	� �\��z��g�ʚ6��.�I�����E �ӟ}����f�w����93������i�W)Z�m���x/�~����Kfʡ�kH�e�|�sjhh������;���h���լŮ	٣�.除�Ĳ����Jg�SRgz+SsR"����\�D��KK���|̄�C��2�ɚ6��3~�տ�t�L7M��_hh�4��֮�Ha&��x]�CQ�#�ޏ,k6S@�����Q�0�S8#�c�*��������vz�g�Gu�D���A�l�|}D���%'ˣ�#6U�����R�	���Q�.��&wܰ��2q|��kb��k�I#��-�;%�](~B.�c���.�����*�<e�����@��d�lxS8R�<9s7�nvp��]�H|B�r�vz�j�� ߟ�����kc_8*�s�$��3�1�E�.�=�ߖ&̵;#���p���0C��gD�����~��dޮH%�#V��)���y+4q�&�r��B�N�y��j���v�*�>�{�s�l��uԮ1���ߟu���I�
�� 9�ۋߚ4�ۣ�:�7�o�?���� ��� ���*�.�%Zɛ����2��V~7]3����>5����a�^�Y_��j���������������{�QOm���3Q���̫���''`^--�1C����C��|;�1A5mgO�(M�7�E-��JF|Я�̳Z���l6�d�	&m�[��we잓A�*�뫋�~'cI���f��Q�p�CɄ+ �Y�S��~��>��ׅ5ؽ��K�X�u��ΧR���"���#C���]�m�����)�%$����
�P)�?YY��	����b�"�m�_�G�GǏ{�s_g��j�{�G����s�2Y��78A0L�Q�5���� ���K-0�M�~*(���&��m)>��߲ �" ��R�%���-�k�`�p{�?/X��)$������T���5�c~�@�8��#R������V���Z���*n�����kÞ��������o+ܞ��	�?���f��hO ���������J��[��ϑ���R��M^
��
�Cu�Cd^���/&Īf1�K�[�y�� 6L_�Q�����R��
��1����VwS+��<1LFV�{8�}<F�����+���j����k�ܪ��M_D3�a���r���
NL-��U�,�؟ܗMa{���fS�5W�uƝ�U���(�<�h�LCd��xˎ�_5��`���D����̍��>p�h�� ��RI@�I�InD|�,?M���)F�wz��GT5�>�{��{��6�[pd�G_�R�G��̊��֟��/2)��6���D���K�M��w�����O�C��T�j��yc��s�diX� ����SYT_�&���X8v#>�6r�*�#oee���q%��f|i:j��$�⭪K_F�$� ���h��n��S����҅�^��ݍ=ٱ́E�A��q����z��Fy��d�UE!n0)*�L�I��D�*	��ŮaU�z�*#��}�zu	5��NG�yJ�(J�D4��S��E�?|��f[�{r�E6�����y�?<�!#P׼�
��=��>��`d/�	~w����VZy� $�2���c �Kӿ\���HH��ϨT���\���B�ڲ��<SƷ�%Ζ
	&/�_م�����KΈ�=���D�ǖ�xo;{ڈ����M��T	�"�7'�?�wz<��"Ɍ��X'6����G�|d��;}�q-Ɯ�a�w��k5y�6ܲ��A���Ûi�	1�)��5��)�IÔ�J��I�N�s=#x*�،���ɝ>�׌}j։��һ듦U�{[#Ԯ�D�)�I;O��R0�o��P(�8��+QH�ڦ*+1���a�޲���6WD�nWO���C�>Qf
�ߓ�3��������/
4'򹀌�Ҫ�h��?$�!�N�꺏.��KxC�n��W�M�R6��D�y>�|��Fj�R+��Sz�4��AH~���B����-t�<�=ۑ�1{��/�C̔t�(�F�ɿ��|{9Nz$����1OtoG�2n8�/���ڞ_�r �y1�|�:�UK�ZXW���Zo�N0c��l�əVg����|�����L8����L�#�k����S����W�G=��r�eJK_&�H�W��B3�F�;1>��o6��śڤ����Ό����'�����������7]�9.=&�r�K0���Q�B'��k��f/��Ӟ�)[*��p�8;S�Գ#�o�p/�x)����C�# :��5��}��|g���)�3m�A��5akp`"`*���i�T���a� �Oh�����n�$�+Ԅ�B�ix;��8���O����'��{،X��D�o���s�n'F�B���Kv�k뢟/��V�E78}�&s􋋓ʓ>H-*P�p�.�锄H��6���E�&�ۦ���AN1���>���Sc���dK�e���x������]�NG� ��^{l�N�!�v5%>�#�>ɍ���S"G0ۈ�^.υ�U�,ߐ��Ti��30Q�E� ��ef.&R�, ��u�ug@]gFN����5������*"�:�^z|5�D�DԿ��S
��|�R�F��{�dV��d����S�ƪ���5a.S�R��=�����d.�5|x�jݳ�=.qݗT����H���a��\#B�E��Z'��q�nM�
�2{�����ƪH������0�=�F���d� ��DD��؝>!;0�1eդ�+b������E^���ˠ���q篴vڤ�$�>������ǟ*ī����`aM�����c7�2������E̒�����x��햰E�X��z7������0;CY�_���rر}~�"]�-3�_����\�,\��~~���גv���Ǒa-#��H��B�a�~����h�m$��3�å��&̷VvhݶZ�,�FnO5�=݁�W���6фP;	�u�O�S!�#��ƎӼ�~��hHٽ8���F��I�����~d���'j�0�$�13�V0Գh�ա�@\ATDMT��ad��uflgn�#��l
ﰹ�,��w�C|��<��N�_����s�0����k.�;F��EOo�$T0��*�=K�����Rm�-�;a���x�F�9��3MΣi#8���\3I&��-�J� �դ��)\'���!7�"��j�k�����yR]d�JI���tf^p1
xw���\�LzhK�צ�=�w��éտ�٬X��	���,���c�J��*��jr����������#�^l�M����ɋ�%b8�-����Y���U�xVo�ho1�����*��HZ�s�F悼��$k�O~���|hg:
�y3�^��:���ώ���K\���g찡f����W��-VT6�\pޝ��gl���{�:F� >^K��o����wV=����E<jy+{2��EMK�ˬ��	�o$9�bF�,�F�>I�oe�,k�Jo���]-����&��+vu9�����6DP7�n]4u����&��*�o���:�5���_�LRpNY7~�ua�W�I��3�O�r���H�ٌ���Lp���?�ƺ�_�����
աBT��\��*dE�"��7@@B�ű�C���Z����7�L����P�,��L��G���M2 ���������[� �n��0����V7a�)$��Z:Uy�>���)��`L�� ����~_wx��R���D M���v�
���s��3O�ht�l�����v���g�3�g�9��e!��g�{y��t�n���Y[�9ҹ���Ժ�% ��>��ybް�w^�9s�X=?����@�~Y�ߟƾh�='D���H��EK\Ƽ��|51ܾ]�L`J���c�S�`�ֈ8�m�(�ac)*V`]^����+��౽.;nV�OcX����Iqx��N	��'��v����A���Ԡ?�~��دsK�u��-hK�k��iR^��5�(k}T4C1,��>0YuV�]����v#E���{��DV�ؿ�IwVf߽�ͅ/R\���ʲ���7�p�d�K1�Y�����#"��%�L���J�柣�#.�~��2�dCl��Q��KD�/�!\�ê;>��f�H��h��P�g�!y�a���]�W�|�!m�](M	����Ϣ�g��1׉�K�&��!��<#��.��&q��݈oB��5o!�x@���v�EU+�;�<X�c�����N��{cj����A�� ��nD`��C������X����<��n鋷�56��4@�ƨR0���;k3?��B1W��M���x�;�q�ݒ�X�A����\��'�R:օ��䆽
��̏�|?��WUK2��]Hl��wN<���<"���eK��K=˝��5mf_"�\����k9�9��}Gq�>�~�:�5�%0��iBjvt�����R�eդ�9�����f|{������lt^�~�_�q��T%��۷/ˎ��۬��{虰���:�B{c��m�SI��
��t�3oA6������-�ϸ��ֻ�=E��G�W�c�︹=W=��Q�>�<��T�����}�-���,���>a���W�����B�*�!I?�s�hU���a^�����+�VyM9��yof��d���^�� �+�����:�]�͏�eGs&����E���np/���.�����:��q�Oc;->5H2e)��N�5�*¸���/S��c#� 4 c�J#lo���A��A�_������������B�ʱ4C����L۝p���:�Ru�&��P����&�@�����Mo��^o�}&�ZhE��^O�R��K�$>�zeHi��ack�07$�̐F�ᕜ**kx�.�/ 1�?� ��=����^��ɡ?�7)���mݵ�C�kџ%|㒯��}���^�`(�z���aU0�̆��:�{���<�c�`��h̡KoOF*ݒ�1�6ڲsh����GM����]UQ����M���j��C?��'A��L�.�m_�$��:��o�$�Mb����ϵ,9���c�]wYX���x���[sU�up]�5J�.��ڲ�G�ᅾ�BGׅ�:N�\��5�������$���'��//d3�td��r����"�Z��Z���[���m3�r���,Qh0��y�ЅӼ:�(ٰwwD���R(���+�_h�C�.��?t��������������-˵��X51�ޤXu{f�>w�q�iC���w��5��U#!w�QW�0M	F�!p��>z�'ة��XmdJnfV�lnB7'���,��Ϗ�f1��hT)`� }-��Y�ٝ�S�jOz�BH܆����m���o��Z?,K�[K��\�Xl��D�S^��6q�U�r�=��7�-����nR��ZS�Ꝋ��1�R����,j�i�x�S:
��%��d��.�zr�S��B��F�1�7���[Gl��8GXk�L��;���/g\y��^%�"+=��A�NF!R9:���|��=���k�X���#�gϑ��=^�	;(P��!zs�8�ߕ���NY�mY��L����z%��d?4�ƻ9���a%N	�/�`(�[����&��V�)άɩ������ŝA��`2Hi�Z�����Q��:ѩ�v�?�x���H�ϡϽ6���*���D'I����v�$]Q�����s��	�]�~mH�D;�78P�F���|�w�6+^Xo�	��5�*^T4�wz�\�p���/��",�@��c��b9,#Ez�lj{N��3�_�!��y���Z��^T魌�0� ��I�U~�ʱT�qcVk���͞� ��z���H8����_g�{#��ٴ^�oQ3e�*�maI�%0J������9�v�����)��ו���̎�Bp����c��; �`��'��M}�y����O���{�
Ń�'�����Gv<W�d��S=7��	6�H��K�/��@w_��L��c��u������[O�X�c�~aC7VC��
'��̥�^������[7�Q�(5ƻ�s��/廱R�����N�{��3���׎��$��B�N�]���F�z����KuI�Vtt)�\I&���6�0x���i,=���GV	�y��ߎFho�Y��(6�N6^�/�{��d�چ1�0����&:�߶XWc��7�{G���%��ko��p9T��O���X{���~�M<e��(u�ȕ\����%:{K��:$� Z���}��/s�{?�ɗ���(�y���� ��wk�gg��ox����N�g�Wӿh���rWjc�k)�<�id>ѩg���^����)W��m���/�B�i^Dۢ�Q�n;g�?�?v�gK�jBwj�3j9w@14p��:�pf5�Xx�]��S ���N�h�9���4\��V���@n0|4�n��up	Xi�Y�o�(Q�Kؐ�5��y�5�*S��)��	��=b�)q��B��� �����F)����M�1��-$��z5vd�\���d,�Wl~�'�7��� �:s�%B����?U�YǸ*#�I�f^�{)�/B0��K}�v9_V���sn<'8�l��%����|{3Pkސp�N������������r��::6L�O
_��?�C5<Rح�X�Ȝi�0 j�G����Ĭ���l�9�VL	�t�Ww��n�����	��5����'�F- �!u�;
��?ah͔��P����CQ,�ؙ׳�;�ѻ*�S��0>��]��ՠ{�T�+�;�}�Un,�LM��2'�K�����
(��L����]B%���Q��E��ٟ/��e+�\� �k=�iE�^��R)�qT�v�1X����8�����.����q�厯�ܝ��1���`�t���h�Adxs��rl�'���׬�Oo�#���]�fQO�u	�]�b,��꒶b�Me�~*��?O�ܜ�s �T�>��]���
��_U��3�Y���|�k���#�/z7�9� E�����R �Q_���@/�fE�"~n��0sR��^zQ��z������4�YR��Hиj����Z�W�����4��V��{)%ѝ�O0/�3y�A9�Jxy�n�״%����J���AS^v�P���w��j6�U�N6����*��/շ��c��_��'dK���퐫2�&�8�y��I�����?���-���mg�U������ң��p�ȝ�)�1N�Gּ�+�j�;��&^�wW/�G�e���o�|��4@�F��[,.��𗸤Oz�/�Os�C�Y����Z��r9j,dY�p8�'�k��;���H��H����$��^�ţ�S��l�:� {'v��<���jK�[1���2/h�}uͷ-��'�/G�oK�Ĥ�-���͒����U#�'�yyG�'�Z����^�q����M�N;G_����\��jCl�K�|�Ri�
�����y|.c�'��8�M{h _^�TZ�݆F���N��<�l��	W��r��	���vk[�u�O��&x��I&���uZ������<�r�H�D�e��qGq��c��J����w��{�b��i�&᫪�E6�Z�����u�K�fa���m��bæ�ł�1���u������Og�2"�~Sa�n�>�#�K�d�QL�@�;j`��[���T�x���<�nӯ���«��}��5�h����+�����l�Vn�0�5m�G�jw+�D��E7�/h�/Q�ʹ������#&g�(����釒�5��H��`2�C�z�_�;�AC�\��9ѬY���Ѡ�y%ɥu�3�7l��냯�������e1�X���`"D����4���1!���S�'/�'z��7Mj��5s�+�z> �y�{��ݹ�;�BB��*�Ȁ�vXΪX�#?3�A���Q�݊w�:~j:Z��;IW��ƫ��{��/�7n���ּMr�#ĂezK�bٱ��\�x��L�A�=�/��©-�H��y�_V�/��kyb�F��2��rj8�5�ve{l8���PK�)�cެ����r��(~�r����b?w+p�S�~�)����Z��O���y���v��7��Iҿu�O��aH��G-�t�#��U�鱈+{���rO�/��;6���5b]Yw����M��<�Q5����p�~��J�$wa��ãD�{��SPg��F�|k�;)����w�V���o�5���8���*ì������ve��3#xw�~I��1U������~��\���dG�}d���?*�<Y���P�W\@,�a�?_J�B*1�lem�%jt��.�3��%��G_�j�����lD��>N8���t�2�W>�_~��w����g9+jtT����{s���;,�u�&�|YJ�����C�k����F>�Tj��|��̍�s(�t����L��i��V�z��=�l��a�=�N���]�Z�"���R�I��k@�=!@�
�H  ��I��^��=�&��������*�f�3s��sϜ�$���ʑ�&N��,��|w.�Z�j����7�w�Y��l�-S��"K<�z�k��ȀPu�*�^?T��h�C�..�&�,�\��sFi�;d���k����a���N�K��"���R	�b������Dު�x]���Մ�_df��s�c�E��cI�{P��i�ּ�~�b�a��^W9X��=L���:d��0�}1�G��+��ۏ��`^�p)����0��9�G�%�'�y�V߅�\U�Ff-��(��/�h���f�5��F/k{k�%w���#�օmV����.��L� �{"|6Ϩ�s��އ�c�ˑu�p�vи�Zxrw�����sj?�6�ƴXy�(j�[�=
-P��z��"�����{N�����߮(��糇�MZR�%k���j�*|^��^�C?Owa�͂���ä����.\2�+[��+(���)V�֨a��HK�5�,��_���զ�h�����jpHl�+U�A"�=7�ۻl��y�_�N�gb?W���&BCW�^�[�0��.������`�K����n�B�q�Q���2��ޫ�_�䥱��
}���>=a�sk(���͂�Y-�i��Q���cSJ�M�Z��DXg�o0�TmN.�:��;qq�3�yi�r�>`W��|s��H���:@�����9�b�]�r��V�ua�E]�'�`��V��t51e+D�{���8�
����I��Ӳk�I��Q�A�zt�s��(愺Ԭ	�@.�nC���p����i���$K�l/��h7Ot���^`�@�^�|/�m+�٥�U�I���C�p��a"j�Յ��ϲ�H����������Qv����u�-�eC?�Rd��tl�ĥ8o7�@Mqeg (ҍ��%��4�������*3��ʮ].?�0��K+'��E�L��?�/�F
w&�Ot�]MX�(}ӻJ$��\��P�:��]d��ڊ�4��p�9T�>�@#�ܸa���!��}h=�Oջ.t)[��9���ձD������[)�P�P4���2B�g�Pg i��v�Ԯ����c���rʶ͓uֆ8q`��Q��uѥ֥^O��iٮ���;�'f�fuU##��s�.���4�S jS��Ō�3x�D��X���4D�.�W����x ��V�{C��*��m`����ԅ8�c, ��y3�u3�LS���&�*��I8V�%6cS%p������ч�BaNl"\��)p��4.L�٬��@��ʗ��O�zor҂��C�~��f#��_��p�j��^�jGQ�-Rh���C�R������U�댑/�J�mC���K�iI�Y���֥`�|���s��V�6C]@\=��T��F�$a�5�A�=FU�-I^����n�υ/'����Jq�9k�4B�^KƵ�a_��Ԉ����dI.�؅ �)���>m�����o_�7\y��F�� �i�_���^��e/V=����a�Ƽ��Гp!�WL
|��l�����p;�0�UՏ/m���bR:͟�ؠ����!ySהnǝ�������o�՝���Y6����7� AR��ʞ)ss���O��d#�˥N\����n�)����|K��
\cW(6�3tx��׈���͹��l|��;�Y����!:$�7#u��gM҇��;��*�ps�D���D:Z~T{���C��$��CW�羪����|H���3������Y��<�X����Ԕ��Uj:��G��{�х�����ø�
��K
���V[hE�b��
�!pE� �}(x��黜��e�D�����Я�&�\��W��)��"J^������d���}��dEY�v��rR�i�4xˏ#ib�<Q�F��0���0!��l	ռ�:�n�C����d�s�&��)R�K�1CE�=�[D�280i�kŦJiv-#����o��i���C���?�w$,{j'�e�M��>���[��������,�W��3X���ğ�e.H�޽��F�ɹn�*��Ș4/1)���8���ܤ�׿hFG�:Gu�W�b�n�ý��[5���
	�F5:S-��-�Mή5s�D�x��8�"�Szkm��..�R�O�P�Ip`����wkƭ�0��y��y�C�Fэ�#��3�MkҿЈ1�X����W6T}R��#5����t17x�@���L�+%x+V�vp��d]~��u�M�U%�]�T�y4ݏ
�a����.� Di?(�g1����z�ق
C���Z!˯(�WK�ϊ6�J:N��'�<�:_O�5�R��^A��3���W��0��-�WIT�s}��_2(�gR�3���
��$ۚ6��K�G�&q����WG����c�=/"Jjj��$]Q<A�L!���҈�������F��?_Dq0Q��C�>���?n7�e�Iȫu�~����2����_�1M����u�
%0��@��o�f�eJgB@�IuY�"�q�����O�]�װ��ݯ1H4i��u��ZKX>EX�˦���.?֥%�%~�h������]���8ȰJ�����:�(Dp߹kE��-���>;X��?G�W���ޱ�41���M�s.��j�zz���ŨM\�� t�F��z�u"�Fyr	��$���oA�9=��b�ԓ`W��2!�eD|T��"�n� 5H�9�,Qͽ�}���>سr�1�#�R�����I�<5cE�4.���"B���.ўL�s��@X��	���̠ζ�J=�k�������axű���Ǒ�R.߰F������4!�B����|�a�N�^�M���#e�Y�	�p���^?La��������h���l�A�Hb�1<��������j0<C�ꠓ8����ˋ�߇�3w��F��~J���<\���ǁ�{�����k���M�����~;nF_{��~Xb��jV)0:���$t�h,�K�"mӱ�����J{��� �z�)	!�͏M���]�y!w#mX@CF�_�A�}���Ϸ`�����+��l��ZJ���C�z���94�~��!�W0r����#�=z��2za
�
�3��?�5$B��t��Y %!^�%o� @�E7"V��r2���r:���;�_0Л.�1���*w'=���l�� ޼�қG5/U��g�/Sjt�s��`Y���E^��/�r>;�pwmC�UH	�z�<;�� }�Z��7�p�|ol�۳W����g�:%�����'}X@�m�o���E�9kE���R����9�/�
�AOE�W��g 1�R<��#v�p��9��1-�9�͖���"�>�r��Y��=�覂i��(�Y��a���L���wFz�r�E ��Ԛ��Hw,G�^j]1̵N��� ������G6Y��.8Q����@�� ��G������5|�1>�kIl*�#Ql�hG�D����qc������}��x�9�K,4�Wp���rG�����F)y��]1���Y�T�Jw�oa��p���̉:�1��S&��R��q{��ļ�����{,�*X�Q�?�������y����@7����$�?C&��Ǌ��(O$~~��� ���[m�)<ˣ���#נ��8��3���
�L��"H��$�P���_�u��������h��IT"M�g��n�y�
���!�Wx�����nu�WMƵ���g-���p����#qi��ǫmK�.XQ�Z�?聜<�`��t���D�и��s��e�<���O𫬈opӑ�:)_�Y�%ʢ�K�h\�d�*� ���z1#��Rqհ��p�ɠ�]@J3�$)�Z���x���=�m+�7����0Xx�t��@k�i��c*!�I}&%���
#Ճ�ˑ/��ת{��k��=�UT~3�}>Y�b��pA�� ��GX/BF䑊;��W(��V�����g��"��vy����/����1�����G�RSa�.�<�Y��z��\S����NA{�+� ������<^���P��JA�Q��)]���D=Fb�)4uy��zx��i�������[���h���M��\��0���I��I^#n2��'�Y�g�=x�_��e�yyG����XJv|���4��Ev�맟y��Kuab|�=�ZP�Vs{�V����lm�����(:���'u�4�/?F���W�r���� �X�C�-+� ɘ>�3ô��U�s�W���az��nܸa>�!�{U,ϩ�9O�
����@Z���J���Sk�z��XdB�lf�4e�+ۃ���Q����Xy\�TP^�V�%:����C��)���0n!k�S$����×�"3�O;����v3�7�Z�0ZۼvG�2�"�(��Z���;�a5�SxВ�s�~��Sr`���-?D�b�u��܉�wdU�/�8,C^�rN�r��G9;g͟Sk���&:\�v�>;˵���]�z�~�CGm�B��j
ԭ�W��ʧ�Y�=��y����k������f}ѪH���Fraي�"N�=HΤ��&��3s ��yW����˕����ot�:�9�-)۴G���b�/<�y��Y�]v�h�<-t�'�:�>���+𩁢:��#W�
x6�i~t�|w�\���Kk��pgke}�Ɨ�=�pZ��q�As#)�d,�d���C
w9_��AQg����ƫ��������O<g�Ѥ�N�]�+�nM�Q\�����r%E��|����Ǩ ��e����U��R����v��zZ*����>m>�G�j��a�(O6���Q�s�}7�0I��'�ݶې�°`�@ųXf�{������Ub!�kS�\Vu�G�8K$�OY
'9���s\�"=���o[�j��S�J��[)�������"��龒`l������K��C�����ڈ���BP���!��8�؋�nuy�Y;�(��2d|�n���$C,#�l	�M�┳i�zI��s�>R�V��֜_3^.=�of�8�P/��)�k� �R��̷��X(*�7�z�E�;i�7c��d���M
�2𜆈k,˫'Z�U& j��Nˋ�U�OPft���R{翑��%R4�*=XӮͷ��@��Dv�􁔢�z1�F�Yjg���&�ݓ���tr²�JG���=��l7�z^��z��y߇�)2�1��;zso���唛Lz���J׮|��9�V~�r�t+v3�1fm>p�$�\���u�qκQA�D�~�MN�qH�k�_g4!��������w������g�ciS�X?���_�fwQ��a���T���Zr��l��-J��7�Bu����|����S�)J����E��9����R�CÒJ�Ep�����T�'!Z>E���6�@[���q������O5E�op��ݪ�Y� ��
�Sy����3�w��d5%��/�5���o�(D��C�W�"�hFèc�f��&RH-60傑mh���)$���Yۗ
��cu5cEk_���
�8�p×^u�.uS�(�qF���nL�����"�wȋ%�Qr1������=��J�)�Ù����h�&��g�]�����{#�(�ې��	�<GM�[�E����z�/��}eb�G �_�h�2<���`؂C�2���$)��!L��lf5�U�]�Pi��	��ޜ^���P��f�r�&VFG�$����kc�T2 n���-�'[�$�F<EhoE3k#�.}�-1?W�({a+��a���\�c��W�!}#n���-_/$f�f��?�G�J$�K�G-ި�Y��6!��Tr�huR�no���kjJN������(���$ �����_e��$��뙱��D/Q��@4��L9��:�sP*zW$�"N`�Ԧ���x�L��u!��)�����#N�STn��aMb_*p$� ���;4�&6��g�V"i��j�bkVD���K��YE������%,߆�a�#�ѱ	#�p_M��t �w3��i��޿�9 }�
��i^�c�&��-l��VJ��I��t����P\���]r"������xe��o�4�P������?㩎:��y���͜mr3�s�̨�U�k%�y2h��i��w�"�����<�6�~Itw� ���GN]K��;^ ��Rm�>�dF���K|�����%����m�F��G*��/8���85xg�It��v�J��)85�{F�"�VR�%p1'OԸ��g����&���`��nO�A�D�
(���Z9�l�1w�{ �H��0�� �ݠ������½��F���}��J����k[��x�j� .)�*!qf����*�x	<W[广G���&�[��'%��+���q��qI�-w��iG�!�dv�o51�/M���h_���3v+՗�D'&�J*�&w��ms[�ǡA��"��]-��P
kz��mj���d���[��z�;i{ݝ⽇(�#ha�CX.1�s�; ��3���/O�V�����E�UNt��k�WR���U*i���b%n{$m�g��K0$�fm���My��,AcJ��IF<�;��0�IvVh�TBuV�4��v/Q��}�[��v���=��E�f@�n{�7�m V��-���0��@�i�C��H]p�у����W�/��.�����D3%�1~)�� �<ڦ�%���@���x��t��T*1�y}����Ow�)��k;7�Y�O�^��za�v���犆���7��??���d �9]E*@E����=b�	��A(Qh��JpJr}m�̞���^$�~��)��^c��<�!���F~5���p���1�$�Te��``e[C`h��ъ=>;�(§�E43�9��^�B'�xq+�x��6%'�����er�y�����[LxߙM7Fם�(�C*,�G����|�j�9|-mϑ¢��HZq3�Y���\@�|�&+
fu�D��>����.���e� �ѧ?����y�� ~�Og�ժV���;b��3�f;G��v9`��)�@�đX�J�DJ/�����(���$,�t����=��31o:�w��yWaQ��l������؜��5V���G������B�m�;��Al��ڋ���P�qP�m�Y�������r��F����^m�n����.v�U��n���g�Tt����K{��qr`��t���AL����2�؅�Z;��d�+6n5��u ��_j��6���h�/�v+e��5��2��7���ǷD���[�a�|�7�G�F�%��[v�'멲�nuo0¡�][��d����^*$xp
m��1*3�
�H9����rOgGl��Q�5���X�_֤v-to�3mJҥ<���<Y�����2�O�a=���Om�a���u�.7��y!C�*v5���v�d��[􈘰/Û>&x$r�D��U��-#���H�*�6`Rq��烈X1��^�\�b6&jBob��F�Ġ�Lg͌��S�j?��_��<	���ZI�!��#Թ/�\�N�4=���.�����!�ة��V�o�:��k5�l2��[{m��&��d
�W�h�=�&طtx�
_���#&??�$���!��P1��^��91?c(?a�{�ymO�b�E%���Q�y�I�N9Q�mf�$�`y�i|-Hc%ϑ���T�S'�G��NU�ZA��f��a]�1z��(�Ԁ�M��=*�l�R4��5ܺEO��_�Q�OK~\�V��5�N���桳����g��O~6X�W����B���	0�f�Eabm��'�� ��w�$�B�Ψޔg��|)��)�~l�@��ų�ݞͦ4��6&}�ͫzDf#A��t��^�A'�iMMaK��B>���lG�;�����v��7���ۗ^�~�-�딦��<=�ᾚ���U�`A�=�@�R�(������IЂ�Q��4t#ì���m��*%߾�����{����m�}�����Q�^��kI�֝���{��d�k�w�܍�)�p���bAF�I�� ����kT�F���΍��QSz�#C��u)��x�}[&���,ҿ_n�c�
�Y���PǤ��nK.���t���j�i�(���YYE$H�ﯮ5��H9�e���ǩ3��X-e�F!{T���Rt0��f��]��e2M����K�g��4��<�d]˽~�O�����7K�C��PDk�"q36������@�_�{7��W`PȟFg@�olM�>_��/�H���f��!�������ޛ��S�aHK���.�ܖ�Q���T��y��?�]�����7��[PN�ò�B����� �"c�;&��B8��bO��k���|�`l����/U��^Eu��}ʄ�8m�	��>"��sR1�_�	óEwf��W��!����5����B{Σ�/^�M�;Jc/���Ҧ݋�CT��$T�8��لZ�[B�ʺ���rt���(���y�!�y��f��z>G��̖E9�;��sX�$�a�;�]0��K0�ޤ��$��p}����]�=����&��9\\�1j�]�����4V�~����l��4C�y-+'��n����]�?�i��jh��Fk^��	��P��B�\��*�<�Lo�������b�{T�.I�%Ϝ�����S:�K}�L9�N�/~�d��	�'xT���[��zj4DD�X�	���ey���u
��(#ۅ�y���S��^�ч���x���z�WM���vh՟��~lt^*3�,�eo�2!~���'��GhZ��_�����6�R�ʉ��i��OZ�%���*��W�a*�c#�@.��_�<�<�כ���nAvL������]���l�d2��h��U��R�������]�g�8�Y�UP�V�����X���%I�����E��S?N%aK�ҠӀ����m/Y�u�<Q4e����tr�@pTX�PY�GT��Z��`�n>ܢ	�����&Cc>A��X۽�_#F�=��
,+��U��>��8#�3�vv��X��Wx�!c�mF=��sD�_+����F
a����	j�^�]��FFaT(QGBe�]3T�ʠC�dNg�B\7���M�s�*�LHu�y�;�e�t�����C�Z�(���9�8q��O���������Kr��:�:	u:C�l�c��mӣC����8
��v�s�$�-(�s�h�����d������ϳ�#��J�殉n�|����S���*|�����*�ࡼ3�]ͮ�rC�EY�P?H2�pu��a�����Js`�c�:�4N��K�Đm�2�[*7f���J�n�����t"+�M�Qb|��ư��)e�ϰ�-`��Mއ��"��^i>"c�1UN#�;^�tZб7d}��/w��h�q�����[fDM�B�0m&C (�mWY_$,��a$xA�ly�m�5xX��t}0|�rY���^m�������⪘��Az��s��h��77?�^��z�i�=�l=���\A
��Z-�|= m�3
���?�I�c�����IC�Ͱ�-4����E���5�Q]�]��R���R�����>T�g���2]����(?G (ֱO��<1��wr_����u�ܚ�����^X�2ʔ�789� ���ɿ�U<(�?13��9���Z�D�5���A;{d\�K��	mÂ��+6��#����s���v�]�-i3��k�V�zH)I�yg����K$w%�w�Z��o�_x~*fg���o��6���u>��v��S�a��y�o�6+�:������~v"9��zG�G��J/[�޹b&��3	S��x�zvjؽ(�2��m)�2�R� kT1Y���c?���ْJg�-�$��^DO��oH%"��꧙�yݲٮJL���}�r言���[ۋ�����[�z6ڛa`hy�)���ɑ9>�h��KE���\��tgi<��d��U�Q(�'���}��*��k�2_ ��\���{=}=�E�`.�2Mi�5���Ct�nq�Gbb��KɋS���y���Y@#����g������Qg��{`�~�����~�\lډQe�$�w�ܣ�(��]ϿTC��>�=A*ܴ�ǹ��fמ�hO���iTb1����WAT?B���gt#1�p��`Q�[��V�B���G(����atW�Yf��aB�\뚪=�����;B���ʁX����B
xҎQ�+Ȼ�,+#1�������M���W��K�MP������p̛�8a7{�G}-��e��7�� �3ן;�R��_sn��iɤ}y_8�$h8��$��Ru��9K�sa�jP�[��*@��iB�*�H��<��
S�CP/tR�a�ń�?�Ө8!�ju��:.e���_��;&�b]i�i[�i�����h�y��z��(1W!P�C�F�n�8])��l�E���������/3�&�$A�	�1)Ɲ�y�VF����WA�I��,��L��يJD�毡!4��큙f�S��?�o�� 8�9��s?�Py�X=���)�8tw��f5d�VO�F�A�~��
Sl"�أ�bx���ys�g�s�o&T<���F���>�����}C������*�.}o���q\_E��u��
Pt��0�[��'����~̘���-g���]6�X���C7�@i@�︆���Y�g�҇��Z���b�G!��kn�����/�Iҥ�\�l�-EN����2ɲL�gy+w�Az���\�2)�gWXza�m��Xۗ�+��M��[2�A�0k�Cs�� C*�/����^E�Xo���n���{����s7\7�~>���Yq�^ ؇":��~�/t�]B}�Gg;7g�k���n5�HtR�����uO���H�\��Q�ٞ?���2�A��W��BW���[d_�Ud:m��A��b�B���&K���.8�t�v�{�b�d2N��O�}*�����	��$����k/���t��^�����I���2�w?ѩi��ZXO���.��*�wԷڂv������ܘ�KM�?M� ��' _y�[ma�+_rTG�)I��?ޯ>������>�el��ͺ�9�P1�K&�J����`\)F/ "j�,ϸ���]�ھ/���W#\NQ��YeJ�P*(.%zn5{VG���<se٫/�+@1��`vf��ᑤ���):���A���s�W28���\q)�_��lڬ���{�����?P]��$~������Z�C���F���53���H=�2|�殴�qa�<�̐D�>ôoNa��V_(��o<6�R�رtwy�g�^����51��J��6l�T�\a�5g�����K�ћ����%j6�A����]�S�;���[�a�r=�e�yk�;Gx������)�/�@<���BT�F=JV޴9)�q�ꂣj�.C���465�N�~��{�}Py��&W%�ԁt�Fi��w5��Ao�*�59�����:ə{�,���Ő���P�K ��U�y��[>�3���39 S���kJ�ڷU��Y�Z����8N��o�����`Iػ�R���Üz���+�B'(^_G�Eo�Q(!��c)'+�8���7x�R��G��JF��<�ps��y�4���]]6��0��Ñ��)��1
�5�?$�g�Z�轭ء�3s����`U���10�W�B��D�O�1�@��H�u��;�R�1�tu���%f��:ҁ:��-^�#lQ�������Ic/�6�e��!���h���uv2+�N�ۋ�ad%�w���y�n��,���{AG������3�3I�/���n�I��Q����)p z籊���_�0ر��ٝ��"�%�vr�ꠚ� C?�^0���U3�)��x˰Fɏ�M#}y��#p��Z(rf���ݑ}#���<{���S�8�yw��u��x
�m�q4���ƛ-n����RՀ2���M�=F�S�lgmVCT���ߛ�9@]�����յ9�7�{˲����f�l���������¡�ퟅݎ�U�'(�w7t�S̠v��������+����*?��h�½;��o�&���=�� ��_ a='��Z�]��2�g�5<<=��p:��(�p
K��_�0�,��헱;�^��k��Y��� je!</�6�%�G����iك�N����{\����A}�����(a���Ə���φ�Q�T��1�ӆk+��Ae�f=�7n(߽��&p����'�x�������7��T����@�H�gkKvmu�ضhj6vIA?k�����_��FVmI�bt#�� GE�vy������6u�(+Ai���FO%���:��F�����#���-�+5�(+A닉o�
w�ID�~���w͊��^�L�K*�g��^����\p��ȶ,{"��^���X��8y�烂k)��й��� _׹z�Wf�3ul����'m�;{x���r+~�ܲ,������d���w�%7��^���G��+����{����/��6����N��h̨�[X�zu�ɑ��D��9>��\�x�Sv~��XV��z���Kdj���u*�IN�0d�3�j��U��|D����V����_��Y��Q򌢴a^�CX����TU6\����A��x��!�̆o@�����~��כ~%^[�o�"__o9k�D`*v�៺2����p u7��́nf�f[U*���D�&�]Zz�{ʪ���HR�j'����F�R�8kD��X���?4y�^QM�W��AE�WZ�)�9�p��R����[����z_ZeS�qE{�ŷN�J}�T^!`��(o�l>u�`ԋoGA�3X�,`�fg�4U5�!�)򒗄>Ӄۭ*|�cT(Ƕ>��@|ƞR�0�ާj?-�������>��W��f���ޮ'��"��nli@U��l8o�S
��"T���n���w(��kҰ�e%$._2X0^��ŗ��/�pIw˩K{@�rWp��30z>�`��w���9�[�������h߯1���ǭ`����2�Ɣ�ڐlS�򶭁ٟQ&V�]��G���n�3r%��tyE�8.��U��� ��yUϺ%���Q�+�⻹��U�� ����7�o�G	Y:��$�b<%7�7/�s ���Є��,%�&�s���)��%9�u�#O��o�ӎ/5�
L�w������{v'_@���*\�J]���6���p�|�4ۅP!"��wn`��=,k��z&ܷ�S�գ=����t���Ģ.��f!�E{�������-U�7�,��+���[X9\bZ��_{󗸝�%Ȧ�.Cc/�:�Y<�o��|	��R|	�z��Lo(?�﫟-L�Q��Q����N~V�x���"^��גr������ʣ{���e�r}3K������*��^�nO�;E��X�3�!#�&�h��̇%o_�	�!0�����X�K\�뺆�	���(K�FY⟣��ˬ�	~� ��N� s?��d]�,��U���jL*g8�1���t�z����<$��u6w�P-+�,�K��\�1V�G{
%�����U���w� �c�º[J����]�Oo�/8�����Cp���l��Ycl�~&�`s�!��xV�}g�/���s#��IC�ߝ�I�B�{x�B���uE��LV'��f��4��j� =���@��承��p�[��ط�溤H�����/�#���-k�I�[q�?!��gۮ��㈮�4��� ����1��{$�-��L	Z{��Tǎ�tH
t�u�E��x������w�0ؾ7�~p��ا�^��N�r+�g�?���$�kQ�\m��{����Q�����k�e
������Ҡ�:�kw�S��-��_i���Y�LĦ����7���e$�ύ���<��ب����J�Xr�WÎ������M��b�래睜����!�ԗ1Ihr���|ex�&�'+Aqf���!wɑTvnu�#�$�j�pg�02U�i�z(��X綩d��<�?���Hk`�U~�cU�uvjx<��0���c��s<�G!�e��S(�?N� ��>�v�fe6y������� /ГR�x��z�$b6�WI��g\�Dſ�h��5�c�g&E+tx��w���,o�Jj3�!1�5�����W�,~d^��-�1�V{��j����뇵3Կ�bY�V���=���̼�>�-�Լ-��R�!.��9�R%KǹNO�-��禼�;�y�Ч�;ū��#�u���}s_�$}�Bg�qj��~m�J�%��J������}�������9�����,��Բ�S�e����h���tq� �
u��.ժwZ�c^�~O�ҁ�G|��[�����õ:��6�;�e�K7
�
�f�?	(��!�l�B�b�����o���ޑ���p���؄ٯUT��Չf�H_)�{����f�,R�Qu�v3训�?յP�>���G��_,��������U�NA�����k<9k>���2����� ��K�˿K��d��:V�P^xX8��87���ء͖{��+����uzsW�����D��q��e�{둕��!�pJ1�d���9i�п4��c.����.q��\�����|ol���A�BgZ4�W�(W�g��XI�\=��@�T)�8���N�'�Й�[�W�w6S��܁�L��ЛЏ�J��s��'�G8��
��)ª�$�5�W.�N��<��sJ1��.�N�J܉�io�B���[�S��i�ſk�S�yq���;���q�+z��ii��~$�������v=;#h��Y��y+ �6}u�ɲ��C�3d�����A�n�����N=-ۭW2���u���f������=���s4��)��_���g��~�-q[��g��v�f|_�\�����JP� ��5���$��M�u�R�r��3?�qGG�y-=�H�0L0�?�p�(z%7| ��N����ܴ<M@>UDB��m�sQ{���'E~��3i��8���=t7A^ʨ8���
�qYm�p9c/�B����ۆX�(��L�8��8�ڷ_�)fĤ�/l�5s�y@�wH��B��$J])�ԛ)�X囵���'i�� �L&��33�K92�I��q���=��fT+���bc��O���W�w��%�4R�%-nW��n����軌����3+��k\n���uj|鸭�wrBi�_ެh�"w���.�oE&���s�]�!��=s6q��A���D�zCAK��`�2 ~s-�Ι9�5�P��)��Q�r�r�N^���� ����~��.��H�Z_2�@���7�4��L
��.y��{8�\3��57�!�3�ϗ���zHg[nn�$�Z/�6ԔG��k�G~^�|�;�l��7�3�� %�؋�-K��|um�v��
���e=����q��Dx��	$k~�����/���ʲ��*BL�����
�
vE�-(>�����|Y��i(��_@:��xv�$���"�C�����Wn�榊�����:s�e�̃�H�e7��^m��$ʿ;���Z����m_'1�@?b����#}8�������X��1���H���F�Ia�+,Sy��^��T��CC��w�o�/�E���-p"8Y�-��@����n|����0�a�w\k�WF��8yVH��m�� Ct^-j	�^Zd>����H<��<��m��WxL^��Q��3?�1"�_��1�_�56.�쉮s���	�@^��"X�*�K�f���N\)Ζ���y�)$NcS����c�	q����H�?n�Ϧo��|V�3X��p�m�]�n�d��́�����*ob���j�?�9U�)������0|cxO�f\t��&��Txq�����T�H�q���8�#>~�m��_)�G̽�����Fp��i�a֩�φY�s(����Ƿ:J	A��9�7A7Ӕ��R�����W`��3	F�@�RqZ�)a�k�:,?�����R*��|��N
1����R�����%��� ��{I�Y���1�[��Z��5]�c�c��kBj��7!�o������Υ���5�v���Oi��Y�� �D]N5<ZA�ʲ	@�R�Exʎ3�I:L˓�9Φ�l���ײ�~��.U����-��CG-<����}��qRһG=ݬE0�J�ν~��H�viI?�ֺ�;!�Ȩ*�
ߌ����(	��{��U���3/�O�0_dx� ��)���H"�!��y��/��VRF��S�Ђ}�����̏�wLwhD���V�H`Q�nsQ��g\�e��a�19l�UD���8� �s ɋ_������>�������_A��4�a�4�yî}�zm|���8}�����+Å�4a�>43���m�ɒ*���u��A���ϥh��.�{�6�	�>/u|N�:PN��0'@�7`�v>C��W���5�s��A�/#�Xm����"��(��gA{;|�kŜ��DeU�P3y���ء��0)�Q�Lt��������վ�4��8L}n�t��;$0#a��4ɨ�>3����>6��'u�'�U_ѣ�P+ŽlY7��s�F9X�y���Hj�]�u�`���ho��yJ�y�1�!�?�Qub4�35�u��($�sL{�"(���2-��&��|��1�u���z��"P�H/�0�� ���/��
ƣZ{���ӯJ��c�[�����IE)tA��D�ߊ\r���*���3�-�TnI����f��.�m�w��n66�����`�=o���yy���շk���S@�œ��_-ގk����W2�N��ҫ�ʘ�q��4�jݘ��S��YV���_$#Ӻ�<���7Jm��N��ʽ���	�ΘbC��M��®�t�<��\�	�+3��S��pl�[!1�0�J�d/��{�&?7(�>j���KߺZ��~��u��8�廇�,����\�������>,
��-����e�v��A�yM{����@��n��6.��8��읔�p�~��*^х5��}z��w��I�PO�vI|�K���2[��6�JN�jDq�����s>��^���"�{����)���57�
�J�>�4��a�Z/�A�pC��?{i��qԾeZ��tm��o��p��|�YLw��a=t#zp�	��\Z�A�-�8�� G=��wc�=&Y\���B/����g�6���*[+�B^�G��RmM�"Z��B�I 7�}�4~�#��>DR.�x�����t" ��`�0%�M�	#'�#��S��{m�M�k{M��mא L��j���K D~��A߲�P}������|>�y^f��_Ȅ����:������_,�
���2w��ʥ�8���F�Ӧ�$�72����
�q+��� s�����=��z�qN��Z��?7p���{d��+�9寍��	8��e��|�=�_uo&km�+qC�
�����H��}د���.iD4,��GZ=���}Sv�Y�mJ����c��)MSJ{�F���	k���ő0�О��o����n�{�V�����z�D�Ck����w�]cqЯ�nȸ"J�2͗4����f^��W���!�ow����M�L��r�E�A���nC�R-���Q���5���Ehl���웲��p8�/�X̞up	��
��DO_�fj��Ɇ�V`w����^�i���B��
�I:�i��|�9܈�nк5zT�G����V�Z�YbV�YT��~�������
ň��o�NWhmWj��z.WF}F�?vx�:q�[��S�t��U�.�@�9�tu|8w�6��� �����Y��QU�+WL5����S[;rj|�i8j#I�K.��%�&�zD��Q8	�[�>�<�K�H��a�2�˃�i�������p΀�t+pe"�c�DC���0=O���	� ��Vо��5���X?��ƪ���6.�d*�6:-�#�&fT���b(Uu��+�s+K����o��hس�nj@���c�K�D&蒬��K�v◕F�`��<U�Ul�)�������}�_Qkw ��3�X�֯�$���kH;�-G�T]���qw������	wx��0<�Nڭ�u��q-[�4�D�
�M���f�wv@�"T����3=!O��т�wid{x�¼��r����y��D[��Mj��6��>�/��0��t\�}��l�B��5a�c$O2��ގ�A4�k���]$�P[������ܯ�y�Y�-4v���<qg��,�g��D�4�=$����,
�}0ݯV��jޝ9��	ZOV#��Ӫ^�0;e=M^��jCk�)۠<>�������>xm�^���v�ab��Zϧ�*J(M-���<*
�^����Z���&pO�/Y'F�f�h�
	���(�ӯ�`�^��UMCg������]��(�6��s��߶��6��{�fU7�o��Õ^���z���@�����nf�`����Ik�E��n�*_��P� ]ŗ+%�dְƇ>O��u�����$���GE�ή� �غ��)�J�i�ܤ,�V�10�]�F�4����-�ѹ��+WM��-i ��H�ش��c�HD3��e�U��0>�0z��1۞����y��hq��S*��˧0#`��3����w��t��2����H�X
�z�<ӧ"�A\���\�����C�8����������vv|��r2<�>�X>D���
/"�q��X	��/�~7b��	�֫�a��ղ���N�����y˵��aF�u-u�z�"&z�Q�B��`����M���F;x��P�	%,���S>���p��JE�>W�}�t��X�T���ɿ	,Ê��Q�}ءj��L"U[�s�e3��Q�o7ܹ'cK��͋_���.�e*)�_��yB@2I� Q�P��<O�)���7#�bw�p���\F�<��3+�g�GR�,,�<�[
e7�薆,��xu�ŭ��y��U阖�>�@۝粉f�����g�˟���Lh
�u�=0�O:h~��Ω�Y��;�R�eK|�*�h�lm�kA�у�����,�&�?���|Y���/2��&k�Q$U%��93Hi
����Nl[Lgܴ�^�)�� �&f�����$�YfrE��M|�!��(�LK�p�t�F�)�JG=���M�'�M���U���p+��V�qݼ9��ç�Q�~�3
��Us��6�t��o������*f�� ��Ӡ;�ڡ����n Ng}�0�H��Zyz����Hw��E=?l�T����Sl,^#�+4��I�����$���y�c)\%L0�k�a͵a�d$�4bIiq�jЖs�0h�������r�u��}3�*�ګp[��8i�a���F�2uRU�m@���&�8��Ec���(��n�j9�E"s��N��q�d�:�-��lx���ψ{�L8�~|�lCمnǸ7+��0ّ�y3�I�}�T����ދ+��?����?����(��Z�"t��vt�+�m\t��#y�����?lR�o�@C`�ݮ:bv�� ��Pd'��~������1���	�yk����r�/̂vɜ��Z>$��lt�u��1c�!�t��eVU��#�t+<��ECXbc����h|%��	l��ô/ ��?�|��-�<u%��u1<�����wc`��[�*�ps�4���SzK"9�E>r�K�Qb���\k���
�㘰w��`.���sY�hֳhi��VM�.���Eq1*<���ƨ�I3>���w� Jv<���u�z�߅}��$55���%�Q�I���	
P�f�w3�����g�l�ߙq͊~J�{5��71p���ZR��4�Jdb<,�0ۦ��r�!t����Sf�� 	����-���;fK�Y�7���n��9Pf5�p~��U��Qowtߏ�����h�ߨ�ƧR+U0���h1I͙3qq�E�=�׫%�A�ּҲ�fS�#�(�~�f�<��h�V\�8�F^�b�:�r�P��f�$N:�y򷞵e6z˦�<C�f�D�h�Yt4�%��`;��&3���Ο܏)�����"m�|�3:�r�w559e
6�Jճb�i����9<�\�����v�j~Fh:?\]d,�.��#Z���ּJ�r�c?�`�¶���ƍn[�����`���G&��	sg%�������V:����s3fuЂ��"��q�F6eBCi�і5̈=�>$E��ne0�]4*�$��t��Z�T�c��yܱ-����J/^&u=�p=��p����!��e�,����Hm��+c�58�J�寤�bA���!J�9�Ѩ�\�M!�Z[���'���>�@b�cu��sZ'��{� H�~���۽�<��V9uR�ɲp���чHJNS�#d�N�b&�p�T�P��l�\��!��\�F�n��8t0lڻ�$i^����]^卌����C���3�2CcMA1������xI_�?2O9']
p?������p5��V|4�W�ݝ�1�n�Iw�:���}9L�����
�-t� ��~�ͅ���ͬ�0+)�ܴb�}9�sV�;��۬O4��&$X�F[ƛ�T��.��1y������Af?��N+"�I��~S�Q6N�M����F��]��R� WKğ�Yi�҈/\n�P�=�D㚊��En<ڭkfL�nE>t � ����3�Ϩ�w�,kY�V�?��̙�.���Gy�p�M�u�t�7JH�!�#���g���'�%����y�ױ��ԫ���>q1̇�B �Abu$�+S'�{�L�N��W	���Z���]��LqC��y�x���*�vw]`�m
u���3�G0�
�$�~���W��}�y�g.�����2ieJ�g[�;�B5k�dk?�������^~����4�Gm�R��p���:e�J�L�+�y����z�ʟ���9'��xA��=�͇g�� T��ڽ&�(B�hàF׀t^-�o(�Q7{M�3!����tw�`׀b>~�����B0�9Кw��i׶��P�掀HzP1?�-��ea�W筮u3M���)�׃�A:�W�g���<^~Jq��I�%�q%�]�� �~TN�F�*�T���vso�E��:�=�@�1U}�EO��N��gR�E�	��&R������Z�ax5��$&ihb����{�	��SCUs���?�ǽy��W��f�u�oh��g�xG f��@����TAc���YpL�GD,�ڮ�B�J ��W�2�+�#���=L�ιY	㪔^S�?�A�x���6xp�M�����
����YoKL戇�-�o`�97i��4��x4�	O��߹Z����v&M��"k -�#�CӨ{KR70o,�)�����es_�N�x"ǼN�/5��֕aXTb���ZN��
���qr��o�d�9���y�e���'d��1v=�]"*�A^R,�~h�Ra麗�!��(޽i���G������k<v�@�Q�t*�uu�L����#����̟/�v�Z��a�pp�8��S��C� �*�c{�����
z�U���u��Qa��]� ��� �v�n	W�1��9 ��h��4RZ�G�9_�9�_ɱG~�IH�.%n�)��qb`j���޻kZF4���<��t��,<��F�$��:8hz&ϚV���N��GvaGlA�m��$���9����̒ݲA��}�fE�����Ē���CS�=�P8w�%o�X �i����/I�Z8���z7T�H�u�	u/U����U&��b$]>��l���Ks�/���K���1�_bmhy�<-O��>2f�����i������A���eʯ�⡢Z�TRx�2��������V��M/$��vCPe���:d�2bO�vu$���z~�<q�W~]�:6���9�&��ӳ��=�22�)�>�ao'=��}W�%���:5�����t��.����^n�z�J�cM�Ug>��5��.<7�n��MW�p�@OP~�+�*ީ6>0���x}�R����/��X��Ya!$p'ҰŊ��ЮI��\�Q���
�K%2.��=-4]p��h�ZyRM������ｖ�A��<�#�ppYc�=�I�S�	�֮Pq1�W9�k�v����U�`v��!L۪҃��4e� �C֖=�15���k��#\��R��dP gt�w�N������͆�Ǘ's�;���e��3`<�jl*@��xd2��Pa�6l���6�>w7����;ƨK�o�R�fp�5��^�%U�̟'q����Ȃ^�����b/(+j�)n=4��V�e���(�����9�Zzz ���:.�#"ݜ����u�̿���U�.K�!��
N�D�������WD$�
d݀��V�>e_�Т˦%a�f�p�a����9���'��y�]fKLn?��|������"8V���|O����T�7CN�U��ݑY��4�.�y&}COM,|MJ��ּ���tG��R=d��D�nʰ�/k����=@�f����M���"��ϰ=nW���_�Y"����W�!h����ݳ���2O��v�ԛ\>Ԩ�kJ��1�����b��egr���w�Ŝ~�f��+i���u�c��5)o��H��U��Ž�$���P�-8�[����+V:OW�]!�/ĻZj)$�_�W����#dH-%�m_
p#/˧����Z�<��T]�\tc&���E �*� ��p���$v�'7Z?|���e�[�n\<� G��T��7Z5%3�Ft+�i%O�?7�[2��;�%�����5�ݻ�ء��K����
��g�*��j�ۖ������Al�%'����BA�ڮ�n��G��1�����_i�+2�nŸ�@s�����I����o�'����J�*�)�o�=&���)�H����Dy�[�.��z�r�v8Li�`QC�FZ-N�2
V��:��mЪ��B���uY�
�NN���HM�D+�]=��ſ��	g�>�|���]/�fѽHW���CevҲҷ~�I5Y5�ý�.�& ZEi�[q�ev�wR����WG�h��b"33���{�t��
��i
������M>��/�Xqfl�\VI~��lm唸���,N�bg��v�,��f��-m�;`A���d��k�9پ7�م�V��Q9P��d\]�9��]���K>=��W��V�ꖷ�Dɠ��1��rB񺠾�U��[>���P�_������<�#	��Y���,�y�;�B��bψ\����c�R��Y��R�Je�LW3�y�1⢭I+�����Ւ97+��)jjE����jo�c1�%�e��gN���޷*=��w�@�'�T�d��Mb(暴�N�}��>��k�]�r�ԋ@~&xD�G�N%O9es.�M�.�ie��Q�jj��nc�0bo5�k�{��V�hgԮg6�{w�FD���WQ69�x��U5����+��T���/���a���30��^^`A$:��aʃ�8��%�����a ��ڗV}�8�-_H��s8�j��!q7�6�"8�-).��ܭ4�q�w��;lH�`�w�Re��������o�!6P��%V [�����-Z\���v�bg�p�+܌&;����xH��A�%�G�E�ŢS;�*��]N�&I^߭	N$�5b�F�>�@�����w�������~������%'��ܐ~�!�徚G�W�soŔ$�G����g#�%2�]�%�Q��D��[����n<�ޘk����
�r�
)��ؑ�jw�y�T�m�|�J��G�J�_ǋ�z� 1u����(��C�mY�t������A����2�䗒_��?�����P��k�֓�i�����eg QC��\gB>,��/�Bi2�~��#�Z����߃��;� �����1+��|�E�!���l��[y�t�Ή���&����U'E\",2�k��)5h�0�]���1��S�K��Z��Bk�z�F�T�y!C��&7���k^@�l�5w�.T�m�Ò��t<qj����_�'�=T%���@�uå"��N��Du##�6p�q�{6Ӕ]�Aف�]V����~P��1g�0!Lk���4�󀒣���:v����YV����q���d��")8�/ ^�w}��U"T�T�$�w��T��[�5r��B _��sQΤMz�:�Z����S�K�P쯇��3K��ۅ����K6��l�fkGA�?lZ�b�r�v s�]2�߁ϔ�����U��c0 /q%�cDu�����`�J��*��"-�������]wG��<�{�� �>�n�ާ&{#������{k�G�Wz��S����U�SS·Z�.���i�:HQ���L^
V�R������7���{j�ΈF=2�Dᙎ#.�Qd��;t�]Yh�p)������=�"_��
`���:����wW]��A%[�bO�^n�"	l4�s�\ٳ�^te{���z~x����"9#I��Y"<��	��jZ�)ů�B\��L�l� ��y���^Ƿ�1&���_b�;���)�^>��(��\D=»M����	6���q�@��c��)�����/�Ctk�b��#b��i����'���'���s�b�d3Y��K��@��37<��������%v�9��xO��{�Y�_3�k7GT!�ǀ��;��kj�J�1�r�G�_/��qy~x���DkL�X$�ù*c�,*����q�����C��yr��/=h��z55��6��%'C�/��)��Y�K��0�ܼU,��P��ʙ�� Q��V!e�ba}1�h-�w�����r��#"�R;/x�����]	�\{9d?BϚwM�0��2���[-�0牨�a��\}����m�0����T^9��}��+�t�꺶=��7y��N�s��e+� T&�د�駸B|�}��I��s����{��ꢠ�ּ�(>�˂�QS���TYh2s�g�nݿHg�#o��l�C�Kr۷Uxc���S<^xj�LT3�T)��*{��y�DZW���/&�mT���N����p��ڞ��>�Ľ3��hȂQ�(3!��c�|�!ǜ��	�1�|����m��,��Ϙ��zL�t�-��ɚ��"+�*D�c�����3�(N�d(�����v�����T3�\=���k5����O������Ԏ���}�F����t���w�*owTݧ�N�jϷ�R�?3k!�T�C�mb)v1�/�Ű�}�zZ�����S��oт�����b�-���C�� �m��>J��O��Hr}��R�R7�,����)8*����F;TMc�B�BUb�TkiA,���Ѷ�7��|�;W(�T�|ܲ5QI����B�����l��4��G~��W,Nq�0�$Ta��Q��%����T����m�+3��G�q�z�>�$$���(���F��A�%ڐz�I������<�5_��ִo=r�޶��,��?���V��_�0���l�h~+�F�Խu����wN6QOk�<��<qN����ep���åMf��*GI�6+-�u��"�k�D�{�$�\����=�ygC��Z�^�����d���<�1������w!��9ݪ� �3��;��ʽ��<� �-�O�?7w�Y:�o���?%�_�<M��S�Q�6�dT��Eo蒮�5WD�\C���455*x&��ZĚ_t��H�x�:,)��,�r{��z��h���oΊng~�Q����*﷪X��T�GP4��Yk�\b����Sʪ�a�7�����t�6��rϛ[�mJԺ��4�)��"723!O�����ˮ��=Z�E��|q�*�������������V��I�cH�嵽x~;!g��#��{7���M��#���R���ǖ�l�nb�� Ή���݅��.X��8f*a`*��
�wC�� ������aI�JK1�{,~��W;�wq:W��w�L���'�k�'oB�ӑO>3�3M!����M隇m�a�Y�l�ݤϋ�58��O�77���U��?Y�9t?3»�8F��
2զ��h�?��F�{�?��(���ޚD�l[j�L�ÉٗO�>�dm~<x�vk�[l�"�+(�"CwG�t<�X�Nh>,L:X���v�C�%�浪ϋ��\�������N_ ��ٜ35�����j�/p�^h�m��{d(�I�L!���L?+P;�Ny�;����RB�(��~{b�3���a�x|�����o�s�ܮE���r��)?���rI��Ka)G�ւEC�5�vZN�������#G&��g�n2n��{e2�g�<k���n�Xxκ�I\��A*8��W)-�"���Ec��*��ؿ�UuѪ�Dm.Zl���Y0�W�S[�"�dq/YS�r�4���J�/{��#QW�w[����@U���Q~?����j�9�}�'�3!�r#�eء������m�ҽ�X+׳��e�m?��Af�SfW���G�c�j�g�qH
��_��Jl�3�Ü{�k�k�R�(P_Ff� �5nټ?�VL��+|!�}"��jbO����]������o�W�u��Y��c��o�
1U���H=�/���}Q�w�zԓXv7��=%�d�Z��k\s&�l�=��vô=�Q���Jq@���;��K���y�/.����J.�'��~n�οiW��<%e���f�X�>�T�(Z~?��L�Cֳ7P��xҳ�x9v��W5��x�8_�#�W����p��Ibk������~ďęb.�dT�v�k�S�Lm�z��f��@`_��l��e�����jTL����;b�rt��cuxke���o�{���c����V��`��~���$ϷU!	��d��q�jdGJه=.@JJz6vܡy�����[-������}���w;;�ب@����WZ"3t�2�]	_�k�	�q���Au�u������(ʤ�ۡU�N���ve������gfS��T����;�4�'ǂ4���^�����r�?Ƹ���4`��c�%{$���EY-:�����9�SS��2鼝����(C�6Ky���>�^��'�u*lRb��$'�ePe|[,r�L���(+*q�X���2�.�Z"��p���T,&�J~;^���H�*�|5�Ǧ�2>Őn�Cͻ�C�HW��R8���԰�y�g*���>���FJ�M��Hjac�(�]f�V�K�dٖ|Gm@h�~��ge��GC�0k�m�PV��u9�rQ<��JA���@�[f�B��'TaN�p'�uԳ�,_��"yE��0�	�x��y:�C��������LWDZ�?I�:,��S�����]�����k+)��:��$����L��儶�82Gfx�A�[OzT{�|Y'a��M",�<�[Sfz� �ij0:��ͫ;H�sAV�G�H�p�!&���J-�z<��M�����xn`bpKqe7���k�ZR?��g����K_{(�������:ɾYM����Թ�v�D�5n��]a��u_�C���ez��g����#���(h������+93Q�q�Π�I�{ʐ5���G���o��p���2n5����O���P���pqC�z��h����~9��t29T�-��a�]��+{���a�����F�_��Ϭ}^�@��'}}�;��Q5�n{eeY��x��2.������E�*Q�}&n��Ģp�����u�<�_���#��w�R��'���n�\���^�N7]��D<�����������g���A��Y����_�W��2Ng����^[�i�<���/t�E��`|3��U����Ծ~e���=�������Ji�M]tJ�Sիq�č?[��\2��?�S���0�F�d���-��j�B�!��Bē����Ja%u���0x$��0����EB����w��K��'_{x�j�<N>ξz<��nW!�ٻLt$w6��)�h���y�#�(^i� SsCJ�EcE��|iJ��Y��9�S��݉��[~�_K����ez��%F�C�\v׿~XB��ڂ�?n��rI�C��[]-{!
W���5A8�,�gN�$��� �S��	�#���JZ��B=:`{�d�f%�(�ʬNac�j[�S�-��M����-�����Ű��ѫl3=��i����KŪ7�.!.������y��}�~6��&�n�ϱ �V%�X�{�����du��#��>�����7���?NG@���/��SK�"�2Cϓt`��޵�u'�C��F��sth�g�p�%>���2S/x{9��o�H�BI��1����h�vW�n5sx���E:��⹺�F�]��G�����ȸ��Kk�V��"���&[�S{DHm�PG�!�#^�bǑo�3詳�
���V�<�~$G�ߖl�o�w=������B���) ����|�m����L?�Kg�M��p��!����N�1���}�����FM�L�X�L�*a5ȇj�C���ԕ����4
�<U	䌂h-�Zo��.�xJ�{�����E�1��k�3��$�r����>��V*pOK��?� ��,�>dg%M�����pO�:�!�\�ӻ�$g3�,B�vӗ����ͺ�4�wV�G}%��[����08����&��zS�-��%
߹"�g-���p5�V�f�$J�~�hc��Ƽ���[�8����oK]�Bpi8��e_��־�?/�	2w>1?��%\$U������㋕����Y��y�]���T/qr�PD{�^�K��#�0�K��$�il(}lZ�v��þ�=3t�?��2���vj:��F�ǽ�D2ޭV�PP@o��6�	]iy�����!�xL,��E�Ae�? O���c��Ik���:��)�	K�hg	�8��e��oM�7�_RP�cp�����OK��D��5���m�W�B��KAU�~�L�K���Sm�&V���%K���]�'����4�u!`���s�Ç�7��0�Ŭ_�k�8o��d�����s�%���Fr+��K2j��
�*=�RD�qLkͬ�.���8e��U�b�%�G��{�;�O9l��EN�9�i�O��*Tc��4W� �V�}�Uތ�2�T���cp)!�(�W�ֆ�m��k-�����}��0Wt'
�#���_��bJ���~���KO�nr����qE!�~���3��e�ɟT�����I?5��8��{�;ߤ�]��s�ed�b��4�r�RZ{�fa��)���N�ZJ��^���ڏ��L�AG��	�x��+~ �y�;�5q�����
�-���m^�qG�7l_%OB�V	C�L�GQe����5VZu���jȑ�U��_��>��'\�al��^�h��<�2��,*3�u%~���N/��U�Gu�͎���˰rDK�>��c-�y�˻�FE�
��p���������L���,K�ݬ�O[%�3i P�ɀ�+�?��2.:Q���T���A\��$�_���-�V��o�p q��%[�|��ԛ�����B��sF[= �X�8S̤��ñ���E����ߝ�4~ᅝ��&�O+��i��ݜc�<��c-�Zh�/�aW^l'��F�nT|���Z􋿩F߾�wP��;%���N��� W&B�Q��A
�dd3�v��Ab�:�6�X>ޓ�$T"�(ì����B0������+�}�\=�%2����N��|��Q�SbкK&vR�s:K�w9�O��c��C����%�$���*등U��ٸAzI�̟����r�D�#_��À�`�aQi37���������al�e�'����>��� �T�ব���l.���3唝�>k����M���ﭭs]�X�w�6m��F���/��f�$M���=�2�&#*T��!�>���)l
Ye�?Gn+��!w��u?{r�luC��uٹ����f�4�譬��f����`�0q*^R��z���M}�lݾk�����m�:j��q|=��)va�&�]ԃ-W�����0v�y3�B�Tw�<�fb�t�M��`WCLZ �~(B�ޖsU���έ�a@s#+��ڢ#m�&2�H�zK#=����~厘2����L����YYK�@Q��:�uuؓ{%?�����Z����/�YJ<���R��n���u#8��'Sf7{�5�\ʵe�~xc�'z���y<x���B�'�m�p�:?]�ws�V�����n�\v����^�k�����l׬�'�?*fi'^�G�xP9�I�Tp�5�"L�G�o�t�s8w�m;��5��1fUy��bu��$��$�~��P�C�|��\`�e���B�g��K`g_��@Cb��c���x�׆��Y��W������.��J�.W-|�njPrL��H:t�2!u�A��#������[�6)�wm���O7�Z�z���ˋ�s؄����PK�@�M]�<,����u�p�z�p�V�>@��B*;'�����ǃ�i-���OEfj�EYF�x�[<�p�Vn-ss/D�L�(	@+Ty9 _K�*�|l��ِē�}�hF$�̥���v�z^��j(�(��qc�r���uU	a�y����o�����JDӆ"n�^���#e�z�Š+����OT>��U����GIu��`H(�Z^=��ВH�,8 $}D���á[w�����4�Z�&&��w&T�aַO�.L��y�#������i���X�sd�~�9<�[g����2mQ��yP+��5Th��߀��s���ӻS)�r��En������
��q��OH�(<��Ow��m���	��H�uSJ�~ݨ8��2OAd�$�/�Z#ok0�n�\g�8|o�����7=����u�M�	`�}ӹZ+%y[��Hlwu�`�,��"�.�&���[����?�ܵ8XWOY��L<W7e
���{8���M)�Y�
���}�XÏ�o�z�0�(�3�ڟ��ѳ��J���oh���~��z�����������}9��z�T�{'|�dPj�0U3�MB?C�6X���l5�H�zrP���] B��6�L�=Q�h�pF�/��b���p7�&8�H�-,��Vu�������4��֫����|�šM�?L�GBE����0�p����K�����P�DT���إcZ��R4���[��F���eTi*���d�5"�:S4����S|S�!�և�[�?�2wy�)ōJ���=δ�Tg��V��g}<۾��յ���SPD�����#��L�z1��m��v�a�|UP�g3ZpOړ(��;{�C�[̪r�â'O���pY��ZtFFG=�?��A@��q�I �.�xX��~ֿ��o�%��44;�*a�>�w ��N#m৿�B��]hk����O_�8�ktB���|ٔs��,�����Z� ^�� m�D��Kho/X����^P�"q��L�L^��;PO��n��tG���7�y-C�-�7W�
ݨ�	r���m�6U�H~a\���ݯ�ه���w#o�Xe�cN��ޥ���<i7�Ӹ�q��t����̣�I_Ğ�{��^�����ˊƖ�.�|C]M�ޓC�	��F�����z��ҡ'�F���UQ�7����ޕ�R��Qj/&WD�9Z��`|�=Ҧ�o�O�h��B��UZ.>x_��}��}�a�y�
Ӈ�<a����O�Lb��%oǐԈ�2��0\
�B�r�g��K�9X��<��l��`Vw�{��`��تm$�E�+%��b��T����T�c��	Y��*؟#��ْ�?ޗz5
��ϛηu��lߵ���p���S�R��h����~��� �5� �΁�O�]����CY�m��x��8�C�8��f��\.��"tJ���g�A�\��F���z�$=�4ie�~�MNN�+jD,��f�s�,�����Ĳ��bj��^ޝQ_$?³ k���IS�N���DE�x��.�6
T^RtuOQ%*Z%G��\�+��Pq�i�"G���d��.^��[^�˖+XQD�uJ7�Gb��lFV���t&���nxi+��۹����0KR��a��J����~��7�m�*d�ѥ��G�~�	��W0B�XoN=��iS���Wn�x�����{�Զzc�d�gI�՝��U����FP O,��һ���F<�c��J|�_"8(���YY����I�`����]�"�1R
Ҧ�P�@�k���<n��S�M�:�fyc�hT�ͪ��y4^+[��,y�ȯ3XgzH8�3Uf+p�z�kR�2L��I�|��M@ȟ,O�gĺ�����Ĉ���j�;��=,eF������XB��rb�h��Ƒ��s�a���ý2�޼���e���t�k���s=i���9T��� M3�n�\Y�^�]d��l ߍ��B�srθag��h.0�n��lwV�_���%�r�vuK���z�`r�����s�ME'�����Z"k��ʂ����Dݖ.�+t8)btiR�C�턗�hUXi�~�3=�j���o=���F!j�����ۇ�u����P��_y� E��H7��f��z�9��-�2�I�:�Fw!�`�3v� �_q#�`?�/��f��X��V�Das�3u�d��J�'M�Z���DJ�����z� s��En��z��1�}���pQ���C@������-f�
�4�}bϿ�X�VYM%������P��7�b�����w�-���i֫��Ul~Cح���kPL0<\��p�'���V�XA��3'q��k$���밚��S�%����������m-�6�~�C����C׺z�+VF�6:����q2TN�y�o˚u���>���u�"���E(�(�;��m�M�-�l-N�욇�;Q�ݶ���N��8חp��P��3��Q�A�ߴ`����݉�ղ�i'�y�]����>�l�T���D�2�VUʊ�:�?+A8������_����l��ʥ��oJ���a��'8O�J6��pwN� �dŃ(��˸�\�������
�Zq�z�.s4��ab42Tփa���c�.�9h�ٝ,�I\'	��^=a�2���~�"-N�P=ӗww�}�[#d��*x�ɅZhSVl6cS�U��*q��(�� ��� ���g�/
�DAG�#�w6IϷ���
c~�{fv�ߏ\"!�=!U{�W��v���jQE}��V�(�#� ؠ�8�l�q�����R\/�.1`Zbt(��D2��[��3O����/�|�e���i�*�����d�ӏ���A*��W���f�>J�Ӣ�	�_n�퐳7@O!3�]eD=� I����#��'q��efQ-�ט���J2�I[F�Ν�����u�c#k��<}|��kx�c&@���;� (�nZq��#����^��Ѻ{�v���=A��ΪX�4z��]��̮�{��Ɋ꫒�S+}�F�t�Fkbϼ�E׈(�t�@*�Z�����>�Q:�[���^���y"~��cJ����=��S_����ݮ$*		�B�˾�l#kBd���-{�${e��d��"{vc����1v�S�������s�u��:�=������X�C��C�U�@�Ild���� �t�D�R��S��Q�\�τЌ�Sl4x��N}���9U������_ڹ%R�!��~�a ��?�믬#�6'�oL��
*!�=��w~���k~ZS&zc�!Y뜗������a�&?$��G�ͭE���a�,���
A5�"�Ж˵~w�h����׬gx0}�J������ݭ)+?o�TA)�q��U��}p����A�4F�������`�=R]�te�4��R�]r䴁��y峥���U$5E95�n1f�[e�El�?֫���д)g}�͖�}g�'b�W`��K�З�b!��43JR5H�۱��
��q5�8t�TC�+q8�`�eQY�[�:&)�9P2]�X��<t 5w��ƿ�s/��f��)��;�5�n�h��t @���mȩ]�Ɲ6
�m��i�>y|�(rJ���u�I�d\:v�r���Yv�x�vYG���«�
��] ^?�Y�u����]F��v_>�(z5�Y��ݲ�-N�y�fh௛����,��e���\k�@�!{@ۓ� ��u��I������]���a7�VE��@�"��Id٧	�s��Va���K�bz H���mߥѨ�?��Y6�{z�;���0[s��� 6Z��Z���21�y��B���iV�e"� Ǩo��������]�Ыs�bu"�ܿ
J�^�� �04g���7v_k�#m�̦��k��ig1(Ԉ��i��NI.n��d�/f]�ܟ� 9g�eCt>�x��!墿��kX��m��&AE�9T�BW�D��HF)����f�x�{�hzNo�k{ a��0o�Z�(ʵͳ��a�8q)�l^�J�3-���[�,AkLf�s�o����Ķ��v�B�i�qg?�����$%*ϑ���%��HF����t��	)��Eco�b��.�K%E�c�|d7#����l;N������\\@�_���惽|?;��f�����0�R��-�|g����\fnxxʠ�2��pJY��1��ƙ�H��P��w�++@��%1���uS~����Z3Ɩ0D_ӓZEy̡�x�޾��(�}4̋�3M%�%#�6�왷6��ҘS�
/� ��,���� ��!�D���U8=W0eNDz
��~��ZG�b���/�р	k�Ը���W���'/_�Ř�y � ��:��*S����d4�+!���,{6�/�:x�-����<R�����Ա{:�p@�3U�c_���/r��O�D�q����#��F��;��x8���q-V?�j�"Y�.l!{7�B׍(.�,O|����ǎ���i55g�J�Ƒi��-
Y`B�+9���#��T{�8��� ��/�^�p�- ܞ<\)u,/�;ݙ�L5����??�y�<�Pɻ�|IC���B4����&WZ�D@_���Hٓ2�B2L-�h������N�u]ij
��)&{y��4���Z?/��y��t*ʸ3�yܗ�k5���v����� 4�h��3��o_d�QgL��n�ݰ2HZ��B{fn���Z5�VE�Hq��3 m��
O��mЗ�W��)Fu�5�����`�� .�/z�Ӂ��Ys譺*F��v6��H���g$"f����RI����(K�OΌݨu�]�����j�
��;��\����F�	�k���J� t��kP�u��ñ�Y);�@�'��J�G���Mo�v�z�~3��-׵g�}9���)��3],��ވ���@F*~C�ʏ���2n��9�n@;z�� ��A6+�۳'j�X�\�&�:x�Zpc!��FOP B�x1Z�ؔ�%S�"�7���wb�ˁ�$��ߏ����/�\����[�{�.�\�,f#�K.���w��B`3�����	s�����W�*�E`�ޜeϪɆK�f�F{�B��/H�w�&�<�n�o�<Y�9�~tT9	�5�)=b|���ߠ��w�H�Id���e}-����|���0[qΕ�֡���t ��J���$ꏕ]U�?��	�Ʉc��)y�ys�T��eo�B� �{�'c��:��Em��^
�M��S�-v��a���v�ǝׂ�}��n�aа���=<���I��npf�Ǒ?t[(���6�Q@��9�XC��-�R3�����g�r;����Vv~��"^�wcfm�S�X?)Nf�]r6�ҞLk��l���hbto:/eYZ�9�r`��זP%WXX�#Ɩ�F'Nh��ٝ��G{�A�j�c��_�͟�&��w�Vo�C���a}���N������"�#�ձgSvZr>À���U]ʽ�ï;�fǗJd��8#��'�ƿ����Ӹc'��8*���a�(����k]0iJD��@F�w˷�ձ݁O��+3�c{P���U0�4��J�B�R�j��A��.��p���E�}5 �Ž-�K�΁���;��&͔��Ə;2]���E%������a	{p"��r�	��-[c�o�o�ىI;e�ٕX�խE�l�>'�����Yr#�fA1�UU���pZ~�3 ��.��-�	��m T����g�P)�݀��i�1�_I-)T*����(�ߐ�f�wj}���	)�0�G��hC��/�C�����vt���C6�F5<�PĞ��?v��3�y;�⼕<
��R���g2̒�<Bn��H�=�X/�2{��TK�98ٔe��W
NN-G9^����ϟ�ZV;���(e-�~��J�+�t0�t�ӛ�Pr��n`&�Yc.�ҽ���QE�3���ˏ2;b�W�1`���&��<?��tx�y70)հ������N�,����lb̻ZK���ՠ\,:�9	9��pPD�i�c3��2��jM��##����ٰ����U�C�n|�ErWS�ٶ�����j���4�+:y R���'��lCK",��\?���mg�'l��3a�ЬXhK��q�5��f4��I�m�����p��7"OzW�Oy��>�-%�uc�{�E�t%ҏU�k�I�=	�sŝ�?>HT{�
�o��\��2���F��[YZ�Y�N�8S�7o���`�~|���8ǸNV?�oXz�WK�� ?�R_Hp��Ċ��3�JԂ+�Q��ڻ��}�������#�9t�X7���<��W7fn8|�3p��f>(t���
��9��?M�O�����6ۡ�FO�$�-w�C��(~5叹r����C�Բ��ٖ��0��V�!c�5Ln9�ь�&~��E�K���9�KP��Wϫ�±�03�:\գ���8l�R*UpUG�0s<��|
��v%�D�;���!D�R���[&���E?h�[\��?�yS��˭�Be��1�n��A���H٫F�4�����a���y�[���%���9����"	S�X���I�)�J��S��K�)��_��g����?u�9,�Qb�s�ǒ�%�*k�x�D��6�ٸ�����z���~2�����w� �9d.mS-�"���{b�Vu�����34a����&,ǂ)Ѐ���?�k57��?	�]1Xs<t�q�rϊݟ���/��x�6��h�;���Mm��(��>+;���r��KNN3C9�)��'�*�
lF�I�!�>����Q2qeUV��#V��+`�F�_���
���]��3w�(��|��������sNנ���l]��{d��i�BI�+w!E<:%=l��h+ROy ��\W�B�2��#��"�m��q����=#y0yEp,2ܽ�+�b�'~�.{&3�w�N�3��D���Ū����,ͣ�r�y�
'<�"����?�$�_b:�_s�q||?�C�+�yGg0�{r�.�_G��Ơk����~E���}��S^��L��i���ɾ_�\}U����p��n,�o�+^x/����ahJ�b3���F��"`������8�q�
���9��xi�PD'J��q�P$�<���FMC����"���S,��)s��Qr&���H�yx8'p�C�\"��g j\���<RH*�������!J/*���4�e���dk�ϙ;+R��H~5Ho��������:ʯ��f'�"cu$͊�w����L�G�n����#�y�5.:�>�@��:�ur94mo�W98#�'hx�M�v��v����N.,�'�7g���,�8�m$��=ợ��^ U�eO�H���z��h?��XG��2ㅘX�01���߻ocC(/�A^�X�\X��=#�?�w���(u�>{�Q̬?fٳ���A�?���>���Q7m�p)�x�!%��G
��B�SZ:������W���������4��Yg��ϫ6��ƛF׈^�p��
[ :��EG�J��\Ad�U8�~��m�ChA��-=�]�@��=zzҒ4C��̕t�M2��0����" ����_:g�,x���3�����9;�i�޳��Sˊ��;� ���q�P�q�g]b�������k��	�L�!vCp��Q���c Y�ghז�i�D8Io��V��ܴF�����j#�g̳>���q'����:9��A㟽�\f$`�>��I���NI���'l�pe<1Eh�^�[�o�x�.����침Z�!ĕbc�S湀�G�=���
臡�1����6Ww�{\�v��>���ʂ�=a�CI_W�ʽi}@�m�l�9��e�ު��W/��~Vu������t�(�.�5n�pj��[w.�}(8�u	�gɓ�r�������TZ�x�)>&H~pc��fV����`/�}Yw�k�w�r����u0�ޡ��\A0��f�.�]��/���6yS����-E�^{I�FƬoO���Ԡ��K=��hT,�~&�ץ��U߅,�+�a�m���a�z�+�eݩ��L<���s�+���j(�HZ�C�@H�Dޜ����oq������C���W�F��� �ާ��V�%][q�Y�"f��;�&F�Qy�ָn?,��� ���E6Й�6uK��)��?��-��aS����!G�D"s�����g;f!5�v�Q/�J���[���M�Y���ȻZ����J��&3R7}�B�	08�>�;m(�o0�I2�!}�{VB����|��LS�@_Űӯ�U��f#`�Ͼ���>�D��{�S��ȃ��}�,Š:�y�q�$��(����I����4���_�Ԋ�$�fӍG��_t])��*h���w�G'�z����� �)��A�R�#�g�	��naiل2t[ܪ�_Zq8�g+�_U���Ea�K�g{Tm����[g�W�;]������Yӯ���ͅ�������3T��R����T��K� BL?�$�V�K�G���FP/7�MFא�#���c��bU���?\�|��H��1_l�'��������lxg0�lӟ��l�2��+Kq,�D�X��w�u1���-Ǿ\�)���������X�5�]�AW~È��ݍ�R?]p��7�S��Zi���,UդD��NX����{"�\�t\pv-6�μ�>��n�����`6K���D��^i�9�F�y_����=j��k���_��m�������7Z/)̨�M>	�C��K��M�0A]m�<b�2|B4�!����ex]Mzn�>>c]���ah�5�0 �t��Gأ �Pa���P�3J =�%�����_-�׵Yy�W�A X+���!ho�T�Npʌ�㝰!�vL �o�+�ĥ�1P��f��� 9Y��ƹ��ȅC�O%�a|7�"�Z��Q��]D���桅��~E�tb;���|�9.k�̿�ч�ņ���~_D=��d}���a[M�L�0�z6����t���̭�������o	�p�sm����7���K��g�&MC�Kt��!+T��	jJc��T3%n~,��k�^��g!ؔ�s�T�;h�Q5w��ÿs���[sս�˾��/��Rz<��2���\�8{�nL�>��_d�U�y}t�GC�B!��k��̭�J�K�}��a�IoʦY�_��=� �������ͫ�2�U����V8
W�N���%p~>m��A���~��?#�^|7�+J�wJ��U��mBU���u.甄Q��h)3�v8ݽ����מ�UM
���}�N�䦔C�Ҝ0?�n	V�	��S�����~��Y�Тf�"�=c��S��V���a$�)��R�gc��|��w����C�k)Y�#γJW_S&�k%Y^�
)1���B��*� ����f
}��r�r���F֚�z�<,�d���oؗ�D�zV3���L��&���k��v���HBYiU�_w�(�aWt~����ҽ����ڋ	���+�FJ2�^	r3:K8f�4{BPջ��[9&���i3l%�Q���?��/���C�2;C<=�Ș�4pD�(��=�����tgW�#�����W-W�t[C�Ĭ���K�}G��F�[��>̢T��K��EĊ��2��AE����g�e�2Ӄ7^4~�_��F%�o��r�/(�q���hU��E�%ǭ� ��Gz�5��O����@�f�'���⥙"Lȯ�
b�qЂ���Sd#>�:d�B'�&�M^"h�=x�5�7�v��9C�D�L�å¦�Z��c��V��m(���|����Ao����^�|�\��(M���s�ǆ�,�����#\�{k��<�IQ��$��q��QQ��9F�}k�N@?�V������댢��Į��|IP��^��IO�u�&Iϐ����z�Vr��B� $�����W���M�^[$��vB�{1\g�?g��9�dp\��q
�3K�Dx%�%2������:4h�^����"9':"̄���k���M�Q�q�Oemv�"�&e�2p����l���We�5t�'(s��~��y�-��H�z��M��,�!'m���u��2ơ�n�R��J3���ԥ+��ʃv>�7+���n�;;LE�\*��ʮ�O����6�Rj~ї���ݗDf�܍�Q�&�4��^p�r�i�æW��'�w�7?>_*J�"O{�1�6��%�� 9AhF>W�QAv;O5�yQ}��ж\��/.gVʕ���"�������}��`$�\W�N[z�K�4Z�L���qHy�#�7A���{��ߎŬ�?Ԟ䉌o���NT�*��Yr��]C��$�ҏ�0NH�S=�#y�~>!��/���3(�Я2q�y0��p
ݶ��pw��^}�����Q0�s%�{	V>j��o���[E9o�Ы:��
��a��� /��4�������]Ik�s7�$����z����CG?Ƀ����v�V,�|X���5no7���D�a�im�ͪZ�����o|�wQ�!Y��dB��Y��~,'��#9���!���O9�#��㖽�$>�^��vП�x��h�8�$�VD���&j�y�������Ҟ[�|��٘Ģ:�Q�Ǖ��f�*������q�v�S��"��m%2�
M�b,%*�9�x�,_�� �G�����܄�xE%�3�Z=��N0��:�vCz��ts��jA0bm_�y.�u�Y]�\���7]����A�����CX��X�J����Џȉ4m��_Q��{iu�ye�;�'�~�v���{�K9�{?y��1?�/�t~S�:4�ƴ�d��q#A�����t�-
gsv/�Y���,�-{�DW��=M��YV ��:W�*䦻g����oP�q��M~��3t��-{�����طA����&����Ԭ�����?w{��]��s��Ikq��-,�o��\�Dw�Ԍ�E|��H���c��~�[�@�G�綢(�T?s�A@(�0�wgX����Aߖ�=��&u{y�2>N��{���ڮx�ǃ=�AV��lE���Zx��!_ӫ�}~�@�٥�N�W��	4�<7��5��d���4«�uo�0�-w�G`e}:��&��]�QM�C��y���㰙y��0�1ɑ�ɽ�ݩ��"�L'�?^�Hg���G����3`�&S���m�ؤ��L>��~U��_Z �n]	:\�i�s�|�HZ&'���[wQ�~^�޼Y��i��������ߎ��؆��VǾ��s<�a���w;I9tm�k�@�siRN��ۻ
�U<Y9����Bp���*���*�y���q��0��z{'��z�����E�T�����H(�Ƿ�u��}��~Z�F�`s�Nٳ/��U��=*�,�Ӓ�҄��~<��WL�G�.X"���l}W�>Ǩ%s�!�7��f���iP�k�?��x��������.[@i��z��6���H�]���<��,�x�y�����u��k��@l�E�&���q�oZ��c�uSW��X�+�Qg�`����\��3�L����j�vS<��7��>0�d��1�y�v>�,�<���v֘�^���;1q~\I����,5z��+t��K��
V�ۙL��XB�s��I�]�4��I}Y�r?���_������%�2�y��?Q�Od�=�v�K��)[�濵���I��g5�֐.X��4)�[(y㻭T(��=(}�%���Ÿ"㯏�ܩ;7�r/���)�V�2��	"�ju�}f`G^/�|��+c{�G:�,��`��G&�_�[QWǯ��}��;:�
s�{�J�S��3��s��Zm�J��mQ��%'�_VX�;���@��'��)��eF��ї<vy��tK��Q+9�xq�E��j#��]9ރ2\�J��뵛]8'�wL� ��F?ux95נue�Ǽ���e����f��/��lX���(g����@�f�J|�(K��q]ۤ���qe��3ZE�����ݰ��]����^\�Z4lW�8�赏�Uf��o���0e���j��E�ޠ��m@Ő�%�ǀ�Ti�:7���_�c��A��!�f�˩ιoSV�K#��{[��UMk�L���"������Ǚ�_����SP߾�Ln���Ȑ�7]���"�Y���s�������\y�f�f�g�]|�����������'�^�N򎷕���-|F)�i6��Zy�����'�^�q__q�T��(�����>�=� L(�^�O���j�(m˕gJ@+��
aӓ)�)q��^4���z�i5�L,����=���AA�$��b�u�#��e+�G�2h⢆���P�I��aW̺��a<�͙3����_E�q���7��Gy'2F%n����?�>��e>���r�N�6�	�E6���TC��
��ۡL����z�ۥ@�\	���?/�д%�-��8�3�o)Q�sB�:��KWFؤ�t�UL v~��H�A�?\�0�+��%W��>�;���Nh��[�`O�Q����..t��9x���]��
^|/Z�K�1�c;?��̙�5{�-�{f)<�V��Fw�t���f�O�e���WW~�\G�D杭���tT��|��v{��1v�3����2<��PØK�	V�!�z9�,�����t��7L:큾���g�K�� �� 4Ӷ�v�.���_r$�b�r���|>�)4�ݕ��;�Zv7���-=������F�vhUĻ��-�Q��>�f
3���TT�%g&��/��R�V�[Km2����%�v��&�l�a}_��n0�H��c�!�y��]M��.�`۴"%h�T��H���a��׵Kqo���A��Ӑe��7r�)������0׽�&�m������m��I��l+�����Փ�LSY�� �<�9�{�h�����y$n��z
�TOv��ݶ;�N�J׺�D�Q4:�U��x5�������P�%���o�vz���q���@����zl��!M�/g>��d��v�BAI�c*@s�����/��E�EBS��#eD�#c�K8����6�w�����*����i��?��������,��7Gԕ�O(%��~:���kx)KS��맼�:6��!�1 N%���ZS�#%P��EY��t��Ƕ0�aOP�kq�͹-r��\>�����5��]TRo̻-->f���~����x�}�U� �L�}�΅W�9� �i��7V:ٓ�Z�8;~�3�������N�@��fNTP���:���AȄ��fI��,�D�i/z�F
u�=b�N���TJ��)���޽���C+�C ��˵���~����3
��#�ߢ���}_f�v��w|A��m�E��7� ~6����o'��L��0i}K羪Îe3 jr(����+�|����N"�1
�F���N�����{~����Y������&F:��r��{�H�=�,&�l4�D�Ɓ!uE9;Lx6I��u��΅��w独?[ցe���
�nǶ��g>��%�;���c�����"**� ��#=��y���AT�sY���-ᕗ4+���z��J4!ԧ9!�u�j
���nwا��Z�U�����_l���'��إ9S�񷲔�R��sρ*e�s��b�k��wтb�k힖�q�kjr�9�4�}�E�E������(7�O��x�?��?Sd���P�4��Цx웴?&�{{�x��c��B(�a�	+<�Jc����.���g�k��
2����ڞ��9�nd]��~*�j�5:���vz-��~m��2�N
����\X���1��k����b���Zmy�ٴ��UX��R�k��iRݍc��JW��Hߡ�9�cK,���o�������r��倯�_�ViY�>Ú��Ѹ�3�;���I�"�/��[KYi�X��4��[��7�*�װ��vh�b}����`��A�2���u���y�����ՑY���;o���_{_5T%]��a��"����Ջ��|��
�	N�W߫	��� 'Xd}?W��r�4����s�� ov�d:�{�Yej�J5?3��cMp�Jݎ��t��B�$�N����b���J�Ӛ��?��2��tR�/kϪD:�����p�).���4՟k(taSһ��)R�ODe�-���9�������}��0M�D�d��؆��i�ah�ff�gGŧ��n���{W	ފ��~j�ެ1�x9��RM�>\���M�z(F'�}X«Xi��E�%P=�?&>SlYw� H�I�j[x��Ȝ�̕ꦱo�q��9���65��QCB*�����T���]2�����i����zG�
��>�
��0�C�]Q�#�r��v!��d(F�w��X�uE�ue�S�j�~	wn�:���FO��epJ�E��q(�b��� ~���#�](V�̟0u����`�?���m����Ԕ��`Q��A>�M��3	�E���Yr#�n-B5̸���)pe|x��h��Ҥ(H��ht�|�;C��Ea����4�P���P��PЭ�洵��K���6T�Q�j��-���J'M's�w%����n�hJ���џ:���j��eu1y��)h�2��M�U�E>��4��B�z|����{��vG����N=;Ct����@͇k?8�I����x/,q��i�9<���L�	/���~��*���TvE�T����U>��2�P��2j�aM�4>"���
w�YÞ��!�M�Z��"��|��[me|�&�[᣻=��/�M��ݣkh8z-.Ӎћ��?��}l�f�}Y��x�}2�B�Y|�T��Y�W�g1�"�89�t�2<;�+�u�^�`��9�1"LP�V�*�gO�����I����𷞎{E�R����v�ˡe�k������s�mY^n`~�V$����bC����ͬ��6��dM��H��������������r��-6z>M#��Qr��F�Qd������J�g�Ҧ��s�K��^�Ұ��J�<s�h�^R�o$�,���ө����4�k��a�*�����[�b��~���b�˟g��*�`X������� 󏒂Ф�^�w�z&���c�Q�LG��$��{Ĵ�S��z@'hf	�[{4,�	C96��3MO��vQ�Bs� l쬿F�0w�lH`�4D�4�㏉F��Q%�G��ٳ$<6�Eq��ХtPmL�����r�V�Pd��N�.�¤'eVhx]�:�oVBC
�l�2�y�+&�g{o��tv_�jsv0֊N�B���$Hl�t��jē��U.rZP-iv٣'2V8f-$�+�����FQ�f�9��jDA�f$����T�w�<�*�X��9��9E~��J\O���J!�����/�2u�Q������Ӳ���}jD)�������|+�+����Y j@B��	���YT�ݸ��6��tI���hB]��s�#N�V�&S+�~��*�!af����q=Hk\R�Յ3�������'�љ�� �/ݮ��;�ׇ�����AK1�f�R�	Ǒ�WO�E
��7OE1�v��&<�{�^����6�'GN+�0��t�^����[~+Eփ��K��~��:�����D[y���j�d~�Q88���i�=6����;i{*�����A����Pm�N����U���IJ�6��*��+S�g�#)ώR���{�(�(�.�@��eڴ�3��hJ4���l��V��du��%|��薱��Db� �������C���_BOm�?�x\�v��"ᶓq��όM������E��u�����cX������[��M�8��l9Oo��Hi���T��D�)��	&�
p�h}E]�j��F���/bld�]̵T���;��%Xú���N��6���`vû6D�Z�ⶵ#�&r�/��V�D���	�5cSg�n�*����+J�J�wQ����q6В��{�]�ö���5]��fl�/�]J���5��p��i3��m���~iMk��s+��C�ƪW���\�>{�i�V{t�U+H���<
p'c�	N�}��0[�;���H��~�"6& �
����0��<e�< Fbu5w)����[w���
����uB�ic@��,�|�!��5��uJo��t�J�fUD�ܮ[�b�Z��MCB�٧�e[͕w_?��l��p�f9��pr�70gi�:�[�<\䏦��s[�	 s�}$�������{������J��^(����~��Z�R���o*}�V:S�H�7}��-�Y����>>���A@���y �r���~)�r�{L�IG����L����K�+9;��AT��CkWw#��f���\�]	]�J�n�c\���}6�{aȩ�`����!��;b�T����@I	�3LW&�ϰ,��w4��٩1����������i�s��e���a����|S3(��Y"��*�n+�틭-���N&��J�ŝ���s�����Jۺ�:�YnK:Y��;+k2Yx#V}�'J*n[��t(���:��^lK�cK���S�9ٮ�f��(�}Sw�
t��k���M��Y8�㧠n�5�������g��[Y�!�뱜���b;e;d�#h�_]�9�mm��4��c�QS�� ��ݕ�����)�r	��6uu�!o5M��ޘ+țӷl�-��"�8?c�3s�:�M�H���ﻣI��c�e��A����~I�����_�Vg�`����]�3뮴���f�r�
%�0;���Ub�{cz�R��3�L���P�\� .n�	e^��& ���������o�ۆ�س�c�y�@1�UY�����������n���Ŵrs2����_���'�����Q#�p������f�[)(�sͩE�S^��&�����Ҡ���l$�B
��/����s!��V_W ���������bk�M��:���6
g�.�`��#���8����n,��x�&�{��/�
  �����#6�m"�*e�"9�m��O�|o�l��P�^�)�k���D�$R���)r�[�I,-��'�מ2xw����j�A^�}N-�Qa�=P�0�t	�d��������g0F��c��c�*�5M|*?����5w!Ř���w��x��{Q�q��K�Na���}����k���V����}�𰬛�zU؜^7Ve����O�ͼ���%�C�$���{}���#��&�;+^y2�xtb"ywW9�v��O��O��!{����	��~ڬ�/���/�����m���9�Ic����Х{���S�=�����Te��V��V�λ:��C[:�b%f#`�7��a%��Z	����ѹ�D<Y�(Y�
��M���; 9w�7C|#�{�-R������[ڴ��0�b;�偬ρ�
eN�h8	M�g��OGj}X���j��L^Ϭ��rK�g,s�p���w$7m��v	���J�_u��coD	5���O�d>��Q�S汹�>;&���I����}͝��*b9sɀ�}��~��$��F��^Z�Z�lE��X�64��)!�%5����+Qڏ����O����~w�L��=0��k��Y�yD܀�;5��-���
��cJ�j3(��o��ɐ���wk�Ȃ|!1��l_g�ϧ����}�T�rgF�4��lVS/qcg���+���X7�J�υ��g�օ>~�-%i�Ҳ�kϾ��~%B��!�	�B�����F�JrQ�'��7ɸ������tB������i)'��}���X�=�L����j��V���: �Q�I�5�q�{�'��������*���X�+k��ɬ��y�)�T�# :݌�� _���I ��Yͦ���>�&:Gw����_�k���6J :rm�����,+zo�S��.h���!�ԛ��
ƚo0�bg�^i�)�� 5�k�0�S���5\������b�������rcQּ����1=i� ��m�����n����-)?�q�4��F��'AuJ/�!�f�|R���o�X��7�m��^�J8��~��7z�_�Q�0i��?���[G%��j��z�Z�r=���z)�f�s������4��q1"$�,�5	o�VEN1dO�����@4}�e|��~�q�4���x�,.�>��J�K~[co�P��b%~1����� _^�u44�?�=ǹ���_��0zb��go�a����/|���Z?�{Y� f�^Ċנ(���s��Eύ�O���E�=EZ󩏗�J�Y��!�	Q)�']e�8�N�!w�^X��i��u��:V�S�F�G��3O�c��C�vJT�����Ll��۝�े�5���j>r���Hw;y�+��/��8�-\��E�CWYi7�#`^��(�8�%��}��{�a�n�q�X�7�����'���ؓ����dU?�ӓ=��y1�.�j~�^��%xu�Çz|{�D[x�P���k��x�nNڶ��[)����1��P�z1���6B_w��!��[N����T<V�ќ���X�G��Ɗؚ6y$�c@�����wm��ɦ�O_����=�.F��N�y�g!�{�L��<!�O�[��)~vn"{�x�{��������'���Z�O/��F���^�1ђbW��1�I��غ�x}��d���~]8�q�ܩ��;�aiz��ZY���urr���-A�-X]���Ig�Oz>�J�e�8�q͛"���d,�!CZ��1��Y����|�S��Ϋ
���YV��~�^�pJ.ӿ��%�����)8�Y�Sa�[<�"y@�c�QC��7b��	�qW;q��i5�س�W��� ���u*P^N`��s�Fs�6�>#\w-v�Tڂ3���z�:!�}���f&<4�s�G�c',<=��f�v�~���J���Z��$�]�����s�����l,�zH��b^\fP��Z�q8l��x"ۖu�ɯ�oU(W�bf�:H�T,��e&c�n�uJ�ɢ�x��
܉�w�K�<�\�D,���Mdٲ�r�� C���� ��s?7ݚ�X,����]�*����
�c��;��;M���!j�u�����)Ǟ������ڶAI�qGp�Or�<4�����e�Q�R��v�e]���WG�=�����琑�o2����mٓ/\��A4��D-��y��w�.�UuuXt��K�Y_��ɇ;I��u|���?Yu�z�X4�i��n�PN-�^iw���!�c���,R�2���،��a+�%���c��^���1e��Ѷ�eGN<}��br��Z����\��;E�{�ъ$ӕG���"�S��E�-������G,����17ç`�NS0wi�W�429g51Qw���϶7�zRf�� ����0��v�P/�ލP��h�"^z�Izd%`�r'i5K��~p(�����PN�9���ޅǓ�m�*����阬�t�%] գhݘX���:�������󫊄 �ؽ��س߿5����D�:�4��Ze*��]���8�c�}]G^���J��x�B�uJP<��/4e�¦S�@!� �Y������G:�
�ou��3hE2�}cj��)j��sd�ֶ;�2YB�Bh��;)�l�qv���{(���VD���q%��oV"hh�!���[P7B����@��UP^[�G>�eJ-��11�#�!PKM^:�?�d��tT�!#`���/�r����7r����e��p�ɾ�� k]��Lj�XN����c�8�d>P��4�Ε��܋{���bc�}�J�u%������{?~<Q�?��$�sq�rs��>6�n�V�~9vJ�y��/MD�Yt���*��nz��R\�*JZ���L��9O����x�ء Ld:����	z$y.,�	\x	K�RB�$\lY�ɪ֊`�:j�L9>b�6�&I��� � fe��U YuV���"7a��܁YJ-�X��6����['kdc��q��_��CW:��7�q>)݂�3,a��m"`A5'QGg ��U����E+�=�^CD��%� B�FF�FM� Q� �D1�(�{�2�����{&����χ�����{��^k����&���̝����D�wJ�*��G=��ƚ�)%y�L����h�&��MKV�I0�acƻ�Ԧ��~P4H�Px�Iww+�(QViM��u�O�[�ަ���;����&�<�ehz�Z���}|�@���J������c
>�b8�Vl�&̜ɚ�5/����a���à���f9�ώ���7E���?�k�*�xF���X|�:J�����ן�*�~ndFt�o�u�<H�}��nNn��U�w��5*F9�=z��z���50W��lJJ�4���C۝�M�m������^�� )�M�~�����\�ۦ1�UZu���N
s4$CgC9�3��M�虼�ɔL�#�o#$�{.�kBwCĠJ��^d�z�h/`x�y��5&�3Z�Ƴ�g��^:�\�y�Si��81�t�����t�h��.�,ވ�dy~��/W���@�Bq�F��E�6��/2>�͏�k����L��ZQ�4���@u���D^-�M�;�M�VՑ9x4S��7���
��t��ϽX��;jRQ���~k�S@~��8����SqIVzc[z��S�p���D���I�wΫ���R2z�e"�N��w���U����9�	U<�u�?�j�չ?� �X�9�3��%�	"U/���E_tQ��,R�U�^�'K��nI�k�����s��7Mk�ctn����`�8%������*0���%G]��;�U?&;+��&H���^�(��!b�{:���)�#�h�G���a�D�(kn�{����<>:����g��`q�4X��� �i�}@��k�
]_�PRK�u2�����s���&�e�u{�)�V�'}�mQa���C�*�(��:��f4`T&�A�7����!���)�s}�)u������p�䵶�';���0Z�a
��tV-S�K@�k�;�_�d���%4�"��[sv,+-k���ԭ��8��W�r��ь��H��v�aޚ^��#�-=�D��§�)&�ˌ�f�I��WQ�I��ɚ��h�~X�Ov����N7%�o��������??�������E�*�Y�ﯦ!�z�V��^���P��cY�@7M�(���j6���H�@|��u��2ì'��\
��Ƶ�o�02��f�$�T��ƶ����}_�[Q�x���~���N�᳓�O�;����i�PT��UZdZ�΀I�|���(ngH�z`� �>�
�M@�%`\�T�Ս�>
�W{��2B����^��7ފ�i�n�ɚ}�}Hm���}�=c�Hm6z�)�>��@���V�!j���)媊�Ŏ%�J��S�V�P� �сTm������i�s�ɭDթ2	�^����IHME����³�%�dH��gD���y+��V��*�&W��kϛ��yT��9�~X�4P����6{��fL�7��t�m�%6�95�@y[�^
�:L��/�C�����#s:�S�HN@�����B��yƪ52(��xh�t��7����Ҧ�|������>�`�{q�4�gX�"*L�|��@�6e��_�aѣ�T�T��'��x�7!��q6�ǡGv]i�XO���K}�c�V�{W�A�%z��[���o�JK��.@����ʱl ��R��=mz.���`}�k�*�nS�W!=f1����7�cv�5�)	r�V��/��<5�M�9R!�9�h���h����5po����8N��#�bZ�o`.�Ǘ���}襱6g���Pj�ց�>���	���;����<����N{{���T&~(ʫ�ѯ,2C�lpF���49�����Q,�X��Q֎	ǩ�4��^�K�=��
�W�h�*p�ϛz�����|i�M#�n�.F0����i��������X�<ӧ�~g,���O�)ƍ�m�iz����H?Gf���ɲR��j�ö�ߢ�?��ϙQ9r�n���:n�Z�;ëN�v�m��}x������_�F�ΰ��E9�䢤�~�l�ʺ]�?�|��ޜ:�c���7������1[�TH�0�7}4w�3ǆm���H���/v�,�V��v
�?��@�5��l>���\
?/��C�q��ö91F���52��3si�m��xS�Ў/0�����L|�V�x��p=�[��-����u_I�J!��\}�<��20��7o��L�;(*���t����r����m�5��9��Tn�)�<��;���17�������Ֆ�N�(�D�
�,�t�;�Y�^T���/Ɗ^�K_ELw�t7��>�����-����>����P��b�/�o����������r�:�A���bҽI�ߡ�}C��d(4�� ��!⽯��zZM�1��)q�����Y�o��v���+9T��D
{������,MJ��t���9�P�Z�,�bU�q�44U�$@0屇�Ԡʂ߇ r���R�r�{	ɍm �W���g]A��F��@8�l�zolE]�z+��C覎�LR��v1땹��FϻLP��;ݧӛ����P��
c%��YE�=J�zK�˛n�g��yZ����*����V�z��n�<ڈ8R��p?P�85V��uɦ��wBo������[O��_�X�4�`_��Kr�:��Ɵ�1����ӭ�ow��P~���in�+cX~���v��\&�͆, MwX�Z���Zy>/��e	$M�����:��N�; 3��)V��A�?N��WGM�b����q1{��#���`x7�Ńtf�a@�:O��mh���^Y}��"U��RV��iL.�_��5�S��������-.*Ldk ��;�b_������Y^ߋ�1N��
��ʳ�� �����e��/������<�bkkk��o�E���\��g�~�?�D�*���F9���s�.ƭ̺,pAO]N�,"�IىC��s0!��p�+��X�2�Z�Q˲h8�3�
�����WII��^���j��D��
�D��\4ZR_<�RR�H$J��p�g5]�)���Yh񼟭%]��%��8rw���:�Y�2����o�)j'��o���<6U��ͫ"��/v� =�~�V/�{�&������^�l5�~b�ؾiȟ���M=�w2�v-Z��*?��$��W�'om��e.H�N�]Ww�J�,ڣ���<�^���#�7E|�mME;����"������/��°o'VW����y��nJ^��̶]�i���X����\� ��e�'�K5��g�=V�5���J����������c	%��Q�e%_Ѐ��[W�P꫚�OR+��F�2�ţ2�j��l����T���K\��E'��)I��Z����T-h���gu[n^=�c�U�G��祺\�����PR�s��E�ξklxPl��鷽j
"�f�>����w5��B;4���"�z��w�v�a���Gd,�\�f*��B�'J[ge����S�^����^=SG�$����������Hw�D��r�
^����*�B�����qz�=�'us30! �ς������v�Jb�N`@�Q9k�9k_pn,�G���~U?�]]eG0(BڥT�a�S*�|?���TI[�X��#��a[��^U*�o�WW]V�������Kb��8c�N_V�B��j\H�Bb4R��c;-zӎ���8��U�Ŝ�,$���O���'oqw�1��z�NI��EM������2�S�F�Ѩ��R�Ţ�ڒ[���s�a�pK��� c�a}f�@@�u��$px�P��Q[�Q�9û����zeff� Ī��1��_���Ω(
d|x�3L���2��O��4I�:q���5���N��6��ym@wOV߽u�	g�1+�C4�:N2#���p�۔�G�aA�C#Vi�F%�����
e3;�9lX����|��`W1rJfPw<� �L�Mbw�3d�:�8w��C1�~ҿ��_cO�\�+��9b@�a�͞�҉��Yв�/��ؖ��td�O��^ת�e��L�0	�I�	�
F��{��C�H�nG����][m'GyݹI����^���ru��}j��_��ѩm�c��w��v�w�^yd�K�f�j�w�sO�Ы����������w>v�\"e�|��7��m�&�����7C+��Ss��~
���� ���������)��$�g���6��GY_p��xr�������퍅���0�b�N����~����3B�K�Sr�D��h+�Y+ �(H�>8�
6I��0E����q��!�!�w�5�σ
W���~��Oд_��?i_�z8<9���!�%�ɏ�s���S��6%A�;ga�zQ���'��NT�ԉ�S�Z�B�E``a����1�Eer�="���7S=8�C�.��ǣ'�t�|��`/֘w�2�3Zi�p�F��"����D�֯.�}Q�X��ۇ���d��f�8�K��򆷐î6��]]Crc�͋���,�pw��K�_S����$�H�J1�qx��С�ņ��I[B��A)�<���#��Ы�Qq�jN�>e���3���Zh�/Bo�֏O.�+V7R��+W���kX���?�:�$��,�u3����Xų����GeS+i�/s�Zc;M[���{��pS�R��"���kSb���eb��|��$:�4o�ݗ���TwTƧn�2ݧ� �3��|�勋�R�,Gv�ܳNJ��5^�Qu����O���˒���ǟ��纎�b���,��%�L��xށR֤��[�iq}���+�U�F�L��Ǟ�z}��١Q��9��x���@�7�ᖋ���R�&��O���+�`���o���{Í�}MlIk7�eo���W���3=�>l��j�R����$���ࠛ.�ݣQ���$=�H��͖qw��$��ҝ�{v��̅O��WYWON��'ҭ(5Ik�;� _�޻ݮ���^��&�N�J94���(�*�֧2����A���g���K�|΋h����R�a�L@ٳF���[꘸�~��!m���e� ��@���_,�@N�g�Y�@ϻJa�	\�<E?\^��Ն��Sٓ��y�H>�{���Kl�g�ύs>�j�h�>4����b��q#L�����!��g}}^=om��G�^�����J���x!��Rx/N�x3薛��?�~�u�q+Κ��&<�p���^2�K�4��`�\��q���;oh����xh��~_��nߏQ�N6x�F]>���d���0TCc!k$1#L���4,n˺��(��7z�i�>�8��_0�x3����o���?ʹ��IՕ*�O
^�5��C^��S�=��Z�g�����,HU��p�%Ds#S��r�i��4e'$J�σ��M=s" ��N���]�����/��n54���Ywj������-~jY�b�G*��k����8&,��7t�Ѱ���U�07m�DH��`ǫW���x����O�c~(�)�)$��#�E=�<�����dny����*��t���W=&�n,��;���m�K��J��]��P�c�FSj��x�Nfq���q�<�PLcԫ.��:T�{���y�阂�}G�f��.ˣ:�uxrb��:�SK��.*����1]�!���Gl�/-�Ɉ����Է���4_=}�x���k��ׇ�������>~ ~ֳ�K�J��pw��|PS�t�7|[%z�%tU���_���Cj��1�۵�Q��*������V��x�"�~�H�^z�T	&b�-�qe�����ۛ�O��︃i8}�>m':lh�Z���Ѫ\��#�7{���_#?6~�i�Y5�|w���?OA�ߍ�ٝ�� �����z�v�Cy#�������d����G�D�hm1*�_'iy���fn%�
����~����RG�����������b��d[pYG�'��"D��̚P��l��r�à5�j�@m
b='�Mњq:�x2�������6N�/Y�d�8�eQL�3m��_J�h�����u�9��1�An�/�"z׆]�ܨdS�b�����+�Y�/'�Z���~�2�3�OFX�%_lÆv�B5j)n��`Q���9��*��C��*����ƹۻ��o��_}�T��w�u����Y =�g1�7&z�k�Y��LԶ�P_�T�\g�cHAګ�����CL����I&. 4�+�-l�	�C����;;]�s[��m�/;\�{LyMV[L�1�х��Ҹ�H@���7*��f���Ύ�^G�-F̠�O�l=��y�CهV<C/�����_@�_��d�M����`�J�F,-`������v���fT,w�k:v�]�z�Yn]}#;�U�A��V���*�罡�R4��`�[]U'����1wLf�y�,�~Sj�d��r�D�	Uv�;�틑�����Ǝ�	���cW�<����!��r;O�v���������ͅ�t_�9�D� ���x:%M`��"�� �鹺13+�LW���VE�I=�R�����tw���M]mގ\��>�g���uI�Pؙo`���.b�� @�F���.(I�C~H9#�����;ث6��k�y��,ZInIu;��F��{w��#O{4��e3�"~�'�6���.;���V���6����C���oGgp����8�v&�y�<sv.��d����h���7��Z�^H�I��i�0�����|�Y��SS��֭��%��D��0go�(�h�mp"n�)C�;��gq��9޲����c`ǵ�3��
��I�Rn����3}��>��>@?TY����a�
�z�v�ŝ�'�� ܲ�r��_�	DY��6A��%ϟ��׹2�3v��qj�}�6����������Y8x
5��D�>0B
	`�����Z��"{��胁B��9�P��󉚜�ҁ�k���MnD��<8���:f���8
.c��^��:߾1�BɡC�H�J{4�=urN������W���4^���:C��3�Ѹ�1音|��,"Me~���ᢛf�?<;�1�LJB�����78��]/�b�\-9���Ͻ=w11/r��ҏBx/[{�_>{�S+ô�=5��VB��=f�g��z�,��ܙ!0P�&���I�
�t�dE�yh� H7��3�WPĄ:�z<�qХY>�'u�I�v1�/. 3���{��r����d�f�%f����n!�Ĵ���y-v���ot�tD%=(^���Q�ݳ����@*K����o�����\(�QjY�Q��V~�t6c3^'��#$Ww�F���7�Mﶴ�Ӭ9Ffgc�Β��$qXD nh�����4v��� �o�b�캊�ץ��L?�)	���Kÿ�|.�߻�h�m}:z�p·�S����}�4C\�q(����w�U�5dV�<�F9kؒ/��il��~Ӈ3J>��m� �E5g?
�K Cw��5d�X%�������2	�����0E��|[-c��Z`�?���1�8�2����u�W�{j/2�[.���ʁIUė�F^�����*�!H�(J���ˮR�>��f���0KO�Ң��D��-��6��=�fKR�0�w�&ˬ�����;M���^sn���Nk���h#F6�o�w��k�rU�鶘F����e5{��Yѿ!�5����>L�Ԍ뵆�s��<J�@)��)���Fe8_�}������������~�f���O�d'�,������Ɲ ����˘�b�˝G?�)�y��_��t�J�nT�s����W�
5��J�7G�:��p\X%ޯʗ�|��v�ˌ\/��="#L@A��������I'B�[j�)�0�x���Mu��(�}fh�dH�����ճ�)���ȝc��b��嗗�2�@r�~�a� nM���8��0w���n����r��9�)GG3�0}��ɏ��.|Q��`Wa�Jm�( ���	7V���h�r���K?�0��侜2���j�HΝ�7��Ư`�h�j��P�0��9AZB���rR�K�䐷*�US�~���|O��/��pU���FT4�9Ŧ�P�BL���5�l�{����ҳ�p]�	��n�ʒ_��N(%j������l�;�?�_>���&��ͽ�nx8.{t���.A��q��m�HdրZ���,9{�yrʐ�"�ɨ��	�L�l�a��-SF	����p��!�㊪o$����7���a�E��NR��,��B~�����;D�> o;N�(�۔� ��k����]�n/�
CkX�.$�]x��U{�Q�_O�y��9���h��0X,�Z5Z������;��U�?����yG�*�,����d���gF�@�VVB���f�ym�g2|�<X"���[�#���D��R�]������&�z�O�z�:��`��Pw�׏�z�?�$�, �����kۓ�ma���0�3��k%�bF�E�(�er�gv[�$u�ۦAy]߫avO	a��m�]ZK�ky����7U�R�1�h�K�UTV��������k�#�C�Gq����5�� lA~��ks@)nsՕb3�p���8����������p�����5��Iw?��0٥#��@洅D�Z��c�����ӈ0�V9���΁�@�ߺZ�\D�=�������1P��MIz��{��'��9�x�tҩa?��ۥa��S�ž+�rʣ����H��S�Tr�f���qP^�3ɏ~qţr��C�\�l��(�3* Ҳ@�Q���t�LXj�;H譟��cc�q`�s��x3�U�m6_o����J>k���RD�Ĭ�|�[m�w�-b2���I�o�-�hg���>�yկ'�TB��%��W�lw[O1{,~��y��\!���� hbݪ�WPJL� ��K�ڀ3Vپ���R�/��6�M���p��<ڀ�g��<�C�����ն�Cnv�%��k& O�khqXY��� <�'{��˓�i��8٧즌2��߼�^�(Ơ����"�o�&���l������Z�\X�BCƸ��3��&VP�-�!���WoU���.3ɅXN�y�M%*ՠ�o<"Aޟ����,]!ȧMQOS5��ȳA5��8q����UUc �����;���e��j���d�	��7�")�Sb��?����֑Z�s?�=P�N�#�2��)5>�������aI���F�Ib�s��t�*Jr��n�!�P���^<���M
N�=����۟�6�4�RBL��Ef�y�Z�x/�o��L��3F*�:5_y�Y�t��A�.�	*�Z�Jo��\Γ�67�'�H;�u�w$@�M)���JP�D�������<Mat�?�_��0^#,�É0mGOC>�n�3�n�W�3��o� T��[Gmjſ�sUʇ�xks7�8/Ԧ�U�����I����������<'%���_�I届ij���}�t(��Փ�)}��e��f}jy33&��l�3����Gܐ _i~���b4Rt��F���Gc샼�[BR�v1���-�O��QcѨ�-��6�u�%x^��w��տʣM�U�����o%���N��;�����Q�ڹA	nzm31I˥�o���fJ�<��y�K{��#uu>�ɦ%_�_���N9wl#a I�Ҥ��H���d�5T0��@쉕��^߬���5����i���6�D��lu��I��hS��A��)� ,;^�~�{3�ЎO|P�ǆ���( 7t�N��� ����T�x�q���Gf���x�(_���%�J@���b�U3���� ���G��9L]!���E��Uo��-����s��J��_�Ï2��+�p/��;Y"���٦�j0%'���`s��xw)���,Q)��֛P��Z/�豯�̢���e�z�@Z/X�bߦb�]6E�t�c�M�j$�=��Xiܓ<�R�M�{�ak7�x����5���d�-����zO���(x��X�o��1�l��O�R`&ݕ|�*�z��+ȝ�]^��*@����{�̧�����e��5��~�H�q#I��a����*�\Ed�SP��f�p#�5*MH���J�h��4u�C*V��|�&�N���$��dd||��ӟx�������g��2;;`���V$jOn6��_�ƾ-X ��11S���[!-9G�\?�#�y����i�Ɣ�wP]!����'zo�]�����An�>d�ߍrT�~%�����`L�c��Ph7���06�I_P��f:h(���M����eP�΋�
895E���"�G�8E��H%�T��'��;>]�.� gv��l]喞�����>y�v�D����vV�#O�'XUՌ���^5a�h��1Q>o�3웯^��q] ��= o�˓�(��7�)(Fnhǂ5L�-��>��:\[������	������"��`GX��F�����C��VM���]�
VV9L�I?�M�u�b����i�����=I�1�ПJ2�d�͚gw�Ԟ��F.�-�x�qK�N��nE�O�К�.��~�o��vɋ<+��_R��rU�����E(tL�l앾~T�����C*�*d 8��Ch������O��]�Xf3��5��W2XO�����_F���.�nTC�|n^==`Ԩe&�#ii�wh���Bܬ�v��Yu߭���O��sN4�����h)�Â ��=�%{��!�O�x]��B�� ��mn����U�wH�!�5��ܔ��$�X�x���Q�fV�5�V0��W��
v0K�=�6?�ٜ-�q�(B��l�B����,�R���7:��v����T�H%Q(��R��0�	�|hk����tk��j�:�d�5M�b�~e9�,���8�8��]�%���4b�ޚ��3xA�;1�t��E�^����e�_ =VgRz6���� �Дi��I�r�w'�8�w���D�d��Rɀӗ��J}�Jp�8���J�=]�X���q]c�x%��uW`T�G�Jv�� �i���q���*fXkƵ������Ų0M}���uc���ٮ��t���*�Y��
/��5�z�������}.�m������)N����/�|:���I�aO��:"ט߮��|Yv\���W�Gw�z5��w�S���+Ot ��d��[u��\��@;Y��tx��Ʒ�sSl�\W�;�����|͖�2G|���B��PR�oo���zlll�9�yN3-j�9Kь'"dh�mh�3���HR��D��<֩�s7��6�#�S��͏��cM'��v?��S���^�AE%W>A,��
a�<�R���6�^��*Ӽ�eO��Y!w��L�x�׫�;ְ;wLк����{��t��8�&;����(�.c���|[`�w(ĽP����EE�HH.
���ny
���xQ'Hc���kf#[xoN���S�1�󱃈���C2ҭO���&�D����6W��3�u�|����_ً��D��m\4�Y�&_��FΜ�u��nb�~��e���DO��W��_�G��k�IzF�7�{I����JM����Z>��F{��C�U�5^�����?*.���hݡ�URR�eo	�-G�*, ;k3��Q��(���j�Q��S�ta�z����D@�m�����"=�b�ѓ�f��S%���\1��1�,�q�.�-����jH|���ꪄ� �j^�W�g[�u�x�Y48��
���[�l5Vj�����ފ}��-M���]�L1ٰ�擡O(��m�w|G�Ff_r�'���o{Y��6b�00Iʫ�NNF] ��#�G1�/ƂU=�,<��$�1
�:{F�n��fyQ����WDd�,��i��}6U��D��΢'Y�X�d�K�|��19V�֕o��VDщ�:=��%
e��9�8_knZ5k6&h*.&nI��H]y�8'���7 ���O����h��ŋ���O�}#|�6�A����ǀnY~t�E�/I{�K t�i@)��L8&������M�߶@���ޛ�9C�Y���x��#W�7�)��\�i�qj���-	��o��Y�7Mֶ6�q��ƲD������0ܡ��cO7�*��1	V˥�w�K��j��Z��0�ޔe,Z ���� {�^��6�FJ��I��ɜYl�
7����ok��)����p��>]��{��syTΓG�k8�^q����Yi���:7�d~��:�����ڟ��R�HI�o�wW�uo)���j+�r���*
� ���EJ�Z�4�+����>��y͖�y��mSB��{���>#
E-�[��8JH�x�U{���m �Can.v���	���)y�n5�);�����zY��Q�	�k+�[p����Ǔ���D@
�����Nem)5ad�LY��	7�*�.%�xa������e�ݠ��E��Ek�[�D���ԻSRN�pS����Ɍ,�qv�)h� �,O9W
��!�s��n����U��/m���m��	Y&m���Ť\0�?�z�'��"!N;8R�Y���s�!?X�[`39070L&]�G9�-H!j�=�n�S$~�n�^���Gg;m�WO�A�}P���z��d�W\p�/��m�Lc��umꌗ��<�!��fX�`�����
OM��(�Ռ��L���V�!�l��+����/�A�0�n�jzu�#�'�"3��<U�OB��U���*:D��ϛ2�c``@#��}U�9�=p����Q��:%=`clN�w�0Hn<�~ qBJ��"��kՎG%w����K�mE`a"��͐�㆛3�E�Ѥ�:���l����R��+{�3�I1��.���)ӑ<��P���Q7g�7_�x�q��[�re\*����c_7��
(���M���q_�B8ߐ�D�a�tĤ���v��f�E��n�KѤ8�m/����+��y�d�$��=��)�@��w~��b�l<�5ZW��v�\8�,�jy�� I�9w���7y�k�j�O-W<x}��;|�!��e%>Ɠ���:ш�,SWl��ݞ��S�ǚ��:5zx��_�

w�|���JWo`Y��p�5�E+@it�k��q#2���9X�U���S���+[�oZ�~� ��Ksp�3C#�-��-�N��]wf��X����R&b�M}0�5ވ�T���w.�\M�����8;�O>P��0Y�1�!�z��xi�B��U��[�{�QO�K�_F7��$L����%��2+��
����T�η���K���<��heԆw���΅����7��/�o�	Ҳu�Lh���ͭDW`O�#��%&P��Re��! ��%pp^0Ĉ3/A��]��p��M�{�!U7���O��1%���BggM��O��JDm?)^JUΨG�"�(�g�J\D���:��#ݦ'������>mt.��yZ��9R�uU�49|���lN�2�!T�������va,y93�r��;<���#�e�� ]�� �����S��lE*�:g
M�u�W�Vvz�jA˽:��(�r�Pm��a��jh"(%C3�m� ��v�ҝM��y���H���z�Ѹ�0����)�+��,Y冊�+?�yB��:z&�+L�؏�a��-+��!�������̑���ᱱw�;�C��<T��H:���۳o�Meu�*�OD=h^?ư��6���~�N4��?>���g���{�E���
�Zϔ�^-Y�|Asa;��K<��,M��8�z_W��Q�Ե]*Y�e2�o�R!��w�#6��ւ9�:�U'&��ŷ��Jؠ�4ژ߿��N}&,L�5����Z�H�y��FI�Bꣾ Co����[�i?.���$�����H�N][[�g�7S����%��
!��`���:�6��N� -�Ȋf�ObZ��8�kG�9VD=?�Wt{�+���9�q}-D�ҒZU��^ɔ_�
��b��U��f�o��ԛ���Hg�YV����ɾ�t���Q�zrOqYb	����^�96��7 �Ặ����K�eLMt�����K�9I^ܗ�W­���~0��Ճ��d#��1R|GG�ڋmXv17�iÚ���v�7�o�%E��������(�%�|V�-$���D�0����wEM3�����O�wtV��i�^�qGY�ɫ�:����:���T��5"Tf��ZVC��R�?r,I��3�qo�y5���۶�^ ޒ�%~I͡q�i�9�ף�ພu2�K/3"�c,�l����m{A�GQgL�R��# nBS�i|�=O��D"������rx!����s]e
r�F�a\
�Zۇ�뚶�H�*�3�y}K��Bf�R�(��s�-�X��Q��J����7f��n���'"���{
�K�ȫe[��`�`�z����P��C�Y�y�f��z_�u�c	��j:C�b-�|4�8V����'U"Zc��7�����0+�6Z�W;��;&;~Ԕ�{��Q���lb.���
\N��`�Ɋ�J�d���"���/z�|sŪ3�SS�yj�L�=�:n��b�����L��IG!0�������a��,Y�q�G���Ø!����g�����_Z��n#M�J��H����K&����z�'M�B��I+����1�����j��2q�妙#<���xݫ��ZW�W�;�&3�v�IE���I`cc�\�uU:L�5�~�86�{�j����`��;�3������a�&~���[��IY��Ϲ��?�T��}���]_f�j����IU<僜Z�*��B��'f���نG�V޻몵6.-o��' *)��j�f�8�Q�������e��aj'^���U��A)� Ą���"X*��{�+��Y�L��@��ܲo�b����	��a�A�^B��/v�:�\tϺ�/�] @u�L�z���6 �]��wZI�55�����a��:\y<�ZL�ۮ4��T�嘐|��Q#��͢�RO���c��gxnܨ����ژKGT��̶��vu,��G�>M<���G>�kó�D^�oH˱v�I%վ��-�o���V�k�q���HA3ǫi�؊��%��O����f3�U-��^g~�l�+3���0�П�+j��\&Eo�9W]v�XƎ���K	�H������H�^�=Ɛ�ۚ���g��Xa���U̯Oy1/��}�D5}����#����B�u]�u��m%�Zx�u��Ο�F鼗�>u��:�s��tx����p�����[�J�!��!�c=<Q�z`���a�.^\W��C����y�a��g'ޯf0PA��D�����v���rd�"�㌮J�k�gY݁(¼�f�X�}<F�ߘ�����L0q�Fw�ثZph+R���a���t�@�(��{܉r�X$̛����޾�F'��_�7�N�ԫ�����0�b�	�Q�����m�cK�Ep�����m|F N����z�������Z[�^�� �ICl��	�^�OC�8�M@��93����ZYWJ�\�M�9�O$�ʗ�OC���\�7�?7��`0�&� 
��,u�l���TE�,M��9��j����f��P�����# 9=6U��5�(=�{���G?0fD n�"?��e��|���p�_�����E�'L�eGY-�v���*z�yE�����.,1Y^ԣ�Ƃ&2<�o	���!^͖dh{�Y4+�L����ђ>��`j��_{����#�~]G�E�ryҜ���,�!|E^'�J�A�}�b%Wl���]�Yϊ��{�ġ|��lQ�\��.Mu5MA� ��?qe���K��mm�ޕ�lwĳ)]~x�W�򔸐D���F���1.dgDF�3�����u�s��
��4�(��~nH�<��{ү7����H�!��'F\w� m��yo0g���|zl�[hT�fO��y�7#s_Sy�D�i�Ϛ��Y�dC�Y��d"J<�+Z	4>��ȇU7A%T(u�8U`�xF�gJ��t��T9r��q.�)�#�@߮{ygҴO1�.u����J�s�b�,���*�^��m�x�L���^�_Q`���ғ>������n��*�P�_d� MB���5��尃$��-�m�\��^��˚1��G$RY"*����m��cR�r5����>�F�����������ms��(��|���YS9��{��BRQ#ToX��w���3ȶu[����T����hrF��C�����yf`���Ԝ�y�ӭ�&?0x/�$ ��,���&�������CI�Գ���FN"s�<==�|�#����~&�抋����v_R},�!U�bob&���䑼\�h@�F��v�xw�������$9�U5�v��-C+�Ku�h_Pu�ؾ��k��^يqBF�Q��tK�P�/��һ��'���|Ax49�ƛ�P;6�/c0M^i\�4��i5/ݢ携V���>����6S~+�9��/����t�2�\PGĊ7��<����F�oh����O��d��VҖ�x��cb�g��H<�p8ܠ���]{�h8S��w�.ҧ����Y����ޣ��wܲ� Ld��4޵3��)��0�O	�h������5&F.Q�Kx���.�Ў��/4nO�ԑ�[���n���v#�y��U�Gh&�Y��[�eN�1㚿������p���V�u
�lzr>;z��^��N�4%5N�����]v�B�	(��%�;<0�`�P\&Ҩ��"��DDD����%��¡�2;�y-��'峺_��<�#�W��w,�����nH20L��.@��D�Ueq�#�,\���dA��������/�?_�u�R$}|�أ��j0ʈ;�E/����j�T�c$48����E�:�ڣ��	�3�\�&���\�
[%9�Ӕ�[r����}��	ͫ8$�����t>��V�")������3�.'D���'ۆ��R����{�e #�w5F�ȏ��,߸E��=_���IQ�X�)i*����3m�I��u�Ѩ��7"!�kbu�X�5��}I*t�Ru�gy��غn��99�&���P����"Z�X�I�,ϻ�,q;bN-�/��zn����e�q?^+��[�o���^�lmA�&Q�7�w�\w�n���Y�X�C�@�� @@�?���ͮi���݊�S\JCqi���S ���V�ŵhq�ܵ8	V��]��y�极�C����ڹK~��3'�.�ee���U�B|����*���������1o7KAU�+��Q�SJ��0�g�.�?X����[	�x	^^���q�^�=�z"�
)s�q^�� j~KU��d��Y(�9/��:ܭTX��0�R�E����{�Uj|�Z�LTr�m����Nʹ�ҧ[6n�Tg6�'I�s��_BL���>`�O�o���")n�J��MMH;,}�`�̋Wk1E��EMN�,�e�J�YV���7;AB�x�V��~��==�_Nru��@#�p 1��O�f:��'}�l��TP�
�[��������$Y�I�ϒ�x�ە��A��D�"���ӗ�$UaE�����}v��O�}g«7���H��_�T��GƶZ��^ �ˤN6~��������@��ab�'q~5��D}�.�A�ĳ⮡�XB�w��@����X>�ήK����!���T������g9p:j�;K���Ӑ����g��������wpd�!�ǌ�	8}\�����_m~��(�H���[	&�;*�~ES���ߜ�ߐ�+�t��,Ѵ1o��ꑀ�d[��z��qWsۦ�6�ZYjeȋĪ�zaT�Nw"��W^{Q�Uۛx�dk�U{�<Fh�����PM��N�`��hU�d�_\Gk��(`�gy��A�R��0v6�կ����Ը�h�{tt)AX�%��ws�4�RB��QHK��JR��Y��o"�!F&5drR�v���i��+5�l��C;��/�=MA�D���q�׬"��U���=+r�P��r���2���O��p�j�W(a��3iz��	ڛ'�i^x�8n������D%J�.���)�rR��Xկ����|^���4�O��
��R��M�Дy��K}�N/A롨�ٙ�y��ll�~u��=���J)nx��A�e��?+�XA�#���v�ŮX1��y�z�������ګ����T��cQ��(u���d#	\�ՆT}�j����l�3�b���P���6��ͫOj`�F'�CP���>=��dX.��o��f,̩��&�䴵���o�W�3�_�%���B��	�s�|K/ ���g�M�y�����	�O;i�g�o��j2�c�]5@�<X׮:�66"_^!��h
j��oA�]�z=b<�92 ��nұ��z*���@,�3�#��E#�(N3�]�')�',��w�_%0�Z�>-�뭇��?T����Al�����y�Wf��4PE��G��,yt��,��H����{�ɅL����6b����udKXH�tߧ�X�=/��LOU�w �Mz���[����7��""ˁ{7��A˿b�}�^��C+��>��~���pd��8�ɫ�#����r��Gx����ڰ���a�ƴ�%.����k�%�-՚]w&<�����Iu5i�r��K���j����-�\�n{B���fӢI�F_$�<�NF��aSv7��d���N3cBK �;O�13�_mv��du���i���Pu���R��Gn�ƪ6�ƮnR#��52t5���f\b�q��9/1�o������#_��Px��s�1��������2�sv�9�2�<9MN)�z�{�M#��A�c#��]����ě�?8�V{��F�V���*_�nB������q(��]���g�6�8I�s[�Х���� �`�V��A��N۸\v2\��qZi%(/g ��Yԯz��#g����r����F����lD���[�Й�Jr-c����FC�(�OD��ԅ �2���Q����#7c>]��mo�.>C���l_vP���Se�ǭ#�O�݅�^?`���z����NQw�\�� ��:���O��Q1UG��@�te�U!Ѕ�B'oG�=O��=�9�����7;S�D;�];����������a�Pd�!K�9���m�N/"�[��ZH�'�-�S�^[�x��9������5�����b����������.+Q�7_�6^jv�
���=�-�We��ۄ�e��BM��O�2����_�`��a�*"�;^�y	�Η�f�&ݖؘ}���}V~/���g^�V���e��+�a���:�����L9�(��g.�|��#�g^,b�E�
B�'3/+ս��p�����g�����DG�5"�F��K��!�	[dՓDS�ry��x`4�J�ޫ�ax� �'mS��p�~V�>>��h"V��{_�d�POe��� ��F�HZ�{}������+����� ���s@݀j�g���U1J%��;���{;�����e�J������c�|�	f���"���9o���%�X.WqԃI}�ڇd��o�i�����b�������L���u�$T���~��q6N���JF#��7#�o�}�ȪAG�uԐPݾ��Řd]���O��#��F��<�A�h�?!�jN^��ۋ��g*o��l��熃ߩ`>Gk݌�u^F����ۃ:�����G߶����8�A���q��{�d�H܁���4����, n��U�*5V�"J�M~k�Z38\���AB���H�3�)k��3R���pe���c�2c��~y^��YVň8&�Lˍ5����H���Y	��=��ŵ�؃�V�H[\���k�����f����u��������||!��{*�{{'X�2e��

8/�i���'�D�3 r3�p�tԟ�KԲR�
Ӵ�Q��$C�&!m���Џ�<�^1����~�~�xL�pQ{�M��
�<G��w����[�ʇ��C	!y�H�Y7��wC���S=?�
)m�1�����u*�~F���b�L��A��nF���d,�M:ƭ����ȞL>jk��}�x�,,,�N|�=xS��y��j{�i��+��虑4}�7�Y�as�����+��?_�i����z�̼g"����*�/jhK�XC��;�)��N�B �^��N�A�ښ	"�vu�F�!X�G\,nՏ��������S<{���>��D��1 �c�U!��-DG���[9МJ+(�sk����s�LKG<r
�p<�����Zg)6�j�-Nt~~���
�6�D�J��h�����`*��d�Yxt�}��II��j��6HS���OĉВX'�z 5"@���IBJ*�M4N�+�=�����r�	lzex��:���r4���ٔ.׮�?W�<i	�k�m\�/�q�4`
`ꬷ����x�ڍ 	�̰�N�󋋍L�jwjK�8�7�Z���䊥�%�_d��U	�B)m���~Y.6�(�{�.�f���3?����?�$l�hjl�R@���B�V�R*�����Ŀ�y��iV���)�/L����ȳ���i${C�䄳��7�P�YgV�l�=��;K(x�>l��mӦ%̽�]��}O��$a"לF[WD��M]��)�ݵ�8�����iG���n7��k�gY�9myy�4I��O�L{�o����9:�"r�v�f�~M&薕^�����
�@A����&����71�2 3�I5��sZ�{ā�9kS��O���xm�K���j�T�u���9�0�F���Dp̄��<mH���C�9`mwiCؕ�6��{fc��k�%�B�\Xc�O��% 
]����魆l��)
�T/K�Zv7���1E�>E���6��9Η��y����ڔ��T����u�ZM��P:�������z�8�^tJ�Ȏz�(2Xj�����Q�0�BP�� �d���ܸ舋�C�����[���efy�1��0�/�8��aO\��V���ʐL�&ǜ'�.)5��n��h�bS�);�ro\������ۘm�� �A��E}pҕ�R�ep�v7~+s+n��E�����Ĕᖮg\�[�>ΩgKp�(�nk��4?L	�aw���RɎ����~�A����[v��o������)��qωe#K>��T#��
u��u$˫��޳IG�&T��_u�����y�A�~ü�k֐�ĸ���Ĕ�s�tZHk����2�����f;���Aۭ�b��\��eX<	l�X��6�e�����S�Hl��W����Z�G��m}6 �X�5���x�h��m�DT��� �>��9����.*N�;V'���b#�p%+kT� %��I�Ml�[gD�&ݜA._���:��O�{~�˥L��<��f���t�~�e�%�6�Jq����zҘ�lW����m��U�Ɨ����jS���S���ҋdۺ�\��)Sᨂ�6L�|
��'�N���}�r�sX���,���E;p�|��F��P�B���[���B �^��M�I`�ː�e%W�i���ճ5�Gx8�A�0�	z�S��L륚�	G���e�zxԓi�~�CV���E#6���ۗ�N&�6�Z.s��s���p�|u�_p"�$nUV��r�w*��Wow��m�%�Y����˴!�k*;	��O�Lټ��5i[�dj���*<��fKQ¾:�ZC\��� %����C�i�| ���"������Y
���t���(2��?.��k 	`���ƿ^��Z+�����R�fk�?��no��ı���]G�F0�D�A�ƴ�~�}|����|���٩�ZY���cԊ�JU1�'�[��13d�U�vY��^��>@K�\L�m�c��h��K�<��I/�3~��4B��'�Z�<��1�;�7;����n��cuC����L�cy;w��]�γuM�~�Dv��Dni�#���W+�o��.�m���oO-˗Q۷"czs���گ�311r���Ai_�c����I�j^c�D����`aqg�0Q)茍�`�ض�(�l�}��Ôp`<�aHP;]Rg�]��lx�����#�k�J�5�4�"2NHU�?�Ѫ�U_��b^Ub�*���S?�N?��v�r��G!�͍LL������D۾����^%t�"�� �'R5R�S�Bf�;��^�s�}>Y�����41����6"����-�dU:�ǝ���@<�'���6M�OY�_k�e�(��
��ǰ�T���@���C> JD9�}�����N���z��gJ�%W�r�~�&A��:�xd���!�i��'���V'F�f��S�/x�O+u���*/�?7��|�T�-�d#���H'��v�ګ��R{�Tm�l�@ʫ<(��8<��9���=�ݞ��8q(�T����M9e�����!W�7��8i�#fǃ�6�{~a�Y��"6�K�ΕW}2y��9B�al�Pp�nΧW�R�4����[�����f��Nl�}�~�eOm-_���6�t�(�R�~��}I!��;vNU���߂\���őD�{�@���uM��i��-e�߳�����1Ѝ���ظ�;S���GJ����Q��K�r����9�ҝ�e.$ѓ�U)qp��4�vN%<��,)�"������h�L%��uz7y�m��`�`�_C�f^b���Fm'�PG�gD�B���9�)��ׂB߻F����P`\N�ާŵ�d��}&�D�/c��פ�dk.O=�8��Q/�|V�WJ=%a���UJ��o���������\�k���B �Ͽ�Z=��"��i��0	Uuu�$E3䆜}���,�S�E��n�\9*Ȯ�ҩ&�$�ʎ0Ɯ�SW�,D�lv/<�����Z0譊���z��LH�q0S͌�?���������f����z����bv����L)1��h˫l�	�V�����\).��3��r�q�W�6ږ)h�?�ʿ���i�l^��T�v���w�m=}�}�i��Bhi��X`l�M(w�Ӎ*y1�4��Ŷ"@���#>Iɸ�#�:�������6_S��c)z��f��/���<��ue���&.bEYY kX�_+3ee�v���P��s��� �{�I�m.)^���f"ޜ�א@e���� r�6���b�ۣ��W�"�c*�k�|D���U�۵�TB��t��+���i����,^��f(�ߥV��6�\>��
��d�?�	[XV.�O`�[GDF�\�� �����71�����{o�٧Fجb����̷�/#�8aevi>r��vN�=��k�B����7DCz�?���pc>�����W��
K?L�����t����O�ǲ�'���/���\�-�0�)���-:X�;ݹT�t�~��,�f�q$�m��B�D���/�R/�������[����%���V��L�i0l�#�@�㰕@��� h�_�������va����YEs��ʁA+�K'�>+[BT��rΏ�/2�eH����2x0xڵ���I���S+�Ab�eDp���1�]š7&�'Ϥ��}��(�Iʱ������fܮ- �Iw�)����'ө=�){=�nD����x���ɼ|ʷᚍv-j����Ck�hu��@�i����F��ْK�O��a�[��['��Z��r�������#~)޹OߛtW��J�+h0�1��Fޠ}�¥��z���K���sK$�*�Xtc5{�o��qew���g�}�HJ�
����(�.ϯ^��,�L��x�5t����,<<��J|gmPN�
8��w����.�@#s*�%b����B?�~�30��Ya[����Ѡ$3�l�E�/;��O�J��F&�Y6F��k9�-НR_X�+6@�b���;y�Yμu)[ŌVP~(��ݣ@I��<�HA�I��'*>n��iH��-Iv�g�!����1=�S����O҃vS]����hy[����DR�R��ˑ�6��c5�ӯ�1�|�H�yFi��F�^�p'	�'��Q�j�.;4��bn9����n2����� E���׍�Q�2��g">:�#H�KKli����/+�hE���B��s\����1	7���Me	���1vx�^��?���X�0}�2�TJO����B�[�f�Q�6_��ч�Ē���Vnn�2Sw`���n�b	'wl\��U6j����6�C���K�tC1b��"�?���f\2���r�9��dL��%�+�l�FQr'��q�OQ�~й��s�z~g�m�v����)Ns���?����<R �m�qCbʧ9�}��#R@W�٬��VQ��*6�[a�<\,��M�V�R���vX�\{V���ɍ��@X"aƟ�A备 �Iaq�t'5��b[���@��P�-���ܠ����7q����	�o9�}^�O+\0=
H���s��qs��|�s�ы�6p]�I����'����V��G�VR[�v�OI�����|52X�b��o���]�U��̄)}�1�'�6���5�W���2�vÛ�a�07�T���ƶD�^��ߋT��yF�5�(�T��m�����͈�v�)���HխA�o�U|`3J�`O4G�˻�~���.%"���]��7��^������X=��;в���oq�f�3��2��}p���(~��	��*�Rּ숈Ӣ.
?P��ԫ�Xf�*�U·�W��Ry$���昕�L�_ ��Bg���t�f���bײ|}�����E�(��aqܳ��+��@�?7�e�dRe�j�zٴ#vJ͎��)30�$X��!?�'��u=cod_C�D8��f8�����O��wlmm�q���lj�e'��K ��v���=�2��b��Y�=�a�p�BG?��0�|�lw��R�g��`CD��}�|v]���-���O�(�"�k>�Cr�
�=gzM���P�NT���<�3�l*ƀ!�R��,�c��t)G�)W�����ץ|�f�C����4���pό(q����8��\�wZ���4��sF����p���gf�R7�M���>�s�AE�a-�q�������D���Ueړ���~zJad ����W"�`�,��+ ����T��l��i7VJ��?��:��Yn�( �S�0�k�K�os�}�\;7&'�=�:��:��6�����
F��3�
��QG�{</=9���'�c!.!֕Os���h��M��p�E������ԥ����!���jS?�LG�@���;���,�a9\��M�Ç�'Zp;�g[�z��I��q8���E�� �qXb�K�/��<$�\<���֖$��¸J����+�:�G�k�N)qS
�秃(���8�͐˭gX�\��GC&`C���8��S�Q��F�1�A���8�;,VW�4�]=4絺^.&�8��X�樏��Wk��{e����΄����=xA|���������QtT�A����ʊ�����Jh�X���kv��{����'�i��c�H�'���9 ��,��3��¶<LNJ��Z����}�O�B��j������F�1��͠n"{V�V��y�?N�j��1ï��UT��>�ꘗ���i���k�л��āI��6��+D]Rn����%X1���%*���qcIa��6i��� #u[�F���$d�g�(.f�$�����@
K��'�O#�	����v2�GO꽯��7UoC�������ߌ���X~7��憨5�Y�2)�&�4P
�VM$~�b�`HB�:%j(c$��k����xbqU�&�q���N�}ԝ|��.�;�e6u�~���`��?[K�x?>:H�*�Z5�M~z�3
�q�u}�f�wn���2�sh�D��D���?c1{�}����D�=H0�]�%���]Z���ᴃ�c��"�	B�=�b�?�'�ž>ݚ>q��IK~�������M�1�B!�������[�]��m��lf<؞<H�N{ZX��x
B��t1�dD2�\�7��7��$2�� ê���E��!dlr�����)G#c�(4-���8=wh��$�B��6�}�b�{�S��oh��x\8��
htd��n�su�W0�b�U<���/�? uk��r�vR"
\�7�u����˝+>6Tk�P�� z)����ӯR��"i�(��V�S�"���f�k1���p%���������]��l���Y9�j/�U�_m��Sa�eqH��ث���d' ?�)/��a�����f�(�N��Ћe�!D�哊4���u� NrYefX�%N����I8�*��k����/�6D�Md�̟��.�n��Mp��8�>���4`����p�r?gY4���Z�V����^��p;���tDb�ͤw�׮ۊ. h�EW��I���7��Bs�:�d��}'�W�Ќ��2k)�����`��Ǻ��x@L��/L����X�"@as.��õNj�6�;͖����t��s��?����眰&��&p��̄:}���,3��Ӡ�<��[��
�T�{�u�ZQ]}�V���J��� T�:� ��]�:�q��%܆Fr��_�����:ϋ�)��4��_�{���(��Š�y}̟@���v�V	��LA��!�H����P�M)0��H*�d�9֩��S'���Ki] � dCV��"AjK�G���ʚ�GZ�s�e8��H~ZDO�P3^�݅�
>�Bs�Q��O�'���ѳ��;w�ąLЪ+�\�P�?��
�����a�)��������ɷH�Q6�ZL���n��T���d/��}���u0��k!Vw{nx�'�$�(ܳf��y\`�(���#sÅ��::C���/}ahHw�9u����!p�ehs��=�_������$��7H�|
�s��ya�W �&}�M!���]�L�qȿE�b:a:i�G�x5X�w����H����Γ���r���p���ǈ�V���0D:�ͻ�jvw	��X�W[�Z4�O�擾����N���U�e�w�cW1�pk�3���4�M4Ņ4�:&��ƛXAl�lHL{IX�[��1 ��Z��µ&}��a�<���^�C��p�#Ϩ��}�Iu�˕J<���)��'���Q�(�+6�4��#<Bx�`�|Dpld�&�i����I�]7}�V��}�@��xA�_ӳ�>�+�m�l�2T#ny�6������f�;௛�"~I�%���� �[���S��aqhh��K�!41�^-���d�ŉ+��>�5�����q�a�0�R ���f�z���ƹ�NW�<���p��	�{i��<�6��s0�3����CG~w��^���N�k�0��K�>��z��#�ں=�A|����d	��@+�����vd経��j$۶��ESd���ZI�g��7��:学>J�_a�zp)�'ڱ�T�T{-J8��X._���UD�]���ʿu�i��Z��Ia~O��E�?�\F�Lr����޶�d�67�^f�y�Z�ܶ2�����}:/�\7�[':::4�� g���p�9ﰁ��o���Jp9'Q��?���Ԧh�'#�ku��j?\�s��^α4�Y�Fv��9�4'�� =/s�9�w�z�Em���}  P�
3�'4�\���r�	19,��/0X�ʁ,g{ReNrV��%6)~ءG$�8G+������rY��$."HJ��E�+����py��ߊzQK�A�6#��@7���,�F�,���R���վǇ����[փ�je,�=���z���87�(�I�T�������A��̍�0�,�J��_5�	��Y�ݧ~"9匘���0�Z[fs������a�$+��[LІF��/(��i�E�ǝ�kymZ�i�Fl���7k~��@�w�+���9��x�utt�õ��w��+E�u���x���<��X���#�|}q"���E ����g��%זTYj�I�wS�?�2X����U�*˺o�6`����[�lIX(�fOl�ÄE�� �,���7h9E96e޳pǜW�M�ө�KOD-b�%y2�MF�
��)��
�����Or�R���J�vu��A��f��)�/�3Լ[Ϯ�W��@W����S�5�ȱ��$F�i��C��&´hG��%�6ȂP�S�z6���D��`��*�-��-�o�c_Ӯ�M˛X����g�cW�R�Y!��`��{\U�2ȁ�c�!=/{`e��_�MŇ����P%�WN�P=��Y!�˅:�Q��
*9���k������#�8ǜ�$B$̝ &g�s6�%jq�i���WBب%u����A�Q�I�Ǜt��f*A��o�E��xy�bM�:o�kx5�;>�* �/�_�|i�ܹ��ZC�X���<þ��[I�C˵��@���.�F�5Q�#ݼ���>`@���EA�g���y�}�solXm����FJ���js"�Ε�P;�E͑\Ϧu�L�]��u�A��L�-�̇7癡_{[���������H1�V�]�k����Rs�g���8���m��GR��A�x���-3��\?��XK4ti{���]o���'�IkI�c&��?f��IL�����^+�8ތ��c~5&�4�Gl�%�ǃX��[9Xzh6�gd���%��j�/(���1��+�A4�թ`E�@�	-W֜S`��� s䄿~�B����+T�]��y��"�c�aR?dQ� ,��)�:Ơ!�Ѵ�� ��,�)6�}�{H��2nje��~o=�W_�Nj��׈ti�e��A3��%s�<��G
!T�{ŏ����hd��Y=0A�P�� 3������%^Odl!J/Ϝ6	���L��Ac%��
�&$Σ� �|4D&���հYZZ�/���@� :3�D���]���޿���I�������=%����G%���Kz?/���E��$�eKE]>*o���OH�A �8�t�IX��e�ʖYe������A��F^ꇻ�_���6��@����E�=v�λU��Yޓ�	�[3�Q�q��$�Q���3����lBA����J��ׄlON/cq�\��@�2�0p�S����y�> y!�Hu��q�������������U�,˅����T?�Z�	�� ��Z�ɡAߓ4
�{N�7��=�q��i<��r=�G�Xi,_u)ι�x�/�6�]~A�ē��!4��F�A1�Ft�r� KFc��Ɣ�Hܵ!+�b���/)��3{��K��6�L�s%��R"%]�GJ�y_��������_�(�sW�q��u�c�� ��3�v��B�E�m�n���`-��
�;+`����d"��fQ���9YcL�ĽF���^-G��U����B_�����h�;�Y����0�*�����b{S_��S�z�3j/���A�,4��ϕ��REƆ�ꤤ��j���w/�����ǩ�Q��
͈��*;T��J�Q�b��]˔����+@��f�par���Pr�Z���f?I�Nϔ��$p`�ދ���F>��⤍���q���2���ϟ/�np�DfŰ�3�M�I��B���/��v���v�Q���R޲�i�`�}�S�	�K	zC����[+#`��y�j�$A�*�ưn+G44�:�@~zzz>�f�Hi~�{Ǚ%�!Tz/v�i�I!�o%���<���ķ�����5F�n~uh*�6S)�]��_Uʂ\ԅA��ĕ�.��V���@*��G���I�w���/Lb����9��9��������y/�:ti�sV	��mQK.4!��A�),�ִx�[�msy�Q�7B��?rz���>>7G���ؑ���xn��B�Ecw.�d�${�*�ڍiW�^V�KU��Ta��r�E&)��p9ʲa��K	���x��-�L��@Xls0,���V�����"�湤�ԁL+�)w���q���t"(���2�ȋ�ܥ�Zy�ݦ.�*PS�Y�{E0�G�@���y�)��4�`����iB�ɜhS����)�������/�捉ؠ�/	7=�huPpJ�+rM�z�[ЛC�j��'��l+"IT���w�'�-�W�-���eT�����[AQ�#+~�u���7w��+oX;��*�2L±�Ɵwu �ް`a�n��`�Q1��j�v���w�����tS���%�����aq��aS[�wv�N��4|����r��%W�7��X�R��,���-��@w��;|��b��ҡ���b�B�E���b�K&��y7AFs�~������77&_��zu�mrqb����;�wi�r�e1N�3a���I���\�5@"�!��QW�"	�=]X7r�9�|�����,|��A� ��p��33������<'�M�t�W�*�t�:X d��E�q������+�n���� 2����^Y0~Ju����?��/l���Y�ƥ�l�G��d��.uTV��*K�.;�}��p�&���[vk��&��ps%����z�?��ٹ%h�ݣywN:<�N��h������ia�/��A��ỳ�Z:UTT�p�"���f�n4�F���e��!_�KC	T�c�N���"��>��1�R.� ���T+^�:y�/H|lKtP��?H9��d{��:2%^�3z��z�%o�#���ZG��W�&����d����/�Sj��bZr�p�S�ؾ�0:)��� ��{ҙt�6x��<�=�]c*ĥTB �n�������t��]�8y �����qe�A��7�LP�	���P��zql$\� @���חY8)|����Ȁ|Q�C{��G��e���� Gr�y;PP���߮]�l"���Z�b��}~'��d/�%k���܂�wj��m,�钸���sޙ�D�2t�;�K8��/���Y���Tze �b0���+� �Ϡ�=����C���KEv�����x�a��Kŉ��0��ǱF��?���F�<3���2R�_Ah�BA;y����+���?ի��F-�2�!�Ï��f��Uܤ��/>� U�{QT�ܡ�qdٝK/9�U�3�
V�N��ɥ�7�y�c=��0"�?����C#9����ӄ��n�	��>?����2��N9Ed��?�X��(���ѐ79��F��IFӋ�ȦN��JU��Þ3��E9O����"�;-)q�}R�x�ʭ���m?�t&�̷êO0��כ>ɿ�<������تb������� ~)wD�2�1&W������9~�{_2�Z�@z.W+��3v̌�U,��[�c�tX�j/��w���.K����ҳ'��b��p	���Hd�F���9���@�z�Y9c	�����V\�$<۠k+�k6�sAFv\����������C��t����q܋-
<$Of� �1�ڴ*�u��V�������߈�r�{%��O��%�7/%	`T��9|����+��G�
ı��SsQoph�T��5>x�Eo��Yԡ� 2Mpf�X^��� e^�А�K-�È��D4�B��_l=Gz�t�����~���ʿ���U<�t	��tԎ�F*���C<�ŵAd�N��S&!1CW��x�G�wF���0������cP?6.��Ǖ�[����p�7��ޚ��&���Nm�)x���
�j\vΖ��ݙ��C.D 7B$�8C�^+�Vi�>EbH�f�[oYZ�V�#�L���s����W�����إfg�xo/ZIi)�T�cݛ�o��cB<YtCZr֣��'7�k@Q�g��Ѫ1� ��Ԃ�h��8L�U?�@�8?Ĭ�)��㆏R��5etB��<��M�^��cfj5�z�N�ww���ju�qR�0LS�P|���A�!�x��n�2��=�(p]�_?���=����4�)�t�l�$�u������{o9i�cU�:uV���Ŧ���.\7� v��ٸ�XP�)���lH��ޜ�����y��Z{_G�X�5�:(�Ғ��S����}@�̶�ٚл�1*p�ճ64A�0���B�"S:�s{+�t؛SkDk�@:�j���4���l)�4c���a8dXޟ��<���سŽ�~��G�vw��M<�I��eiw`w��(31(9s
����s����(������XѾቃ��l{��Rn�\/RG�Yc�[ϐ����n���\澴4�ޓ���LRx˱���F��,�u���U>:���|!H���?�.躽T���EѰ���"f�L�n�C�,-FU��O��n����^r*�pL��7�@T�<2�>3՞u�	�ج�wZwgm�&��]7�v��3�y%����7��X1��rNm*��լ����M�KMD�t�0��}�+���$.�z��P.Wu%� qzɲ>��m�R�c��Н����~��മb�a�i�݌c�.�y6;���-*!�A֦C�g_��p��@����4��8�z3���V+�[n�������h��Rm��`!�Z
���.$�W�[T��Mr��/w�*G �gF�4ۈ��8jJۓ���\nPݥ�rMQ��+>5��wڵ��v��R�>m[�Vf���h��w�'_�����{�y^�<���������$�k�~_��;�mt��>��H��H��e��?��SP����Xw�R8�PЫ�~�Lg��}B�C7#8�M���U�b���V�¬i��D�B�{i�4:uP���Uׂ���R��<�J"���/���E��a6��f��#A��(鱐%MH��Ĭ�E��ó?ۮ�*9�P��կ\:ux+s�C�X���T�W`;��sN��'�R q��hv�1��8�~Dd��q?*���Ӎ5��j�+�4Ҵ�"/-2�F�X�5�)c�X�S0�
/�i�g�=s�*A��V���zNj~��.а�E�[�~���ܦ��޲@^��\=����u�cqS�����x����,c��q�;C|�!�-f�N8QbDy+���h|�I�}e��=#�)?�"Y��v�@�ʓ��'/�E�|�Ghʏ�+v�dM����$���Z�C�m���X߂H�";]��j�����ȝ��.��&�;��O9�W�Lۅ(�vK���l|�0܎#���g]dE(ɕq�&�̶��-�6[��`��3��;��2�g��&U�&qSBg���r��;��m�9��;��8O�aP�C?;�`���+�-�zӬ+[��!qI�8)��s3k+��7T�WWV�)��+������4�[��7�]��6�o�J:-�N���@��,�M��UѱnI��]��P���g�cx���=�K�=��E���E� �m��%����"��8�9��kf�+������֓�;���?�L 
8�ŕ�҅��V�H�����H�����e�܉L3���T R��Gl9;*�@�����ĩ2����"��A8`�eH��0�oE��|� �|�H�E��S�MjK�7��d��P>/ ^��:WN�K���������Iim=�&��Z�(�qt�In�ڕ"F�m6�Ra/9�����͚d�]{{���`��v�}PIB+���[#��4[��A�EZ�U�A��!����>^v�W����lې���!����s���G�ru��N=��>T;�m=����K
U?�J�0��-�HLyG'�,�.�F�5{�]b�o]!�(��%�v(�e7�W�W�����5>�͔WN[�����R�&��:_{����TǍ~�7LUL�, ���������֡���|"H��j5��R��m�:e{-�c���P�%9w�y"�:)M��ra��U&�PO`��\��^4�[g�O���ȼ�����C�ɹ�Y}B�'��ƦI��ձX���õ��q�7����l�����	�? �j8?Ĕ<�{X�q�\:Y8HR������� Y&�i�N�̅��p�8��/@�&)p���V\C&�Cdl�wM� �V���I`:7A�-*��1�����aM~�� �"H"%-- �0P�S@iҍ��(	�����56�cҌn�F����|��ϵ����y����_��<�9g��n۠ϛy���G�M����j�ӇY���R>�����u�z� 7.� �[�z�9�� �L}â^<�}�޷*�g�l=�Cdu_�F�E	��4�]{# ]L��/�
2�D�-�e5��l���x�g�JzN���V.%�T���5�G|9�� �%�#� �fI��yxe��{�����~�����Mءl���������_��|�N�;��^s�WI��(�[��ģ���շ��*� \;�|�v�?9��1J�f�s�?K�8`�ĢMZJ�򬨣���B���f:��w��ּ��o��~��{�ڟ�g�A�ݼKݛ�?:��z�۶VS7�`��sj��8U�邒.^�H��(xq�V�@yyz�m�-�I)�A,ǈ��
vA�>������[;Rj��/��鍫�x���7��'I�Y���1��˂e4�yPږ�v���a�����{���i9-\�J��n'�{�����.��˷��	4�ˠ�HJ�=Xc�%��ɭ��m��ݍ6S�Ԛ(�~�O��������u�(��x��S��}���3LDݳ��p!�*�;+��	�N�u/+t��'��&~-�Kɽ�GZC�p��E��	���	h�)��1c�:�u�:I(#sz�<�M���x���Fz$��2f�>���G���X.��� h�/d�#ZT�l+�;�22y�I�'�Cd�m�g����{E�|��=nq����z��ѫ��mC�HD���;L:/�` _�n�*�9XÂM!ȅq��0�ĐK�t�=8�\)�ޓ���?���J�}�@��˱ǖ����5��h�,:���럒}s����u$�u��}]��摵�`Q#�ȓg*��ۛ�*%�������Z�!G9����� ��D�I�@��NLB������C������z����-�0iǈ�4�g//��Z�?LEz���
9��#��'��a��7��L�5ng�_{uC���ւ�[C��W�i/.O��=���(��J�h��Oz�H;�3,��NE|�Mi�d\�;��~�:/�5��	�E=�.-P[`9qN�W �8=n>prT�ϸ�:�����9��W��o	y��Y�t�qT��߂�V���0R��Xn!���ָR�B���r�.Jw��^�gcI l�N�4#>}=e��r��k���:4���W�0>�^p͡D�3�Ӑ�'!:\�XbkŻzjh��G7����,�E9��ID~�,�=/{�A6U�����7{cz����0 ���¡�,@R)q���\U>Jl|�����I~s�-s'8*�;n�n_�s�}U��ѳnc�w�r�ҵ.�<�$Ty�x[�o�} Sg&b7L\��dXp��.���
�i���]U�?e3���oC
��% a�<+5�j/r�O�=�2���ѥ�yr�}��%����&
����MY:T9��n��T��d��og��Q�5�6�W̌ח5���M�*�OB���]V}m�LE�B�����Q�L^���j⋼9l��Y�Pwe?U���I��f�4|��5����WeJ���l2e��I3�g�z0��r��^K.E�������q
Ċ^DR}�M��܂�Yk�%�_��uKىrQ)����[Q�B�q���Ie����/x�{$�t��z�az^R��E[!9�������y�a	݇�{��E����a�Z\���Ř����k߿��?�v�ͻmd�=�}���n$'��S�T��դz���Z������
���E{&�>%j�g����������o-@�R��j\�HJ	�:�I�qљ�S���QҖ�!/��ǥ�T��S��Ý+�L���1�}�����3��n���kF��[�g��������D/��-DD��)�{F*�e��=�%����7l�8�*�HY(yj�1�$igw�sZq�0_���3 4� ���ο�������8��h��P��6��H	�H�[br��7�����N~G9	�-N+^ H�8�����1D�l��D����X���囈Юo���Ogr*�ˣ�e*i�M��o�sC)ԧb�]��C-�m �%�Y�z�fD�g���3�����K��^���=Vs�"����\��u��1��}9c/�[��N�z��X�?�eF���]�nF��>�UkY4�9�gψ�ˈ�YV�����ڸ݋t�ͷlI���}J���gMM�8���.�|x?��Y�힟���k�憊U�qC���A$��ϰGֳ= �e�+��i��ހJ�2,��ac�ޖ� ��ė������'�=��_{HJ˶߇x�o<���U�|B��y���j,���ݲ�`�T��H(�n8�V�&[qdx�S��\|��s����w�G�-��ϮL�yx�y�d	�%�w���s�)tzo�H��͹?���6���F�[�$$~,�~̴� 
�.��Tj�n�,���`�ѲZ�7��"�CO�:f$�����D�����-���d�����'��⧎���m�i=a*}T���o��'�L�	����w�0c�rRN?)���b�G)�&���3�]�3��,���9yZ$�����KjU�a�w���t22�V��F2����l�9_�{�͠�i�J"d,[(i��YfS_d�N�sui�̬��^κșs�}��SPa5-p ^�I�s�[9�C㭶P�數zvw�����=�l0�{�0�KCbr�l�	�����j��ì��*�(���&��\N��8���� �	��>��L>h��"��RIE�i?�;����6p�gQ2]x�J��N�($�'陙vo�5p��#�
��Q3r�Ch���2�QU��W���vf�:V�����'��/�j;°�e[p�^��P� 7d"���ǲ���sxPis��%�絷���ˍ;ɲTQw���8���^�Ϯ����w�Ҽe�w�-���sw@�?�`̷�ZI��j�i��$���D/4X�FkfW\O̡86�ԬKЄ)
)`�q
�e�B��4�}Ob�e�;|[��G��Յm�aq�g�tPDGb6�05���)U	��.+���!G��5���O�=<B�Y�O�mm�@�Q�ȁ7�����]�z<;	ųLBS�k�$�Ԗ��?x�[�YcF��_Y��o鐜�M��q��څ:Q�J3i��p�~qJ�Y�;���@����K�L�#��S���|�h�����d������F�zA2㊔h�}br &`�������L�����W�x$fL�f��/�ǌ���S���s�%���+ �/�����Xc}k�R��*&���F����z��g����zc?��)��.Dkh��� 8Uj����#^������h���q�-��&���?�,�s�>�o�,xI��e���is��̦""4ݳDz{�H��~te�\rY/#Pݴn�5�>�u[T��+>Y�W�e7'�7REI��H�r�sF�5z�=�ْ��nw�<��<C/�6�Gb��_�e�ܴC�.�[���
4�ɥ�T��]�Y�d����А��0�9PG2	C���̑m���N\̞Ϣ�^���K}��w|�t��U�D�{�M~5��V|$�ɴ���*R�W�Dk�ݚ)�&��<�:n#�����z���B�PS��J��G.��'����x� �=�Pm����x���5.�v�l���l��(�|g1�l���̅�.�.�������L��խ��ݚ2�1,	!��l��!&<³��"_G��k%_�9vN��1��z���.�oc�x)Έ�6ņ����]�}�6,^�8u�~�|���X�e�
cJ}��-_����ߗ�뻗�;�R�[ 2��q��2-���'7[�9	�c3N6e&	�s�i˲��S6�m�!wM�.�aB�Rt�O�R��[T�L�\3��m͇l�����E�n��T�z�2���#�?�3�so��I^��]jFj������¾~�����h9�V˅�n��BHm���F�dn��^!;E1'jkm tR�ߦ�"#�S����zC�@�����ȧ���ֽ���K������m�o�aDYc,�O�؆�G>y�y�L��h�A!�B�0�aFT�eS
F�1GӤ���'U��@/{�<?.��te���8��gJ�Y�s�z���1�l��$�;�QY[��_LN��.� ˖�Z&Gu���:�pR�S��ޅu�犜��'m�ݏ���g�$#���""�b&�/f�$���[�r�f�j<��x) p�d���ϛ�,���S[��"v���9D���χ�,�I�m����R���U��B� P�oF�U�3�}M:[��)2��d�O9Xx掭��� '�t
�����S{� �{L\L)��o�)"`���i?+��z�v���(<6>��ώ��-��B�G�/�^�џV���yTS�Jͷf��T�pU������� ����	o�	�V>x�/�����*#�ڝ5:P'=���]�ݖ�N%߳�#^kA����xT����!��?��-F��r��G���ޖ~��̙�)UX���IV:V����tS��y��\���>L��Z��݋�vgv��H�����9,6FW�U�6�/�v辞�y��ަ��m��/�ʽ�8f��1x)�+f�?쒗i������wy���kJ_��� �3�*��Y���^�z+�]fa�D�\x�?��(�y���������ß���+PϢ��nߞ �̈́�`FJ��ֶ��4*uJR��u��x~踶*�+�~��k�/5��Z�8o���<������k�!�H�N���������E�-��=[c�7t��=�ǝ<���������gW��c�Ԗ���D���Y��G�E�DF���7��Fy"��ワ�%�kL�&�1r"!�f)e��ǋ������co^x�e,��	+�.���sI������s��~��E�-y�\A	mFM�����M��&�vn�}I�w����r൥�]U���{��.�"R�HO���兔���S��r��&��/m�0�e'y���;�<0�<�I��VW���$F�,��!���^��F͙N|�̶�.���o���s��&�ϙ���M PjH���B;�������cpl���U�;�*�����tfͩjn�U��ڗ@F���{D�AW��#$���o�$F*���Pi9r^�.�=�	/��u?���{��qZ�o�s5_޸�}�fh��#�
yߦ}� ��Nt�Zs]���4�,�u_A�:�hR�'�j8����<��.�c�l 

�¶m�ͥ�T7N [0�cE�GU��UV�ќ����d(~APl�l�Oc79�f�rp~27�����m?p�������z,����sة���xʽ5�n�ߴ��	�2�0��砽�(��ʐ-�V�� ����޽`b��;�])�z~drhh(cWW���K[��k�'�p���g��;n[�N�w0� �'UpO�����ĕ��W���d��^f�Iwn���+������ey�����z
��w�n^�bK�r�s�"���W�B��x�'}Rٳ�&��/�(�}��t'���4)���Qg)ה�P�ѷ&��������Y��Qzڨ�ٿ����j�O/xy��Q܈��(�Y0��ݠݚqW�y�j4R��6_��2-���3v �9;{C��|ܯx˙��������{Ny��x��6&��:5�A�;�w��?o�lu�V�Rb����P�����M�Gwg���:�r��u�fy���S5Dh�J��E�m����o 1 %󺙏�h�G/)m�l���#�]f�<4���[�G
�Q�ڑrMe��<FNe���Ĝnx�>��^{�d,wz���W���UĘE{����f�7�߯d2)�4�����Uv�Q��h�1E<�a����W�	�[~Y�=L1�}m:WB�H=�+��%#�ss�S�)w���[����m}�<yl����`��[ie&�0O}Uzq@w�f�SCWdсc1�k��*b3�n�S[
�^��P�Rz�Jfǲ&".�Tȷ�Y�B]��f�f�Q�,�bhRM��o䋙ἤ_��n�o =!�R ����MAb�
$��0r����? 9����<Cwg�+7+�2ԥ�GɵF�׾Yvηb��#�Ut���dk%*?;��k2i���JE��d�=����S�[�\�v�;c��N�%/��V\,<�Ҳ��< �߾�m����2�ڶ�Z���kɐ�^&ܬ8��]~hχMXG�hL���W��ߩ�@xZ������Ϟ�����Px������BKR$�U@�~/�`]��Û�$e9b`����d�25e�&�L
Ƃ�Xh�����3�_(P���u��,_%�d���i'�M�k��RP��:��DS�����툰Pb����ßO�8�iv�䃻��M>_$*��5�_)͍9	NW{W�[iox�G�7KEZ��=ܡCo�
2H�����ޜ 0x/�tϯd��(1:������d+(�A��f�e��
x����L��m�ܳy��D���������0P?wn:<��c�r�Sc�.lr��=]�.b�M���Mϻ3""`%�>"p�&�f�F��nR�<�k����*V��ms���>��\L�ܑ6�n��p�gR��*�G|K�aJ�����;X�}���K��#���M��<gY:h��v�2%Z�T�#vgE��٭��k �t:��;�_䖑g�4�9:�����n��q�C�U�v�;X֬�!:��r��JD�~�l6K����kF��V�^u����T��B��F,Ssh�3�-�YT����/~��ސ��"m�=���w�a�ڣ֬��Yc�Z>�� ��}�r0��L������J^���)C)�s�_�r��Զ��p'1QX%�!��)QR�2�Fޫ�E��Z��$b�1��W�t�E.�"��=�(��[o���@ �%�p�a]E��̫l�m]��I�T��]����O�Sx]d [��x�b�>�JP�"��h��tP?���1Ҧ��lE^��(����o5*�~�&���w�m��m��0)�E\1�}$K��C��#(u����J����gd)��;p~�t
ٹV>|�#�����=g��$0�,��#l�z?�㒝�նb�������(Sz׻�'�����˂r�\/����LH�0�����=9��]�aO�/��tn�J6|O�׳�"`C���KF-��M��|e����5��]��	������1?�]qD��iTu����S���?��@%<���x�m�%~�bB���-��Z*��	��^�s�د�f���m�m7���=Y|���h�׵I�4�7�ѥE�H��aR��f�*$b�������Nv�-��3y�`S�AD���/i#��S�����\��w�3E�pj
����Qæ}y��NN��d���Zz�~��ސ�߼�wې'�j{cV-F�c�O�mX��o6�?iw���k�:P@#��d��1��۴�
�m�x�>$J�-�Z^52S�ߵf�-�P�ճ��D����������cUx�6�k�K�+/�t�d��W�:�^':�{�j6�>���v2�;�x:��
DԪ}.�M�y�@�:�QQ�����Vtmv�w�e���л��}�=�5��R�����9dS�������IEj�d?p��w�=�cQ#���gW�k�4�;���[��ƽ�%E�or�[�k�K[�.&����{��ҵ�H{���������ly2�k�(dv���	JKC�����]j�k,ң��պ���X�,�hH���������̓�mz'�t㹮=�`k�����|:N�|r>�C����7 %3�z����{�QT��T��w�O[W� �ڰ������R=����(9���§�M�DK(a��h�qZ�A�����	@hL����vd���Vћ�ƛ&b�0����>��'zbh�K(���s���Et�m"�ɨ��կ�QJ���XsZ�_w��-j�O��'k�e'�ss��ÜQhC��O�'���}D�A�@-|���K���ڸ^�>����	�o<W�n;�7i�|�5�'_3J�>��.`�9����yL��uL�B�{�RlB�s$�@b+����NNZ�� 2db�qJ쀯���ƃ���	� x�+q�>`4�{��ǡ�%m���C��/;8�_�G�]aE^�t��ж����]ܮ��w���������+���#8��P֣�/O�����{��\D6@u�bꕖPmd��q�%�����S�}��)*@�0#G�4:� OQ�:9��ν�b�Z/
i��<f�����!����m�+��Q����}~�)�ci���ޠ�l�Ԁ��!f/�X���"�A������X==[j�`7&�DW�<�4�ֿ�C`ߚ_�錴vi��k��̱��/4Ɨ��^H0 �ҢR8~��Z���"q9gr?4,?>�Z�E��aF.�L� G�ILKo���y3Ju�f9)o�+T�`̊F{�jJ�<|H���C�~jK寂kT�^��<b��}���h�q�^0MrA��<�)����M�@`2����f#�^����¸�$�����$3���:3xZ.}���ͳ�юvM�ƕ.�M-���w+���� d�C��܎�zp�~9Z�e��dR%�E֙5
�D	@9K�eib��｜����'����{e��]-&�R�X�6j8�RƎ��Q����^=M���s��O����"��m�rE���Y�#^pc�h�h��D=Zo���MQ��4��x�A��'o�_>BN�(�:G���0-��߽-�.�뢚_R_�ܝ���z`��9>�Պ����>&U�n�>��(����;�q��-20Pt���x��w9�Z0qN ~��N���u@�7�����Q��<�>��3�f��yHF\w��%Ә(�,o��R,��b�E��)�e �@�5�TB��:ne�B��j`nC��_�q����5�^4��M����GͶ|җ�֧\��'��j�U�2#��%��3�<�;]'O�BL�ڟ�O@+*h�p��II �$�n]9���{�eU.*�O�^9;漬V?K��=�2~��"�����d�RTf1M�����tJ��G�6o����^2D�;��ⷼ���_;u�B�d�s��%D�e� �G�U����t�F����?�˨�'9����΃�S�t���O41���c�<�ڈ�7N
�R����Q�u@S�}��������y���[�:�~�#V
����N�@�lK)f{M�6',p��,_����+�+�ƚ�'G�h���K]�8����(3��j�9�`�_`��ޢ�0�,,�{�<����h2��K�&[}���m����v�s�)���>��?ε,�\Ze�>U{hV.a�B�c~3�� �I����]kXw�Kw4��Z~.�F�t���[���?��ޒ��bC��:_&c1��������M��J�����4&z���^�Geń�x0���\��@0�y�66i�,i��SQ%�r.�子&�p��/o���ר��{G�����s�i���o\�<����\"�˅{Bj,7<�-����h]�B{���C$R�+`>�¶���{ ��8���^��引�K��ׂЭ�ߊ=;"�w��������#���o�d[nu_Qm�Tw����T�*�Z�Y�
F�b��]�l*,�jx����=N<�ѣl��KLQ��SNNR^��<H?}2�UJ�5Y��?�������5��PO<̐}�dS�@g��6��E%���E�q�@��1踠�uFS�	��DϘg����5�r1c|��/;a��1�e�T�x٨�/c[k.��f���U��7b։�3��̏���G�R=���KM�(1�H̺p�b�w͋�����QCn!�d�@O���3h0�x¤�EǠ��&+>�&�Qlr	���Fe���lWa��Lֲ�P��{�>�B\�M��bBrmUD���_����"d�#g�{�q-?Fy���������	�+|D���,�l<�A3q���<���lz����T��X��2~�����f&e��P8Ru8�z7!q+֝M��,�	跼+��gn�^"Ϋ���?�ژm��Z�?��t:,ifp!����`�4�5��A��~�IpRY�߷��j�"��7���������O��;�Ӻ|(L��ė��%���nTS��,CGe'(Pz��)�YK�k���Td媳�ڏ�Y��N������i��wr���~R�ֵ(d0?��_Zs^��9���Y�/uk�q&梁��ż��nv��b�te:�7/�NH��a-l���sssOn��D�`U�8�/M�
1��S���;��#sqE��m��8$���M��G�B_}'���~�a�u�8�iq����I�nG-�{��qttR��7׉6��Z��a�_ �,���+8j��K}�8H���'/��O���}äs��sW/�l�O��5˱�݊�2T3�^U�o��,9bD^�j1W7�������@=H<#X����f����=�"Os*�K�'צ����� �����Oacn<���ṅ��,A�����jq���O�wd_�����7�觿X��"VE/��lufOl`b?D�����酡ܞ˶�����e?�?7 �͒���w}_�E3Mv�Ǹ���i�!��_��/��جt�Wԏ�*y�|OЩ\8�D�[�6o��o��'��B�b�_�:����p��B�nBL��Y�/R`;}W쇹��#1�I���_ѷ�7� _��s5����u��x�CT��B7����#���o��0���2ҽn�t����M+�|.ݽ>LL����h������r�����F��gF2As�-�
��Ʊ%���=�۶����+7+�s� ��M� nЖ���Y 5Yx���7���}�%�y,�b�l?�{����L��d��Gc5����=L�b���h��v3O��L�`��)���;��a/8_�y�\R뼵��_j��tk))LJ��i�{�	�>=*�\���غ[�%������-��(�>���pm�s�0�����%x4�7M����z�����b�2'kĚi�3����7����z"���I��#���d,ҋ'�|��5��D�ZZ�u5�� �{���q܍��Qw=o]�F��^�h����B� �}F�1s�c��ToUlK��^"����^�ǩ�������o���^$2��T�[�#����,nZC`��ѣU���mOE"*�9���wd1&V{����%���Q~T]c��8�Mª�('��=���]A��7��H�.-���������JQ��I���M��QM�"q
�no�X:F?�Q����/��{0��=?��-	\�Ab$YM�V	���^oN�'E��7�g�d��}I��f�������:��I��3Zil���S��\���[ 6�>�]��?���Ay.~�����[�*.i�)����>E�sM=�=�"Ke���gzi����j4�<3����$u��AD|�����j.z3 �#��Kg���8�:��d��{v�C�v�mcF��v2�/�0��˾�1�d~4�2�N;�����el���G�Q��c���r��Ͳ���y�$l��_�)ז=�i�~8�5�
��/�� ���ȦcJ�9�T��w�';����e�ͷ�$!ϵ#צ�9�1��KM"�iN7�YZ�a�V3>���U�mݽ;?C��?�x,,����M����3@�r+=(��;��-LSJ�L���#���7�ۑ6i��I!/��>�Gi/�j*�ҿ����bk�F�n����W������g׫yq��?mrA��T����y��P���rCb0����}Er����5t�9�	�:RD�R�@FL
�W���tA��]j`�sO,���]�F)�A/��]#��bDq�w�>��<B�.�cI���Wu��ݘ��x��ȗ�5��� Ts���%~�p.��eޚ���!��0��]N����^�c����\H�b���p�q�g#넍3���?z5����\�^=� 8D;g}/�x�mf�=zWAy��N��~���3Z%d��Q8ǃ��
�ZV��
t��
�����>������a8mp���]E���_	$��B�AM�^g���E&�10���jW������`~$��<IH�6�l�ٶA��{��_#O��?�#�E�F�8���8'���7f]��A�:'��Q��][�g�ƕ���?��nv&���{�^�x�X*�=� |ʟ�<\K�����_sAH-j�|���N�ֻt�yc�f+�XǸ�CH�]�Xw ��fK�yx]qR��G��φU�Oq��SRGj�>���wV�,g�y,[����w��*���ZI�U�`�K<����K�P�vV�9�TM�U}HY��6���7b%��Fq<��pSͬ��gxw����̞!����w�Z�O[�4��|Ѵ~p�����������}��$��5ȿ������h������Z��C�d�6�\3��z�>�O���٨8A�F��U��&�����ѡ`�J]�&�� 4�$���\�N�zoR�UU�	�Z���I�L*}�5"�x�}�Ӷz��1Li_�ќ����7�HD��P Q$�jv��~��j�pV�L�|{���c ���W�I??��T�ۚ��P-���M�=�O���!\���S��ʛQ���s��0�9� d���ydF1����,&)R�ϻ_\������}���_n4/
>���̖H�t'a����<*O�M,�R��ڲ�Q��8��9���ɐI�"�"���v�¢Oh��8!d��w7��H�0�����.NK�����9*5�0c�rb|�pO�D�AV���6�Wd�LD�Mt�
�ӏ����M}��Jd�P�=i�v�R��<�lu�sﻬ$hdN�K}����:�B0%�<>��/��E�UD-ɥ���������8�5�/�D��Hش������v�e{��{�
'b����j�m�9�~H�8}����*�*-��qR�x�3�.�;[7�<�a�~Y�T'd#�ԑ3m�s߶6'��3U��s?�Ts����e^Q���~w4v1k,�f{ Q�$�����ɏWMG��	���jO�����*���h
Op� f���J*�����r�_�W�(%����q ߪ�7�=|�2�Ӂ{c�rD��t4�YdcF�u�O�0P���(�8w��n^|��3)���Z#2'�5J~
�0<֭t�����V�m���mމGzlI�M3���j�@����`1,b���v���(J6��P/,�댄�a���;L%o9[Ju�d@��%�Ȁo�uI�&s_}y�] ���9d���aTU��9ϥT��>0��Id��j�3��^���&K+>�����"r��J�����l��U�F�7N�֡Z���f��Q �G/�j��c_��N����������s�|ا^��cT����"?�<I�Y�E`��cO��!Ů��2���{�J����E����@w��W�N�1#�:!��
҆'�d���bB�M�f���pY�e6�9��#
i���@^M���-��*�Έ�K!`N�VE���/b�8�B�kj�����֨2��#-�����c��\P��O�h1"�g�~�֤�qөP����NI <3>�p�^@ʹ�3��gt4�=�B9-6���7ٮ�
]��)��j�z8�\�hK-�7�jp[�+��z�����:C�N�fEA�ٴ�q���X�����ܿ]��|�W��wc���T�'{��z[���IG�H���uOU�Cެ^?~�;H�X�X�z�*�e/̌$����Ÿ�E�Qv\�2"���V�F��2e��cK�\D�$�Օ����Mz�Z��l�TdW�B�\ū�e�v��כ��$��yLU����9���(��������5q�̓�+.#PKj8m �I����.v����jЧ� V�@���G$�D�����҄H\��	�Z6��9yN-��l^���]�bG�F�B &��O&b�'����L»�e�kU�L7hhHc����sW�����,��-^���j�����h�uF�'}���f���Q�k��l�wgO��W,����I�a���m�3�&tQ=11ڛ���?@����w���V53o�\� e��5lǥ悏�K��i�tde*�N���T��,~���$nb��;�n#Mw�R}��'D!��7��{V4;�2t�*z:,��@j>�D�a�YI��C��짬�c�;�Q]�Z��%CE��g۩&}��Ǜ&���I��eC�֊��.�N3���h�$C�>F?K�F&�����*�����XY?�>3n|���S�~�s#~�<3��fk���|�m��z�[z�J���b9�a+?���$��V$o|An�y�.��^�ힲ���3��;p1�wp?����G����{�L��X�x4N�u��q4�o�?����Gj�}�t�Np[�<@�[����f�'Y�]AS�C���/c�v�HH�����a"�,�5z$��p�7$��K/����a{����[�V��$iR]X�e���읋P¿��,7�ԕ���ʧm��W&�|.�V������*~!����o̫��o�������ם��S������KW�I}���'�s���JgR�s�f�$�Ӿ�^p9�#?���DR�p���g�g����,�,[��݌�XI���h@�1���o�L�->K�dBkO�c5��^>i���YU^nU��ͪ��s_]�
���I�jh ��S3����mV��k���$:U_\λ�A��m2 9>����h�"_f�Z���H�'�����R{���8��'Pc���W�Yz#8���~��e�����8>�,\����ʒ���c;��J[�K����B��b�cE�|p�X�'k�p,��� �ε�27b2���S��^i�P�m�|�}��� D{����~D����}�f��7h�[2Ǻ����o<V)q9dW:E����,�1��XRi����{�ֈ��%]�?365�$.q��p�ߤ'܁�rd���!�<֛q��>M;��&��?/D_�IJ�"��g���{��\�� ^���U.R�_3|K*t�<"�>Y֕tH.Rs��P��3��[�?�V�1P�b�̚�q�@���OzT	��rH籱�R�0��[���Afoo���(�	*IĤg�놉MS�D�o���ǹ5��[��0[8���J�&�hF�f��Og'��E��I�2Tpio���S��}B�{���|����\/N��Ib����C� �S�0�38::��/:a�k��3kTf�fs*y��Ze
����m�],a�Rr��HV:��_��� ?]ز�����\wI��<y��r������)(<�h�7��lK������'_b~J\�V�y��L�8h;C�Dl�o+Q�'�	��Z{j���¢U��jDm'SN�Э�����K^�:&8�$�\��q�w��+ �k b.06s��|��_�B��_5A
Pi��/�	�ޟ�4�z���sΓ�S\�l|X`�#��ŭ�}RX�_(@um~'�:\_��d'0�+�`a=����� �z\~ٯw�"V_�7����ٞ�JÙ�?(��O���A1�s��e���|߯Ƶ�R�uS���$�r/��@f�Ag'�Ep�ì�A�$��d�|�b�q��|�o��Ywbh>ֲ�[=9e=lh=>�`����z����nD����N��D�
@'6Dձ2���-��?���z��Dv짟�\��G`��b)��wD�>����Z#���Y��$���#'1�VŤ�rɝrb�6�[�ԼnUͦ��a^��z�mg�iȻ`�z�գIMBWq�p�xc�N��5-�j�����7��uj���C9m�Ҿ`�)�~�����T�4t��Ħ������#��V��a��tӍ'����~�+%�mҔ�&���FK4�6O`7���Q��"���J��A-�	p6�ϨaO�R��{�`uK��V�,����t�w^�D�UN�����^tܼ�S�۹G�b9��b��Ղ���|�+�K��?+xs���yr�}va��u�+�([	�k;���l8 ���O�I�+J�j���w|D�{ǪF�:��hU2���*�1�LF1*\�I*��$&��l�m�A��;���j	s��/�o���m��~\�ZmXT;�����-��~4��S�Ac$̗�Ay�>�Yr��ˌ�.K���ջ���\���/�x^3����_���њĝ��7_,�Y������ ֭������)߉��Z����z-v�Z�3.Iq�+j�J@d��nhzl���m�C!sX��`hz⌅/!�̮"7[m�K��Ȯ��Ei!��E߸���B����̀b\v�D"�,�WE�l�D��B?�(���;A�.�%8�`ae1����rc_:hHm��0Fˡ�ݐ��uY��5�f�NͿ2T��5c�M0F�^�~�M3�׆�
�,v��3Z��T��׳���EC���,� ��`z��
�O4�.O������7U�k���6��]��&�n�J����JM_�ϝ�i����6�wm�t}��^�y���>�,n��ɯy�;7���_�9����ɏ�u[��޽o}��)C�	��(p��|�d��`���34�����`���_N����o�������)�	 PK   �i;Yh`Pҷ!  �!  /   images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.png�!MމPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  !?IDATx��}	��u�WK���hF�h4Z@�b��-˖B�b�����!���'�|b�CVs�3�q�#�lr�y/��`�1D�%����/�e$�F��=�VU�������Qk�A�{��U�]]]}����:.�<��c���7��;�a,�4�֭å��>M����O�Υ��KHQ�O���3)2�d��<���*g��{��y�>��2� 1-�C,χI�!z�����P	"�?RTbA��C��Œ��_�I��T�j<��0z�J�W72� ��O�Ua=QQ4?,����,�2>m!6��+����I�Z�U�����˲�	����?H��������'��@�jڿ9>�Ĵ��ʊQ*KFS��ea,�z������S<��2@!:�
j�Ytʍ�sc�O6wT�8҈�=�����{��8��w�}�V�2b�ب�L�"룐�,T�D0sb��zz�a(��.�sF���0�O(�	����a*k�p˵;K��_�#m�p����%�>Ҍ����6l؀]�v�RK.@�	���^ȅ�{�8_g֬Y�����&�Ju,�����'�Pۉp Ο�Ce^�Ч�9O�8?����ޡ�q��Ӓ�Qۅu��8':k��D=v7kN!P�J%C�6mb�e/HL*���7sRKe3��Y'��(�?�>�����T,���� �($S��,G���0�
Ź�|O�f d	'�?�"��_Ob�V*g0�&��Ϝ�_���p���~\<a��P��J���\��s���`�ԩ�6m��p���25�J������J�ta��J2��aZi�[� �<����{��r���`���l�[6`F��d_��-i
��G��3O�dP�rr�0u�g�����#�����CKKr�V������{0g��~��={6�� 
_��לƲ�0�B�Gɘ� +c#�nҫ)�Qt
�BTL�Bl��^�}w���ߢ�M
��(����AX����F��Ə���?�#Y�h���_<����
��u�~l!NuO��-r�*ʭepp[�n��/��H$�Wǎ�թ�\�w�u�~?���Ĩs;�r|E����� ���̙x�n������R�H��5�� z��T*����X���<��f����z��o�rV�L7ӛpk`�4f2��P+�4���F�{t��%е�[���R�r�-hjj�������9��c�p�B�}��B��d2�3UU��x
�3EX���gnGyh�H�@��l�@״��9L��_5|5���~J7��`
,�m*�<F��p R���6Q�lW���?��0�e����V� �\C�]�C����e��?0Ps����lm^�#�3�A�Ȍ��c}���=�Hs����җ��G}###�����g?�Ypu��X�-���"�=p� ��������9S���g�٧$P)�l��L`%h�P��f	��T� +.ML�moJ�+���
������
v��?1o
���*�����9���>2sC��� Fq(��"��`km���N|��8�<��OÄ́	¼744�֫7�,��������/�; s��E}}}�E�)�[o�%.굉�����+pݜb�b�޴�����B�@+[Fe1_�� H�l`V �L@<L��Ҧ*�Ӡc`J`$8��a�#̚9���yG�4b�e��B?kH������5}��ս8֚ru4�|�0Ϙ1#�����+��k�axx�� a����ǜ �������wމISf ��:�rS'����]aY�c�����V~��	f�6	�������	n��l�ထ�6n����[���SP�����ί�gYqGl��aa�Pp��Z���F���}������w�^9r_���l�2����"R=x��R^^�q��Lm޼Y����_��{()�ƒ�q��(���Ri��[�Į�EЫ>*�QP�M�'�$s bf1$�\yؑa�4 �!�4;0��B������S�V}3���`��F��(���n��=�u���������ß����o|����׾�5a���M?��$/ �E�>�o/����֮�]�E�<�:��ZrH�"����K(X�M�^�Zx��"&��4� �ad\�F�������L���$`�ۄ�?���V�y(%Ka���n�s��(ߒ�?�'�o6��܇��	qW�x��c�쫈$T޷��$P ^vp4�g����R��@	V\}�S�b�*�L  iE�G�j>N/)�����61�$lP���<�ʹ�N.S�M�O��bbQd���(A�p�!��撏�
�ޗ�;|-Ä�(�������W��+�濵�[innơC��`��Q��9�-M��ٳ�[c�e`�h�Y��#���]�l�"�$����$lF\�ZV��0�I�[�,v�6�
�P�;�c:b˄����F�X��Ӡ(�������Cs���>i�l�H!
�� 1===b��;j����H&R�1%6 �(���u��SE�D�C¦��5b���������c
�i�d���d�b�1%%�c>	$��F��$��$"1�|O.P�ML�H�Ϡ��M�)V�p$��][����,�%S�� B$x%t����M��`�hE�#��φs3�x��J� �k�!��}���|Zd�x@������yhi��h[4��%�1�����,A�����gP��Pb�x���iX�������b��lSŬP<@(�o��EJD�
�D���1%��S�����gkºoi�J���p�����?+�Ԫ��do�j`2�q39o�3�n��	0"H��'0�b��
��*%�!v��43k�d����
=��!|�/k���I���)g�km���S+ېH���H�+�uSX�x=���]��~�6+>LbH��a�l�v ղ�!@�����]"[[�O�X���nJvc�!n���n�h�9�����F$�D�3o�2���5Č�t�F�]	���e�Xb�1�aa�C���5�UQ�rE��e����>E�f�T,�~m�q�昿�?�+���3�7ǦK�`�[�������D��:�W�a�>�`xDT~r������}'+2��$�͗Б�8f�Xn?Yq�{xu�d��|�no^\���rP�(0�T�kn������}<�z1m�a�
Q�#�|��TBWC����K���KM��**K���q���'y�-k�܉�o���p��ĵ�Y��"3������v�n�d�`f�0CVj��+�u��N�VةϝvS�eN'����ἀ�^t��V:�s��8\/E�z�"�u��%o�ʦ^�������N�ZD`��NW/Y������k��`�	�����B�Ǎ��D�j	92r≎+ ��d3���긏���t}F�3�J�M6]
���	��:����͹. �����q��3�����
	3�`�A���zi��Ӷ���f��n��t��k��wh��U��~��e~�Su���/�>��z��,���F�N�5ı�wlv�0m�A�T͓ܠ\c�e��X�M�e��d��U�j�Xr3R�fȶ�e	W�/�[V�j^͉ɫ5��}{9��d�SU�,�(��`G�+���Xr�{9���-���v�_���ӧA-�V�<
��U�����z�M�q�&h��K@�@\�QU�����f�.�h�꒶���Z���ŗ	
}��fd�H�-EqYb�Ĥke�b�zI *�@t�M�% �t���3E쨧��O�߸��pDTLF= 8-����Ǔ]���?�2�%�m��R٩��Ldd�b	��T �!.�&�c��R���2�"�F>q*%=� b���b_-����.��Xܜ�:zز����5�-�"���z�\١.�z����4ؙ��a��M%&� 9[ٿL	L�2����Y<u�<Ҁ��m�t��<S��qkq�� 1�WZ��zYU�\D����.D �N�oM�܍����x�E�= �C�a�j��U��r}e�Z z0d�zE0r����L�^4	�5t��N��v�39�K�+Ki[/MT�ws��N[@��"�[P�r_��$��}���i��fk)���e�V�[_�1[z�NG���%f&+�N�1RĒy���]+�֨���J0 %�d�ntLUڡ�b܅.ƃ|Н>,����O�أp�{�;����֍��hZ%��&i��+S�+-��CG�ME%�Q���ȮG
��W+ǧ�f��IT�R'��$�O��?�&Z�_�宴/J������so�@=a�"���r�-�=k&��&��*'��}-BQ�Q���Ng����������&����M�윬����E��o�q�x^�	�v뙛&f�ˎ�҉����~����f���^aw��s=�WH�0 ����'�R5���8/�e� �C�����J)�)v:;�Ap=��:˭PLGY<|@!("r�"L~*{���sv��ny*~���:fHE��t��\�Q���S�4�>�BQCp+u3���H
M�!��" �.�3/��$d�D�{Ve-��!>'ʂ7�R�""�N3F��(9:�Hl|��e�����${԰�!��NH4ݮ'Q�]uR������[r��-�)��[i �¢�����d�i��+�t13�i�]��t�1�("r1īC�)s�In�2C��T8��a��LCދ"J�p	Q w��O��MgLKw�v ��&\թw)�y�[5bOn�U(Fy ��(�4��$]m"���b�Ʌ���cTF��V6YG�]~�͸f*#����""�.9Ə���Ԡ=(˔I9�N����{C^˰���WVS����;m��G(��*�<-�(��p#�]H��kY�#(6Q��(�TQb6���D<Rw�.��I�~v�9v����kKrx�����h=d�\A�423u�"\�۬G{���fQ�Q>���~$X��I���p&P��C�g�H�F<ڮJ����)�#J�o�$���L����R�(p��r��m���z���l=�v�El�ퟏ�.���p��;G�=������&�趙�F��mU��tB|��r�����Va‡�`��<f���Y2����&�ɹ����u[�ܜq]�#�${��\4[��|�L����X�yݖX'M���V¡��Z���~����>�v�J@�R�hȜ�QN#hDx�~���S.K~�$��OF��H�{/���ȏ�!h����S��@1u�3�i�L>E�#�H�ά��WH���9Ч��~"�����T>��<�D2���S(��T4[c�b�"wRM����vtH��~%�[�D��Uo����idɒh�I�Lj��Y�ODt��6L�o��N�9��?��^"�_P�MeQ��s�a��J��-�$��&J2��j́�b
s�MXv��ZQ��8fKSya<A��{fvu}?�~��z2��"KF�*A@��"�%s���f�)�5���<�� ]���/�IC~�	8r/?p�&T����0���:݌��K�,���ò(a���-bG?��(��RAgOr��gZ_�;3��n��^��Yb��H!�����3Y�I��Єi�O���+�`w@��y�x;�c�Xa�a��x��*�����cO�
��k�+�\�����8���������I[��f�Gd�S4]҉3j�`���y�������|*v��w�m2���Q��#q��C�x�~$��^�aH�c��0��M��j�H�o����R�x#*Q	����"5���YVh ��ޖ��I5�o`d;x��p[3���&]٦K)I��WÌ� [��O�	��J���h뙆�-ܦ~l,�'�$��d-n$F�ⲥ8��4}Z�9�~Y�%#*^9N��U��H �M�^������X�-�`�ѥt|4�U���R3p(�i,,ya4K�ܤ��T�[q��[R��
�V�$��EU}v��qŶT&�=�]C5bպ|2�Dʼj���M����$����+>؇���jε�rƓ�����`�$�I��X�:3#���dO=���GN}l�>& <~��SvG�A��P�r��>U�%�+Ἣ�t�M��
��>Y���~���T6�ALۮ�e5���Φkؚ�'�k�_�<���#?�t�`T4.��Ay1�c3R��3|r)#�/$;4ME4����CCMC��8�5���-W�+)<�J/ΐ/z��L%G�[��~Bt?�d���2s���3z�0W�nf�^�gxVe~�B4���i��_���2�{
\�ȂO7��π�)��!s�l��|��\9{���\Bb��Ǔ^��$�1rL0#͊���|㇧�u`�lnb*�b�_Xi/��W? �ɟ��դ��Q0(��.��ߌ�Y��+����"�T� �G$�_�����(��?���;�8"�^YY!th@�� ���o�.���;@���w>��ddX�RN�|xb���Ce�����)}"�Z��[���&�wx8���t᾿8�^�u7�Ry^�����Ւ%K�q�F�`b���IL󋵫(ʊ�&$��S?��-z��7,�M�f�K�}�����ja�L]������y}�,��d���_��=�"�����;g�]�`^z��&M��իW�W^�q������}��u�ҋθb���81ԃ�is��.;��[3f�&ḫ��t ٿ��a�_��0T���|����GĢ`���Xw�5q�Z ,/ ���%�(⭷ފ'N��^Y�?h�����3R9�,�٤b����iW#PYw�q!�$�y^D�F<�����N^�������* ��9��}�D�y1I֙wAIg��|��Çg,L̨�z�>� �}�Ylݺ����� �������r��%A�}H-J&�B��6" ���+�2Qpɡ]0�����������$�������ʸ�������^��1W���O��{7y�Ռ�=*V�v��M|��p�u�aӦMhiiAdd/�
莖��?Q1���^w�(v�o����]�U�k@�j�����'pD�y�~.�Tt�����<Y�%��)Y  m�|>�����/�CQ�����X�{�ʕ�o�C���F��;Ώ!L��_��W3Pv|�ҥK�x�bqq^�o2*Ƕ����4DWռky:�p]-@�r"�Փ)T���[�d���ȳ��e�Ć�#�G>"*�Γ��c:����/$���6a۱e���V���P>/�̫l3�׽e0����j�cɘa/3䩧��}��'~��qH������`O!��{ёX����Q�wg�O�0f".�_"�'�B�W�fb_I%��W�z/���Y!�=��L%a�/c�`$"��\����(5}����#����q��A,�U]�s����\/+��'0:::��}c���y�Ν;��ى;�MMM�B-?�c-�;���|3�o��!���9⌋���c=g�m��<��C���'��|A
�|�39�����Sܒ���c%MzxLڗ�!X�Ӯ�L���y�'	+������m��^�X2�P�����Rb�Z�[�l)��}6)(1lmm����E�6}�t��B���3-�j=n����(1*�/Dέ+u8A!�@�<V�0/jƹp&���y.�������=���b���DL����_W�� 4u�Ykl�'08R娴 ��ɁJΡ�l�����K���~�m��~1,	���V��LG����(�9�`��1�uK���aC'��v�?��%�F��܀�X�{��W�O��8|�E�r�N�X���r��*V5�����(����2��xy�D>��+<H�?HS6@�b������F0o)��Zk��7��zWW�w���W��e�������U�V����?Et}(�3^���{�?�)�f4��Ť�h��
��O?�@� �����&F[�Dno�ɞ��QZ�`�J��)J���Əo�����RJ����.��vG�|��$�!Z��CK�)�{�^�Ϗ�	�%�?BZhT���|¡��vv h�"F�<3cjK�T_[�%+c�&tM΄�\r�!z��֭[�K)��B���5E���Du$�
<���ϕ��<)���2R�5���m��Z*���s1ip�0m�項�>zwG(�����F�wM���_�� ( ^QCyz�_�:܏�s�GI���˿s�E!/O�9�J}VGʭ�RAʦ$E�c ��2B���P�$ :)�kD8L�%��;фCgk��hau�@Xt5�H�~�}oL��5R��Q�N9D�����O�	$Y�t��	E�`��E�o��R�]�<���p�]� ^�Z�V�yoϓsb���gw��=vƫ�[@
���6�y��C��&E@ƙ�0Ǽ���b�    IEND�B`�PK   �i;Ym_D�� �� /   images/51bdce1f-f35a-4993-9bab-5f201461b496.png @鿉PNG

   IHDR  �  Y   "���   sRGB ���    IDATx^����e�u%�o~�bWun�@�HA` H0��H������xy������`��Y���(�%J�AjH�@�� Rt��+�t�����^�n��.���}�~ᜳ���|ASNں��	&E�i�"�tP�.m�q��&��
�2Ĥ����[������yY�mZ �}�ڶE�O�?���A���?@�^�u�����iZ��'Ŀ�6@�� ���0Dh~�6�
�4 � ������\ش�D-�d?�C�]��
�A��x]�?/l�t~?�e��ދwǿ���?�w���;�Оݮ�>B^YW@Ӕ��������}7z�E�_{os�ݯ��a�{������ҿ��hN���{{D?7|k��5���-��Kγ}Þ̭��ﴍ�m�uԠ��[Y|L��&�3�+�w�eQj����U��k�^7n��~܆h�\м�6l��7�+�m�u�'5du�u� �����u��l/�w�S����9�_���d�>��?��m������h��nm�6-��C� nn�%���7[3W����q�4�W�Z��8*v-޻m� ����e��q�nm�\�#�cݣ�
3$��-���w���a~;
�s�b���ϴ�zC4Q������N��k��9Q�몪Q���'ך�M�r=�ys&����6"�g�ƭ���}5��ʱky��~�q�A����B��~��:�pv�Fi�a����	-����z^4D��p[�}�v���o�k["׀�'��m~!�����"DQ�{n�U] �a�j�rL�>�s�SYV���[33ݵ�(�j4���=f�5[�·q[{~x�4��n�i��>���О��\��]Z�`?���֚�љ�������Z۳K�%?w|F�k�S��uQA�Ɯ{A�����ë��,j̳�md����0 �I�8@���ss�!�5���2��ՙ��p�G6�&��Y>�ۈ�ܽ6_�\'3�5Aۺr��5A�R9��1��ikp�E�l��8E�5�{�H4�fC���+[�f����0�ic9�������6"�b��M[h9�M��M��̖��Y���{�u�֣�?�_|o�pQA�%[��D� �E��o|�8�w��uq��5S���!I���)Cń�k�{�/����,��dk�W�\l�G~����1�pC��1�{�z��k����;�J�����G�N},���{Դ!�-T�-��G�C=�l~w"n���6�ږ�[��|Έ��~����~vǓ�-�"�'�[��],��p�U��p�qgv�����b�]�Gq�Ɯ�T�>Ӻ�6��|��=��<U�a�"f�B�K�>���l�-��xW�ѽ����	Ѻ�|��7��c2�*�4����f��W�rwO�_��"4am�=ȵX"jKĨ�cnkLf�����o�Xk7l|`�YǼ�I���Z���`����L�yM�!�:��{� f1&�#�MČ�I �=W�0��8�w�.`����8������� ��*�Q"�1N]X�3/�ęW�71����	1�
L�y��q��q3+ps��:b��(��m�*𤡡�]@�4�mY@E ��Z@�� ��₡Ñ��Ԝ�1n/l�
�D�wZ���u\ �E����\M
 �lsו,%"����������َ��-d����!3T���j�3+PPİ�y����,(��e�.s���h����lЮo���?l�R���]`�����{:s��®Z5�L��ؾ.�lQ�rp.܀984Q:D3��fp)4�\A����6��R�$�,pS�)i�$��s�����;I��9 �n�hfks^�[��@�g�P��ܬ�'A7����E�����n�(t3j��U?�ygK��/�:�q�@���$n� ̯�ȁ���lɿ�<������\���߻�psk׭���f�ޓ�f���]��e䜖�LD���]�9s:<�XI?vČ��%�O�F;d�w�uE�c�-�#���5�L974�g9p�CG�uG{f`Г��m��Fw�@J+�����St�fc-�$�@������9�=8xz��5ϭ�����^��7[+;�n�h����D��@Gv������q�������r��{Q�N;N�D0�cUi�;�S�2/��� ��XOPq���EM�"�d6i7`�]ʀ�f��� ��Irɓ�֩_��� �1�-c�H{Q�����o�"�V��$�|�[������d�AD�&`0��#�Eߚ�o:"I���<Z0����n����Tx"�|��ܶ�V��$fi��BA����Q,��<�k@�'�8n>`�����E�]�{y0Fh6���8��0�O~�no��k4q�g��pu�� ��?��jm����F�1����^O�ПTh�PD�=M2�`���#�I�+�rĀ{���|�fI䀑Ɯ�����W�������M�R	p��kx��{���M�Ua��j�� {;��+��ޟ�~r�����v��|o��;8ļkٍ��5}� mS#!@i��K8&�H��,;~��6�=>��|(�A��V��>ގ�,޵��)����p>�u�V���HdO�r����E�����5Z.��}��9���@	�5����gv���Ϋ����p慃��;[7"��"0����j5VF����1F��A0/�I�(D �A0hc�����f٧o��h�:�!#���S�C��B6�|Qu@4k�8���Б<Ue>P�K�_�	����vF�FVh�Z��{2�CdQ��6���%R����&@D��o}$�4DK��Ϻ��M2�y�</0�u�ў�c������������C�������(Z2c�� �=��峗����ǳ��`;o���� �[rC�y��b�8�y�G�9\a����	��8'�@��`�
+�8��<X�30����|��4�m9�
��u�BFfh�{��w��wv�DJ�ᝑ�>�pѲ�'�mP����5�r�E����+��`�f�p�Z�p��(l$֟�bW�qP�5�33�͹pL��7���߿.X�=�׈,�1W�
3*�z
:�F����{5 �0�e���9�h������[/�,��Wmn+�<
Uٺ#����U�PY�Fl�۴b��}ɸZ�3ny�f��5 i��ׇ�Ψke`Ќ�9�Yf�u��GC�2Y~�؟�Q���kL�ln��s�G��
Y�Zĉw4f`��i�s��E�8�g�u?��܍���1��.�w�K��n�9c�||����5��{h榒��|s�� �b7�<���k=3���q�-��=�8���itE6��D� eϜ}�s�,�W�(�+��ug�eLH���J����~���%�H�3�zM'�u�t�=ݎ�!j�sU��Qda�(Re�<(8ڽ���3�i�S<��a���`�^���KS���@<��)�D��Z�Z*^��9�e�UWs���m/�̮9�N]�쀦�����1���wl�������-��2�K�Z��N�k{����8#=�(�;��(ɭ%���JkC٪�B�@����|E�?����d�"6{;�Q5�t�	�)�bdMe�p��� �aS�٭�0��_�;k�>vgb5�3��槰�\��n̤XP�@�0SV��0U�)K�ا)x$]<�e�v1��>/g���k�C���0@����j �� ��5>���$j݄!��elv�(�ǅs�넱������"��jF��K���!m ��|�Un�:������-���@�;���A�TP0��o���_�5�j&�Ke�0gW�.�P��Bd׽
P�#������ ���8���{��v�E�N�f��H%%h��Gn�+�v��W��d�w>l�k���u_ԧM��z��|/���0�P�E�������q�(1c���;��E�^0��1F�H��@��A��o���P
�*r*�ۮ��3�z����3��8J�<��.���YG�x���1BѬ��k~���o�T�_�Q��#��Y���|��sD4H�i.��ܜ�Z$��l�1H�M%R/&��%�
aU#ikt� Y"Jh;ZI�u�57������GfQ5�&QS!hJ����G����KX�eIfmմL�O�e�gN��'~�^>��* ��K�3tjQ�"����U�:/�Ԅ. � �}Ҧ���.���m6i"�m���[,���8�&N�-tg�*��A�%3s�[3d>5���O�X̧���vR�Z[��ڝ}��3I�{~���9iJ�,�$f]�ܓ89�%�]��I�L&dN��MDA�7Ϭ9P��'I��`����⌳չ�� N*�`^n��@P�mLη����0�"����,�m�G�V�L�~�OnƃT"�̘$l�����ǀ���L�(f�AODx��L�� jew$A �a�vd�f<�;�hs����g��X��,�"���N�m�8�Y#?&rVЅ
�͘{q�I.,���ƞA���n�٨�޵���f�x?r\&��=��hD ��46M ��FgA�l���5q���*�5v|�"(P������D0<���?��;0ʴ���R?�
�(]0�2�fC\�L2WG�x��e�)Oe0*0���=}'�q����á��t���S��x�]R��XF�<���8e��/,��^WF�����7Y��q�x7?&�Ծu{�NKv��[o;7�;cmw�AFvB�N������ಥ�I���"	�2���v�M�Z��n��y������nw��;e��L����f��'���+���U2u'1����eq�ސA�e�f���"W��>N��u����Uy�~'�s2�$z@��42�d;�w��������n�>|��؁�������$�n���}-��$�>3�,�,��e�c��֍�n_;��3I�@v��ŵ���#�O@T�J�j�͡��	te5�-A�+d������_md������A=c#΋����S )��	ۧ�W��Io%a������W-G���֤���A=��#��+K��C8Sm����&ݓ�`v�)���3��~y��Ͼ�.�'&�}=c`P �v�#�'o���I��Y�2�
jxe����d����K�',�˖��s\�t��v���޿ъ1�L����l�=���Թ�)e-�+3����1�U�������d�[æ�ޑ+���N����g8\D���'34�����'�l����[q�*j,�K��u��ʨ�sꁙR��
c<O�Z����~�,1��j��ΈFc��5�NV�������W���7���sS��9f,l0I��
�0�,��>�&-r�������y%1���E���FXh�Ct�˽.V��X���I�-�/�c�?/�a8��R,.�`ny��{�,M������q����ay�I�dG��M��F-�ԋ���'�WPu������Ho��gh��t���H���65QhN�Y�C�tQ�]�j���\L��ZX���9r�nt]U%��cp�*1#I��\n�8D�2�\`b˜�L�2Nf�Q-��rE�Mr�~��g@i�}� ���S�ʪ�=�)Y:�C�<�X9#����8�ƨ����{L�e�/3Ƥ���������ds]�� ��/bq���y~S*��>����zG�c����!x�d����ɀ����9���1��TUa���F������MkR1�.p�����;�]:>ɚ?h*����qA��>���nKT��-R:|�:�d�?�i&Q��.=�#�.�'9Q�9��I�@{P�!��b���6�2=�}�e��E����,S���Z�1�Ԝ)����M�"+f
�\�A/%�\�*��<Tp[YE)ڐ;�������2NB� ݂v��
�,BdT���!*2�A��1��)��cKX+s�����4���I�<�f0U�y���U BF�C��$S�&N�sک���}�I�]���?sf$����Y�(�%[����㺌Bd)�c@��F�Z��D\w^�k7m���aV!v5)��󙯨����?�Cx��	���,e IUàp�)���EW�����O$�k@F�9h�A�O_���i+��\���S`b�8��p�_$I�(LQ���@_q'aa��D�рܵH�ԩ�|���YA��������"0�������z�@�j���i�*c��f��\��q�y��J�KBF�X'������M��LYAU�H>���zU�I�M6j����R�����aj
�^�"��7c�I�x��jB�$ޓ�30HhJ (���w5S��������\��7T��⅙��KU�suB��5�e�A�$��,DuI�B��U}ͼ����'���FMͼ��c�2����X�Yw/7�Y^��Y&À��]&�e��N�!�j�$��end͛,�����	rs�_�80��EU�I�̦ٸ�mV�1�	�����i�����O��-Z؎<a�X�ZE��)�2k;) ���$����򪓖��q�����$�;�$���
�(Z��rs�&-������z��N�`��I�E�٘+��{8(�i�l"����Dn4{�2�;*�$#v̄��Tm����H������ �����O���%C��Fዲ��L��;J.{I�m|��BL���D`PkS�;�� �!�?�B����q��|M�G5�$EY�jqY㫵�3��m��-�rI%_�s3�>�T��b"���U�bT�m�F��:�����e�v�
�C\�Qc�=G,�"
�����M���G�TZ��#�q3z�HpWrj�l�%��[�����Sg/bc4E������1)	�S9E�8���[�š�=���h�)<���揟ŉ�[(�>���)� A���|
$���&��@9� 1�eȢi��J����i��2@wѦ=�M�,�g�~P\yW�id8(u(�P[�a��Xň�.�F&@-��e�ʂ�H�	�����Z����� �Bp��Ě��a�HGjX�z]Q:c�-����}��Z��������k��5�P -�y�#�l��G2�b�by�q�#3833.�g_#~�p��i�-82c꫕��<c	���45�Xi	h��f���	�Y��WbH7��c��&�@�m��*Q�If̴�k�]�HP�&qi�
e3�s�,���.;���A�����9�6���@)z#MU ���GY���d2n1�ʘ󇖡�5�sv57��n׬���{#�V�G�9Jc�u��)d�8OaӠ��	�E�1�ߚ�� ��T)�(5��l�m+�B ��r�����[��d4���Xlk���#:(-/f��5,H$?t�ED�͟$rN����S�CY�@ܫ5�� ��!F�'Q��{+�I���͸�ѳ����S��3��k�"���A�S�&��%Y֙5��Q��H\��$����C��/I�%1:�l@V(�bD5�a�,���T��"UM�j�M��A%�`M��Tr�&�"�����-�T65�4ӓ��O'�X��#L:�f�a�Z=��v�d���J=B �	c����e�ǜ� y�+�uR:�d�í����@�e��fIE�z�Y��IUcs2FAO�aƎє�^��(�zИU�5��U?���W#YG��?6���Ll��J��c,���KT����昌��YR@�$�R������2��B(�k@�X�W�rA^�5�vL&Cl'����&y�ngE^(ê=(pod�����>��ÔkV�V��v����d�A�#9�|?E��ĉ�OA�.�0�N����,`��`C�6JP�gQ�3�6_Wi@J\>A#�I�4��l:���t��Y3>#�t�e�\h�p�$ �i��m9E1)�!I�L['�`2�%Ϟ%��>��ye�E�kD$���J���Y�O�5��M�����D�*��H2"�L̬���%��\>��0}��%({���0�w��Ȓ�t���u�.�릈Bʬsۇ/6l��)�nW$�dRPg�߹    IDAT�����������de�E�L�2Z�q��}$�u���8�V$V�(+Ј�!)��L�ѡֽ.PLG��JDp
�	0K�s�e�N�����tjrXI�mM1Q@�ᚆ^��J�U'MP��S��)7�]ٯ�k�)}C�iaĪ�]7�U�#)�k�f0���,D<�d �s�8QV��?eKI҅R��;c�@��0�4��Η�ҘQc�2������$�L����*.q%N���%��y��5�����YXܧ�y#/����J�F�q	�y�_�"�������~����3I�5-R�о��D���S�:�]>��+U	$�U�n�Nx��۽gv�~[1n���$dgH�^$AJ̤��AkM{�0p��=];Ÿjg֜>��1cEK���A�Lѩ����^ܴ���+,f���,ߔ{�L^��	P4!.m�̋����(��}Qǩa(�WSa!�p��U�z`	KI��Jն�.n㯾�x�������a�2MV�,6�#]��hi��#Vp��U�[�G�:mW#�>ip��<s�U�N���%����h�i�Me��)~M�%#�B�C�c뙕�!�G0�����ԀZѦ��U�
�}a��zك5�4L�2`��%+͍�(JTt�Ijr*�����Y&��Y��3���OQ�NH�\x.R�dmcF��d�sw�I�j�`PG�F�M�K���=��sY��߀��C	5�p51; �eQ|� i�oZ�@f��u�d��P�K�%��y�������Xy���i� [f�#7D��ES��k�V�?�ɞ�+[C��+*v���N�Z`�dָ�k�ƀ�&��M�`,e�Nb���&���@4@o����n�����:S����d����u���'o��=��:�EQ��f��P�|{[:�N�"g#f�C�cՎu�_�2졉3eb(1�εH b5O>��}+��9>t�W�/#Mc,/.��VS��� %3���T`�=� ��3td��5)t�3���������J1�<q��):iY��d4(d DCe]�H:�%�3y�:�KӽhOY���M�S1�� ��./
t2ʖm��k��6��x �&G����f���M���	�2�t2��H:�J�f	̮�!��{P6!F�J�c���ZǪ5 K�f0��T��H��������fӄ��=�[�a�!Z�5�����s�*@lj��Q��.JL�2���� �& �� � ps�2&�hJ�P&�I-����U�8룿���CG�]T��3b&C5���@S��S�,`��|�Ţ(��QӲ�F/
)���K��6I��Y>AU('�(&��[���x!�]�˚%�q��=�""H85b�wT��X7���(��a�:<我c<���d��g�X^9�����M�}�d�$�\p�ג���H��$u.+��W������k�g�N��q�����$����N�$��]��/�ߢYoQ�G��QG	�y%��@R
2�5����G��vj�|&C*����*��@N�Л�4�ޤ�4uR�j:Vc�|�
�|�~��FL'9:�.ƣ����9�ң�l�(�
�k�O���_��)�G�WV3$U��m"�4���!����-`�Ү�m\��k����Q&Ԕ=��X�d��P�:T�Uۜ.�/Hݵ�~	m1a�F5��F�XYك4��P�$=qYoN�RS[c6�v��#S9�L��5�#�ڊ�˭7*BH\3���S&N�U�Z��2���ʒx!�|�N"�R%G>�@ܔ�X+�6��"�g�&%�� ����S|Xp-$��R��$���JFԌ��dmmU�����"�dEӢ��68&��*�\�e�,�����X�o���Le��i��������PJ�T|��(�(�c������;yߴ'$���+(�X �$A�9�ɴR$59$u���&E�1�G�B0E�o���\ �7˘��y!�R�u)�ZO��gL�"�H|�W����L1߸h���Л�#���P|L�zQ����,M
�(@%%^e]��q����}�O��l	�-�h�,�ȮG�7�>r�kW^�?%3
eU�GBVe�j��`Y$���	�U㟱�&�Y�+��5�>�������2�V��f����|�G�|��w1�tY�A@Ǯ��=tk�e�
Ah�6Np~c��ً8v��Ճ󘪜�FH��=�s�A^�#8�]����s��~�<�#�[°�/BOB���9ԗN���o������pd���.zdP��L61����?9~�?�#�x�<��%�i_�a�����1�w����I�#�hܼ�NG�����X#Hcf�AA��>�ԶI�#!Y���e�EU �µ�d;�3'k�F(d��M1�L4	�n��D@�o�7�5���v�ê�e��΢sG9E�O�R���2�j<!@`JKDI�.���N���]Q�6�k�j�Zx�W��,ZK���ލ߰B�CAsS�(�CI���,�):]cӨaF�,�R�iG�i���V�Rp�4�(���Ν����5�d�B��n��QլU����-�5�qWQ�ƈle��Ac�Kb#G>�F�ʞ5�D�,��2p�(��0@�-��I����l��o�ο_uz$��`�|ګ^@���i[�L���7��M�e�~��d<UPJ#6�e1z��I������G{�Y���5��չn7�6P<���(���hIaeu/6�'h�2KG٨�%1b���R@��=���͇V9�����H�1�Y'z^fH�8���E����g�
����\�����2�5�I$��r8�.�5�{�phU�C��1������`6bWc�e�4�6���2Hk�nf ���)��%�z���#J,_�G���H��mTέmakZ���A6��ز0b�Yc'�ژX9���o5�6�)6�\�\��}�K�Gc�>u
����[X���E"��g�1I���ٴ��M� _<��n_���j��9M�I{[c����y\� �L�pe����>�[��&��>���^z�*DؙGuP����5Sk��s'�qMƴ?�]��d֑A�u���Y�|�(ꑲ��Q���T�� !� {[�p��2�]Ğ��0��k�)A���������X�"��eY�l��B��y����&��I�C�������3Ǟ����ބ8YB^�n�NF �sR߸�_��b�R�L1D?S[3��{W��<��{�we��6&���9�$�y��i�O�
D=�iM�l�k �f�W�l�U[�F�j�WW����M���)�����HEO���*h�E$P�l^���>y׽�~���֦��A�`8�`��<�~��I<�싺��-U�)KE��#W�F,F��B��m]A���`i~Ǟ;�g�9�=�����u 2�!�q߲�F�{�����+JfR����������iK١pk�zI���zn;��NԢn#nbiiQ>u8a���+�����'�D4aA2�6$�kb9���#�[㻯-Y�A��8�4���1A�-���
Ty��3Q+�ލ+�~��[�c.����G�)uD.L�H��_~k[z��n��VC#��{y'�&�@ھ���b��Kq��b���8��8y���K+���7�!�2����������@�Pեn�^m]����D�p����m��������enl
huY���"�#Q��7�1�� 耐���#�ОiA�5�,3q�^��b�H�~���j�����>�k�xA_c1��r�z{{z	)�O)�ml^�`a^1��p�iCit�)�w����Lvo�w��H6����j9?�gM���7�\g8aB"!M�t드�������
+�1��}5ݘ�r8Wi�,e��!�Z��Z��37�D}~L��2���٤�C�Q��V�j�3��羡Z�*�4���,$�<��r�]܊���b��LAa�;AE5N^��c����kۨ{sh�L��X#.K̷5nݷ��ً���Ϸ��������*���ɚ_�C'�p���hGW������o�[�ހ}+KH�-Lj��7	1�+i�+��{�8���Oq��kh���̛�ѥ4M{�B����^_m�eM+�3I36[PF�OQ�Eg6(B��"�t1�i "1�{J��DF�|�۞i{Ս��1&�T�͸qk�m5��u{�����:���Gjkd)�%D�N#�����F(ɋ��Ϭ9R��8@9InÄZ5�`:ޒa`g��;u�YH�b ���I����'�SF�@(3R���`��mw�
���C��v=+����+3�K�>��Y�|:cCKF�Ǎ?�y�W"���{�S�N�8��&@��e9�dﻝTO=�^G�X�i<���7XP�QH��%s���w7�y3�R2�%3�l��%�:��?�:)ºD1I���u1�Lqvm���lI��� ��Mb�	���b�gM2y�+p�j�X��#L���� [��ʠ��3Ȃ��%Ƒ��I�E����O���IEl(�7|+�غl��9�㸻n�.~����A�~��:!�������ay�>�i�&D�#lت:���)2ʫ��*��:��?cK��	���S�^���B��sI��o��(�[�c;�$x��������6^>uO��iK�/vl��U��?r��;M�d���J 5f����CY���*��_7.���S昛
���Q���0^��[�/�ӟz�]�xl 'c3���d+���<�/=��sd{�~��81�a]��~�>�7����ա,�څs����{ޅ�<vPw��7x�����_Y�0�0�VH;}��`�ߞ��Ar֊V����r��ţͦ\�����M"7/#nj���w�#x,v1����߈��6�?����'�!�[:��asf�R��xT�(���732�hR�H����W'P�m�VR�og��Pg�9q��ײ:*����(ЖCt�|�Cx��7b�\�4d/�V�0����|�+�����[XF���z08���Y3Ʊ�K�D�W�lm�����W>�.�_����|��{��6�꾛P5	&U�ub٤j&�rM3�nA�/J�r&
x��P+��/|�8zd�$D_26�4�bZ���[nڏ˓����F��}\�)vG0C�{������2���r���[apC),}I!�A�!��ɝ��J���D��-0�!߼�<|/~����sz��)(�j�9ia�o<q_}�	��,,�Q�l2-L��n�.3$noG"*ygȵ>�x{Go8�_��C8����_8����7q��y�ϯ`0��iEIv��k,LM�s�(sg&�1�Nݤ�F�0x�.�q#I����[L�6q�u�܍{�ΡG��dv4�N��U4��3�����q��t��2����qb&eV���]f2R���L�@'IQ�X�.�],IP��k�'�I1�g��3Ui� �7���z'�z�
z���1�j{VE&�>���s_������ ����X�˽�sC�đ~l2�i�oy�w#��_8�3�wϝ����x��x��O�ճ�%m��������*%Qw��8)���d#�v����ͪ�9.�cL�[���A<��{p��9G%Ґ�ۂ�V4��?����ޏ�AS��� t�G�^�2�p��%���1��9�1�LT$��/��Wm2K,����)3�,��xF�c�r�{n:�;oڏ��H|��i�^��o��i�i��k�8��il��4�I�3���UT����#3�$�k��Ǆ`�,�qd�
�u�����[ǉ3�a����������<��H�7��ן���|�h���D�N�6��;�}���>X��xErV3Z��m����m��)�8S=5�B,��r[�k)	/'��	����>��&ܵo����lt+{�*��Y��s�=l���D��'.���O��!��?@N J�WۢS�n��o���}������G���Pu�8��b��kx�Λ��w�w܋�5�t��&��94�T1�)Ɠ9ǡ�bcR�ϼ�?�ܗ�/��[�fu+��E>V���n�yb��A��:�鄇_4J?KJ)͡u�JY?R4H�sb��&���C4QC��V3�b�3����4Ġ��D��ֆ��dn��%���HF$M���4��͂y���tD�M�&9@SNPO�8�on�� &[��^_���e�,kk%���s�2.��+�T�E9/�J��2���YS�m���|N�j�������jc��Qb�c\w`�=�ՅK�X�fny��QQ�I����ҩs�!LzVC�Z�fJ�k1���%\�#BȌT�m,R<���ʼ<�������0Xڃ���:ds$���As�����g%�o�)��sJ��#Y�����\|���o�/c0O�*�q�w3�2lll��N�O��\�31����ޡ� ���)3[Z�?��d�W������B;F]n�_����|쑇qpe��!T	v9h}�]��x
_��OФs���`1����9T�	���]M8�^;���W����ǝ����=�/?�_���X�wM�C^d��� F`���� �B�ް��,밤�2q�Obu�ŧ��c���:A+�kkT�]��T.������O�9\��љ[Q��k��5��g��l+R��13;i���|��:�\�ٿÈu��2N�eŌb��9��N��o>���?�����=bu�Z�+r�t{��Ͼ�/}����5�ܞ����_��fj��u���ˬ.�ɱ�~Y{����?tV�p����s_����+�����i�I	L&$��,k_��YYWŚ�G��ڥs��c��]w6�����?�� �{��=r�[�a<���K}�܏�(�ƨ�_|�kx�[?D�pAweˠ��&�ufVr��16�O�q�"�KNr�'c�Ĭ3
�]I�*H�.��]7I�
���F��&�I����>�n�'���Y�1C@��(�t������+�E��Y7�;�QA��9~�*�)���T	Дc �D?*���	<p�5q��O��/>�w�xe��GnƘ�tMY�N��ݵw?��v�+��ӡ�Ǐ��0N��8����}�8�w	5��k��ވ��G�������6F5��I5k�Y4I�D�n�/ST#0�������Ⱥ�doiw��T���9���2��g��}���{���O����uz�{l�FE�3g�p���={Y�Hi�y��t�Z=�|�������̇���طo�<t7��d�'�]���u���+�9,,BP�i��N#wΜ�Vݏ{?��Z�$��u!60HP��O
T�7\�}w\��1�;�R7Q�ᚒ�^�����<��9����Y5�/�Ŵ�����'���j"�kשR�www��4<\/�EK=(����7_�kWI����h�)F	�V!~���n\�Zacm�cJ�kTTE����/}�;����}��?7���H�*+�M_LNN M���9r`��y#��������r��:IHO_����%{�e��e�L�LU��z8ex\��]G4ŵ?iк�sQXf�5��6�l�d���݃���A �<�81l1�1@�����ʰ�6�G�e�;u�-u���\��?O�G��#"YMm�j�w��oiakK�H��)�&�I�ޖ�!��w�mx�7��"%�tY��cH�2��zpc\����ϟĨ�U&"�����.�%gQQ�N�Cz���-��o��F<��!���va�?��?}9���ͩ��(�;t`�U�������C{�/t�U6Tc�����M��p�m�e�@ f��}B>�>p<���M<��i���(fc�Dt>;������2y6!��'���Cx��qC/�<oNieg�[#*�����C���⹺E�����y	�ׇ{��|(
�sh�����;nD����_�/�]G�t u�������y	���,��z��G߇ۯۋ�4䱶�\�gWݲ�WkK=sO��ir�i7�k���_�~xb��2�Nߎ	p���NU��X�� 1@ο`��z��xn9�G���,��<�#E���̚O<�\ښjS���    IDATP�@���Gm���0D�C,ٹ(�c��D��[o<���	��-|����6��=HҎC�o	����I�3�u�t��٢�V���h�$��z �{�[T䙏�X]�c>������Z�8ui����7q���lUd�uk+n2Q{:��Ѓ�kq�W�����n��[ ��0ݾ��������G��\�o���(1t�9_6M݊�1�տ���ď�W1��c4)�0�w��80X���a�D���0Z������o�Ƈqp������ߕt�������Fdo�XYៗ�����*��q�G��{���st#�φ��
I���>~������/,[$W�F���k�@w"��]����wE�`$�t�,c����p�~�S��/𝈚�W61U�Rf@����ŵ1���s��K����'�մ�Sa RDY!wdg�q"�<���>����w��R?=�">�ů���[܇(�����ց��Q�k���৑�JU`M[L�([I�Gp��w��{����-\xYr�|�-����q��=8�^����?�ٵ-A�`���f=׌�������u;�/6�dx_l���Еd�N���nº+6��S��J'���Tf/�9���y�Ϳ��������ҋ'����W��0.J��M��\Q}S�e:?���MWH���xV��Z��$��na����wޏ<x+����g���_��}�8�8���C��ol���1�%��WD�YY�=w߅��k���SGH6��r���r�G��d���9�,/`�qE*�n���f<��{���������a����JjiM�h�x�F)�#ILK+1�KI��A�/s;�����Ʈ���j�)�}=�V����l��kx	��o��/������-|�����^:��W&N��4:�8�m,,�|�.�F2{� N��\��j��}m�{S���^�͇W�ȃ��=�݀ ���/_���ckڠ�zaw�����&%�;����1��dV��
6�I$��n�l���P�0�4����e#���5��	>����nƅ+c�o���=z��Q�&@;�'U��G��Mگ��zMh�k@�^��u�]�n���.���e)v(}��#��D����ת9C5���ie?��wI����Wx�'?A��I��*�qb:e����ED�+*6�c`L`�d��E�$9OFp���O+4#���c����ᡷ߉�N��^:�/|��x��3�[>���>�q-���b�B>�����H������}�8JDB)�h�<�xsq�=�a�c}�2��ߏ�|���}x��6~�3�1�����&�2�g���$+4U����ʄ9Պlc�hݫV�㒲��q$�,�τ�T'�lS���n��K~�Sƍ�V�ұ���|�d���b�QUԗL����5���YD��Z3uͶ�O�������tP�S,�Se�����|�ux�w୷�����W����>~z����}M���PF+0���|)��j6�prǯ(��u�D)���1�>����L��^�wc,2��-Gq��2�]�}��dǁ��N��$�b�'c�<��/w�K}o�kr͒�[	�����nT՘�Q��8x���d��{>��X�f8y�>�<��
�8�� 6F.o��>.P�<D�ѳ�®7��q�n�T�1+���H�6�!:u��V񮻮�у{D��|�2~��q�Y�����1)3�:������h#��L��J*���"��4d���2�|`	��Ht��Q�5\YRό�k����Q��`��,w�8k!#ׁ�k�[L�
�-�x�޷�W1��n�u���vN&���N��,�"��em`�zF�� �N^��/�A�� ��1�v��X�Z��Λ�����m�-b�� �|��S��i���+����G���5�i%+�Nݱ�D�v�t6a��4���?�\i���Hc?����o98@F�6u4ar���f|�}w���d���E�����f��3��x��Y�	{&"z:2���*� )Dd��|��b�����ɇ1����'���ë����ωIf���S��SNd�&o��K���-⧣�v�>��3E���n�G�u?|��N����ؿ4/�ܟ�c�8�+�����'�=����H,����_��l˂^�úK]���ϒ�|v�5��f��y$�y�a�҇߁�4��s�u墤,����+��x�'/�_A0[��f
t��ՃA��g�m��l���I]`t�<�{!>���x�;n����{�>���ǳ�ϨV5b����2ҁ�;7nH�ӓ��y4S�NpV�������Ƙ�����ы�Cf�e�2���>��q�[���M����8�]�?��+2h��X��D3�kl�X#������Qݿg�L�hO'ԑ�J�i4��/�ӿ���܏������*�_\ǔG`t��[��mj�Qg��5b��e�ծs,��.��[����8[/�p{z){���Cw`a���������Wq��Sr��8��q�Mצ�6��ba��ؾ����^XC'�-u�n IP�c�t��k�$�=��$����~�W>���}�4�_��qik���=()���f�!ٚ������h;GGӸN�t��~_ '
إ�d�~��Ȱ�Z�I�D�[�J�d�7.�=w݁O��'�gy�ןǷ�������~�@\�O)g��Y��Zk� ��X�ǔ`P������F��w[ (����>���p����о>^:s����w��	�v�_XAv��5F�pZ�cfq&ӑ�b��}�ܾ"pl2y6�4%����Q��s�Pc����?:?�=���5�:!>���W>���,�o��_�~�OQ�<wA�
	�a�^%c���(�ţ��틘$;��&������M<�Kd���6���F0<����{���&Ȣ��s(���/��/��wނ�N��g>�G�ǈ�%it��L�N�xqeE�I��E�y)��f�ي쩮,�����ވ��&n�n>���p�m�
־�����.�2��}�
֨��q&ɧ��3��JjoZN1�'b����P퓗�n0 ik,�u��y	M=�o��?���;��k���Ǹ�>Aw� �{lR�c���� ��L�� ��ݡ�G��!�f6�����Kˋ8��i�<u��(��&�r�q�)�T�D���������z/z�~��� ������(�F���`�{���V�&�.�����>���9��; ����#�z	�Y������Y�c�{��.5�y��Ʒ�ӗ1n;(��+J;�D�t,��U,�i�n��e��гL�Q�T�l��X`\�TX�t��o��O�-���S����Ҵ3�ge<�]y��ڹ���A���Megfv"�c)c@�
�UTXц�ΘR��5���AqX��^��G�����qh�
��ޏ�g��(�	Ke�$�E��y������+�����ŕEDY��$��e��P]�s5Ya�ք�����,�!9�4H���܇;�r�� �2���Oq�œ�7Yo���3`\'Y��f�D��;�{;�֩�$�dY��=#h�)=�r��yKJ1�)�1>�����ť����?��1;R-�
{����J��Ѵ��u�F��?*�l���:H!�t0��fT%Fe�		Z�Y��!m�}�ށ��.$i�o���ޓ���Q�NoI��&̨��w^j�)����o�cb|'��]��^��K����	�Y1A�-pӾ=���F��̥;�*^~��oM1��QET��8�仒S�B՝�m5|ڱ/��$
�u�o#"y����|�+�UN�j*x��>��q��y�m7��7�S[�4C�n�jb�J����:Ɔ�*kJ̵>���pǁt�Z��ߌ3���Yj��d)�
����a��4��|���y�J��z�2j��m������'���iÅ������n�b{����x��;�o~��8��,��3��2�q��5 D*'�̏-�I�Sc#�I���s���?�9��^�;���;;����j�g��eJX�hGGL���'����c����c{��ؑ�w�
0,*��G����eYW�"uk��c}ץL ��p�!��бD5����>��;�нo���N��m�x�,,��3XPZ���L����Q!�X.�:�����*��}&�E�r;������<ҐuxSl�]���y1�w�y��������Oa���j�@�d ��UQ�=��U;�N��9�u����+̐x�oV��S�9)�$��d�2��&>��Ⓩ�]������_8fݣ�T���Z�&���@YҊө�Q�jpl��}�2��D�ɰf���x[�ypu���<����w� Ͼx������g^@6X���1�XP��v��CD=�7;i5����3���H�G�v��(��t1�V�9�{P�?Z��4l�/�⃏�/�����3��������'�U�f�$ۖ�������]�جN�ζ2-�"����7����Ui�,g	���u�4��?���ߏW_��o����̹�:s��-S��$�<f�>�rd�����;�/�p�Y��X����p)�۸�*�ۿ�}��b\���̉��'��
��:��~Q�F����]h�̅r_�-��
�)?�l(�d������՝D���A�dζ7�P��K5&mn�.�ӟ�4����4ſ�����X2K�{��ɯh�E 9�;�m1Pg�J�-:r���ػg�}���35�K:T�S�y�d�����B�%���t�����f]�|�\\�P=��P���r�x�j#b�L8�[�:�GG^KVg{�d�V_�9���Y>��|7a�u�[ݳ�[n��݋*�p�Sx��il��(�,U�q@�ް�塜���m�i�L�;*�U6�!hs
����G��y� / ��FX̡�v�<n�
��(�q����{�%�����L6�`'=f��e����6y�����q���xeg�^T��t�J��~&���-������|�ͨ��s���,@�o�]�o��_»��O�������� ��E�Ң�8�*��޶�>����h7y�#�5�l�e�*l�3p�V<���1����f��'�[nYUF��O����ᗱ6�1O2��N]��nHܞ��8��&V�`��B���$CD��gI��D5լ�gß�&븹�'�H�Ư
ﾏY���{�W�oan���Vy���ӥ��`Н9�J9�Y��k��=�D�b�����[n���^\8w��<��x(�>�W��J����El�B"�� ���'}i������6��t y�aڤX']l�h�Q��#%�~��(G��������7�1
�-��Ո--�Qv\Op��}��@���/����>�\�d���@t�'�x��{�g��X�h~Z��BI�n�kY\�nV���܃f��M�qHh��b5�*&ه�{�+K����կ}]��
��;�џ'�)A�V�x�
O`L`�5J��3������^>)R7�0��lTq���E�J��lM�_y�
�d���[o:�_�������p�������feĲ��@Fڵ���ue��.��*�-�gH;l\G��D6���:�G@�M���v���#{���=����6��x�|����3?;��3'0H�G$�`�$�׋u,7I����޻�Dj�WR6	qg*�
�^O)�D�&m�_��O��w���6�{�g���4� ��G7X�.;҂�9�&�4lhx%������������� k+I�IN�	&�W(�����x��w>�������o�����ɚ�=����f5��qS�"}f�0�y�1�ċ�$��5E�H�=�=˸�ַ��Po��Թm<���x��l]Qwv��Ų�zd�J�ԫ�2p��T�:�R����8'�<�!|��eLV*�s�u����w��j�.�����ùQ���N���J^XcH0������7��'M�G��/�Y7�D�Ŋ�<aA���s�2�'vT��5ns5�Yx����!�,.b�c�؍w2��,����G���k1�m���a���<���/����l��&E��1��y�����Y �vDhى��ga� �¤����/�"겭tj���?Sc�}5��m��b{���E���݇�������;�/���{:M�A��H�0H@�$@1 L"EҔ,��I��ϭe��\�.o�kmY^�,��(["%1��  �f�3f0�:9m����v��Lw������9�y�}wߠV7�����cg5)���.���l�<��M�l��B�����IM��d�U�0V׹�e�[���w���.W�RуO�w~|�έ�Ti.�ܘu1fD�Pjc��&�C�y|�޳3�Y�h��g�2/��\���ژ�ü&����&}��[U���������o��c�)���n��0y�G�.DM�V
O�-�CGN�f��N�x�����w�<ų���U�&9�辊��6�O�s���>��5�����ͷ�R}z��㒧��������Dd�vJϮ��@�Z*�W��l^����&�u}�w鎛/��\M�_xS?�уz��#*U�4�.j���W��5��n�3fH��SS�&pF�(z������c�2���Mz谻�Q{M��w���?p�=T����V;c��R�E$ �v0*)h���b����48���J�"�~�oh�k�d�ٙ#�f8�������y_��X�J]S��6WN�Q�7>�)}쎫u�tK����N�_�0���J�a����t�q�z�M�3��U�����1�N���Qr#�M�<�Y>{B;w��S���n��J�u���Y��~�_yC�i�(.s��*M�ޘ�Y���n�(��la��5M��p��|nNM�e�����5��om�+_��5j���_��_腗^���N���Q<��hE�l�)��r�S�f�!̵ZR�8��鳺��+t���ޅ��9@��$[	D�)oּK i��YW�r��~Gk˞����jj�i�jh���+0����,�p(ò��W�`�d7b�K�R�LPװB�.���M:&X������E?�86�hf�{�bJ�|۴��Η+[̣5�D�#���k�)��qP1�l�?R��'�m��J�ٲJ՚Ml8S
E���H4�� ��e���"�^����K��G���MU���@�����N����S�`�e

�D��:GC��H��l��O�릃�t�؊�����:r��D���[} 	�s�u L�T��o��A#P4��E�Sd�bk�egS�Ϊ��l������۫�D�?��_���{�TƁ�d�1A���LNq.�J2��漕��*�J1g�u:m7ed�A�u^Y>�z�����gt�]����X������z��fv[��9]� � GCȲ��5��uE}1���R���z���|i��/?`��W_��ߵW^�=�3Z;V�	 LDd��!~�}{�usEc�0�M�i��ٳ�����&�t�@ˎ�	�T袽��z�ͦ.8�Pega�RФV<��Ud���$��]�V'��njfz��U����ZG=���|W8�5H��Ӡ���$�J@O�x<�Ȋj�0��H��ܷ���zݾ�5���=�5*��� ��ǻFVfl�E:G$E��*2CW����KG��֙����[��?׬�7_��ZI�Mj���ءi(��+���k��]jNխ����՛ E���B�z�|��bb�$`�h6�hh�'�p�Y>,�ij�{Dx�y�P�����ڿ�.��J�ݿG�\U��M��}Q+km�D����H�_b�0��S6�yR�`�I�5Θ �S���V��U)�\fn��O����%��������卶r��ƅ���|Fޑ-F�1H��\��ɢ�l���%�ԅ��,<�d��c;����4��IFK�IG���J��n��J}�Cw�93���{M��{I�ϭ�x�R#N�lO��dF�M2�b=��Կ�sa��<�K5�/������r��j��v�-�����0eo�7����N�L��b0/}�OB���l��d���(|0��AC�h�!��3    IDAT�.�i��3&�P����X�3u�۹M�RQ.l�ȩ5m���3HK�B���1����.�MMB:�c�f*y�F�H���HS�̽6۷��jnz���&߸GE�+h�_ҏ~vH+É
ͦz��O�nKs�n�������x���f
S�"uWO��s�����i}���tv��}C/kh��A�/9�B%��rr19��O������ʩU�\��pIg%Qp}�S�}$�v	�fc譜�=7�O�q��Zk���_����8�"� ��D�*�T�Q,,S�/��C8r��(�����@\�ǝ.�t�y�.޽C��{��~�E�zz�W/�'��Ro�<�Js��Md{8r-�Ymﲨ���˚A_OP�|����_��Q㦿�82��N���W�x���~����g^W}q�&��� >���h�F^�C��M�o�P�$E���"Ԇ3#��ӈCƘ�nO7�fp [j���g?�q}�[���������	#w�3(��3M,�v�UvР&��]T&��hx��6푆#��؅
�z���_����s��8x���6������_��=���/����r�WL�­.����S�s���Sa}&���;Sݠ6DX+a�vx���w��%�v������������;��r7�,�)���l�vuY�aK���6�Ц�/�R�^z����z��c'�O���i�hx�l�^���»�N��!�I�2p^uL��x�N�݅M6��l����#�R�Gc�n��Fe.d��d�K���C�5��]���7Ӎ��场�5o����ڷ�"��/i�����	�v#pvQ
���̂�94i��=Oh1\���=��F�0g;v�L�^�h��,k�LS���4U��0B��n���ښ>p�-ڳg�VV6t��t����p|O�q�A�;=���#x��Ţίut��Yu(�w�p���[oӯ�q��4��M�[4‧)-��Z/R�06�aQP)��y���n�A�5j�G�� �����d��qԈ�A��§�b�������'���������8�uF��Y-��F��(��#&����m��,�	����:�DC��\#�7P$�P��\�Hl�4Ѥ�S)�=)0% �g�;�H`7�6^'g9&�1{gU!���'�`Or��c=��z��'����h�3P���Żw������4�Ex���;|KR���U2�f�[C]w�ڵ}^�^_�>���,o��C��{�1Iأir��Nd�rk�)�+�9c�3´)j�j֛fM0�m���t��[^����X�FE������'���NZK7�4-�2��j���;3�鑽�gs"���+��RI�jM�V���[��L�QI�?���+>7%(�Д�t; P����f�YbPo,iy����k��T�k��]n��?ip��ѝ7_�"O��
�Gts��A�8Ss@��v�͌��5-6�ذ���d�̎s4u<	 :a�z��Q0Z#�Y�&�LXb��h@�>Ea� /�N8��f��D+Kx�G!Ip�`���4)p`x4�X��-;�:���GN� 2�^�����Y�N��b*�55�y�\��G)���#.�G�&?����1=��۪�/���U�t�Go�5��Az��AC4$}"[�L; � @�Fq�:�v�bb���f;DX9S{��M]wDm�����gX�B�a���SґT��{0�k8j�X.�93�R���h��V���FH�kg���ZJc��4 O7~D{���﷧�A�6H��%��?�Ŝ��V5�l��+/׾=۴�1��yL+�6c�u�L-��ME��Y�nQ?y��2_CM�	�)�����]XV��vN�xL��Hs��T��}��L��4���Q���κ���v��i��=�֞[���چ:�\0tCNF��ߩ́ջ��m�?�%�c���ȍNn�^�?� _h��`�2�N����j��� ���l��u���̫ݦ16�M�O���B�d`@��#�M���4�`58�����:���I�8O��j����d0@�C�>b4v؈˙��FZ҄k�H0\���^/;�(��b`-g�s�����!�ċ�(2�Iy�-]��rw��?�fvh8	��F-���	�;���o}Q��x��q���T#�鹿C�M���MJ̔�@��8ו����z��YMJ!�5���<1��n,	��ni��#�p��e}��7?s��{e��?��^y�'snvrŘ�P�f:�4�ϐ�����	�}�N���"��6/�Y-ic���.{�>���?�[nz�)��?�����8ˤ�O�?�t���q���R� �4��u�H��tvQ��w��M$�vsY��:}������?��Ͼ���.�0󢍈Ġ1慨� d��cN���lj8�	F��¸�ː��Ҡ�L�y�K}O�{6� ���*N��O߫�~�zmn��_���z��զ�5��Y�[��9�F���{F=�F��Rz��l��9�Q7}��I��vN�����潺���t�k<���;zꙗTl�)��g�F�ç�ie��02c�:�p�f�I�,ΣN
̤�`,O�<� `�d�����.�7��Վ^z�z���X��M�BC*7��*��/�詣j���^��7�1]��}J�_s�5U�!�h s��j��yL���������u���fHc��R(3��3�hƫ�Yp��I���dN�Qń��;����3-�x��,����K���ݵ���T��
�PT�9�N?e!�IS��X�[�K����	5��:�}��k�>RX�+7v,�}���s2�HaG�:��^L�;P����9:#������&�@���۲��Kgt�����ߦΟ=��jM�q�gu���16�R�<$���?�䚵9�=��� A*�:�҆����<��,R����f-8�a�r�w$���L�M��,���χd��%���v�`S]��Ћ����M2$�f<a�s��vw���t� )�mv��MG˦��I�9.��քI��n�n�9�Є��n�9)��@#_P�ԺN
����p���xM=�+�S�ޟ�Y����꾻���ن��#U��w��Vykn�0�*��s�,׀�|��ZU�r N�ayc��N���V�W�vGC�>�e6���#f �A�����9�z��SS7�JEƜ����f;��ّLyUj쿙n�]��V:�/ҵ�D�sD�H�71�K���E&����t�4ݜ҅�uOݺ��� ���g���F����5�����k�������~�VZm՚5~�ڴi���Ni�bC_��v�[�Uw�ci	�,�(���jJ��l"��b5�*�qL�r�S	h�y��&�b=�4�w7��ݙ+�<���\�5�m4eDb��@a'��-��h�ASw�=Ţ�@�p(OD��i�Mb�Sf �0�6�p�[dif�Jj@�Z&p���^d����,�����٤ܗ�
I]���>�?��R�S/�O;��㟪Z���m���+ߣ�o�A�ٳ�n� E=g2 X�ub����;�O���E��&��;B�fތ0��1��2��f � b:�&mhpa�:�3�6})�0�Rɩ��P��I�.gC�`T�V7��^��å>A&v���whqwjW���:�ù:ӧ�z�r�ӆ�q|ΩV��Fލ4�D�w�ub@�
!B�2�һ���ajv��b^����~�U���k*U�U��k<*�Vo�i��Z\h���3:pQMA1����2L���?2+�+����D���:��s%�(������l1m��ƈ�:c^�j>C%�Ρŧ9OS^� ��}�d3	��@�����)���=�4�,2��腁�����2�F=:���}p�w���(\t=�s}zΞ��5�0�V�x�[@�p�� B.@���vj�N��K7��:���8��~Z�ZCͅy����J^���.�1��G���NJX���QЎ�Y?�����������eitf@�hmz�\ ���j��4�'r��?��Bg�?�o���+����2��h	٨9�8��d�1,�L��O�����řM��c�4)�=�b",r훞�R|�`�U�К�,�a�¶E�A}�V�D���P����n��nkE7]�~�c�%��+G��W��;=~Zx�z�^��1��v����9�n�h:x�5��۲j�E���x��Н7�y�ַ������f&��k�E6�Ս�����G�ۗ�T(�!���;ZP�R���Ҹ< O�rc��,xD"i^.�Z����鑮��j�t����z�]XY�a.�F�
:o_�0jӔ"c�I�b��6�&�P�fQl���Dk++6����Ԯ�;�mzFo�q��� �:���Å#�s�@��EU�Sa��f����z��M;�+��l� �7�F�R.iccu+;˓�Z�Sk2
Aύjbv2���z_��?�W����uhJ�A��l���Ю����~J�����p�Z��^=44+*d���z�[.x��(&L�A'1`s�5��M��p�˰^�|-�b�ܶ&#�����_��ږ�ߝ�Ctp��-1�"��`���t�S��BX�MC�U�
?ш���w��ȶrd��XPNc�`�Fcb7Nv��ݴָa��?�=|�����������LM'/t�������6����:~��v�/�K�����r�z�iJ�5a�� �ds�b�� 
�?�:�~ ��J��F�I,L��@�O��~���b����2�g��'ԍ�ūi��R�=yH���K�E��?3�	c�~/���@��葘2��b��fj�Xr�����6���+�.���E������X��<���8�lT)ώ����9i�;���^ՃO>�e��K���Ѡ���}�u�]и7Q��2X��1M�FqF#���|�Tn�N��͈���sO<I�ЬcP����"����})�h��` &�x��獽P�O7hq���X�Z%�h��O�EԏcU��(!:[�pb�y"��X3�fW>/�gi�������j5���o���R���M�0�2%�I��ʳf��!��脏���O��]�8����7�ͩ9�4�t��Q���/��n�j�V�r���/ �� �5��j\d��lsφ��Q,�~��sO٭��z乥5�A@�l��M1VއaH���]���T����z�}��1�{������E�㘞��c��,����qc���[]�&j�бX�z�d&j��iO���YtybS�hb��R��51��0�����酦ά��#��ĳ���Z��x& s��>���u���ڝv��z�Cd����4Ғ7��4r �c�e��t.y��k:o�l��|Ͱ< �F�:���QTi��#!��
��tidj7ϊ��{�� ����Ga"�r���d��3ҭkҤ�K 5Q���`�Yh������kk.a���3���w4�����y��N�g�Hb�0$˅���o�4c���U��{�F��VVVu��iK.�8�n�����PP��iX7��0Pmz��k�ǋ{���0`��R��~G0��F�
�'ׅ�4Ti��3'VAE�s�M��z`_*��	�:C������	�r�Q��Y�~���=��ҕn2<1H�O������GC�1n�\�S���NF�O��f0�Y�<-M�3�ݷ'��������T����W{(�ⅷ�С�U[X���ڭ��iS��
�M힭*����O'��}B��7MZvΩ8X��}峺y�.MA?*EKFs����K��F�����ԁl��������Ot�'�,0I��VzT��vc�
w{�|SKӞt9qF�!�s��Ć���k�/��ǰ�&�4��c�͠՘B:o��Ӆ��u�
��K��ׁ��ja���}鍷Nj��
8�����GFR2���(L#���
�5H���<��c��H��9����Lմ�8gW���~[=
l�yݤ�b���]E��n�g����G^��]�t�-�k�\����Ac��!.C;�w���=üՙoF�3�q���""�� ���Y�%����xN6�	�ʛUz��c�#�1��4>I��#u�I�_��崹����k
e��P)_U�����f j��a-��a/P�l�1�>hR�Z���s�Zр�Pxqh2�z�Ftqc�,W<9d���9�6�M����~���ñ3u��Nt6���/j�C�o�}w�"T-�.�)�'L��\�@���P
���C��i���l�L�(d��pG`F6�֢�󴾐[O��pY�����eLDb*��hr����]E�5��)(��6�A����aV���O�9j��3���9J +F�)�l�@\L�(��䝄j�����;�]��)G�5�9t�v��{�H��>2�T.�����0h������7��=�v;ZڳS�κN�9���y�u�]:�o����*�@��z�� ���f4�y�Q� ȜCȮ!�-G.&��n2pi�j���O�F���@^���� e�yAys�q����b4�<��0c
�M ���QS��@��n�L�"?��������M<���4k B�3}��,���31E�s�u���6M
b�M�k�C%���M{�J2�
�Jw�C�����|B+ݎQ��zC��M6W���~�b�nW%� �gEE��t����d��4 �o�h��� Ş�B��]�F8��aF�S\����X�5��T|NP�r�ܴ�~�����	�@�K:T@�n�����Eӄ�L��P���~����o)��b���Y�gAa�!�;]���c}3�q�
�a0T�Z��w7?ѤD�T 8�݀u2Ԥ�S2p^`�_r�ȳ/����%�׍i�������_��>��K����n�I�="B�����H��q��cc H��hf��f�+m9�_(��D�)�|0^"�Z3�"~���^O#&4����%˨��`֬�� �`1bbλ�������翳O1qc��K$>Ҁ�hh<�J�r+�Ћ��i�<NYf�9��0�cwr�3�n��"{'S�-�'a08wT�5.���[���xXO=��'�3�)���^�O�u��혉�l2H���@KL�������W��M�D㘏{*G��Z&���N�M�m�ul���`�xR�15c�q@)�/qfc����Đ�>a��/8��I��w^�8#3�+��]�^��*Tb��G�"QN�v;՜a����"�=2!xk��V)�9(��2�\v ���d�׏���|�n����L�f�MD�$�����{n�΅i��`<�d�̗�EO��SNeL�$�[����y���9���3����@��1Zz]x�����0�P#��?�k&:��-��w��w�N>����ɳUL60ķ�Zۛt���]��\�D���ϐ�i0�и��ǚH���ok$��^Q	�q}��,\Խ�y��M5
����P��������4�}����f� �7j�W��5SQ�C��N�i����dC�Ɇ�'�[�ݣ��R�j��08��h���[]��� �ј�#)��`��Oc�����LE#�	�D�d��z��,�Jnq��z������Nd@LWʘe�}��%�5�������ُ�'*)�Y>��ڝ� X��"�M���ViسS$��f�6�R��2�h0�N%�LcQg����H�P\�;���m~�Y38 �;�6��6E�03ӌ9_T��Ղ��,�����ʛ���XӤs^��t�n>x�����>��(f>	�ߥW���*L �5�/-ޡ��Q1/#SXhRl�SS�*��j��2M�:�ٽQQ�B��)k"�>�'��M�ͽw�ą�s��EÃfC�����-���<@S���FЅ6��0�f��a�BL*̝(�y��4��CY"Ϝ}�[�#���Ȕ�u;37�s&��#��C/Y��+�4�4�|q��g�v���OT��\�xsӚ�(��JKc�陼}�<%�@�ޒQd{r������>;��=A���)6SA��f�D�♘�Da�o�i#Bl\�;��ԨA�ϭ{�o��LT�~?h�]&��L���h$J. k�.��h7�)�Ǝh�cp�>���Y���O��9@\<���XgwϢ $@ۿڭ���hl�����TEO��f��g    IDAT�����U-�ޡI~�VkC3�Y]�ޫ�s~��{�=��8 ��6��9\��S���)ӹp��^�X�����^��L<qH�U`�B3�$�gĴ*�%�I�So���[O�d��D0
�4e(�?𾆮�����,	�������`��0ô���?�u�t[���p}n�)�t����+�5�|i��>x��?�=G}pl��b,�H�m���q_/���;�+�GrE��u�]��W��[߿O�M����� ��.d*�.ф{ ƥ��jL�K%��Tx;�&�?���u���=�eɃ���pVMЬ2A4c0=���t�/��hL��h��w����dp�>�w�*��<�r��U ��p�	 Ѵ����AM`v��ek=i��g� �˫�n�1�$i�:0a��#�549���Ey�xT����V�Q�?���#IU���i�ݍ��؇oҽ�^�B]�N�Lw���u{nP�8<:#�f@*�K�4N��  ?��l$ �'�,�w����چ�,�����J�n� ��@c��\��JT=S���tNq���t�{�Y��&�K�fu�Fpb6�,)>�+�;��
zH Z���~�|f��k1���P���E��y	�av�� ��ꉌύ4�a�_�6a\էT�.����w���㜪����ڿ{���f��˜�w�F�Z"GDf�q�4�����T�g�erX4�"��Y[f�"�3���q�Ɍ�Oc���w�&�Y��;Gv�����d�~K��;c��L\�����k�)��9oFҘ�G�Cd�Ǝ�6p��En�;�����՗�B�5`$�mͷ��<3t�Pȁ���7�Zo��˧��w��3{���HS��Xڮ��m�����)�q�:x��ڻs��~��=��M��J%h�53ީl�a,�4���c�?�k��P57��`Ԕb��S�8����\���aG0�SC�&�64��~ٰ!�8C�$�/�8������s)n|��6���D	�g���d�#��s9��'	���'�b����&�J��V+O�C:��1�� ;x)��n��ה������K��z�ͧ<T��Ӊ#���wݪ��r�v�+�@�{���X�c�GN��I蟥�����x��elhF�݁ʸyY8J�7rk�"}�f�k�����M8���������Aq4���D�6*ĝ> s8!��

)w�?�/��-]	M����2�e�������
�[.�f�N����ʊ�`��7֛~�ٌ+����C|gA�v���]���-yjc�tg�Lj�6U���aBT�Y ���g���GN��|�����'nӎ�%;�q��^M ��R�/���r[��|���;6;���<x�)䍶чR�R��d*f�����S#���@>��	�x� ��,�T"��=�����I�D�8¹ȵ;���1z�$&kM	:/]4JH�i]��j%�2��7Ek�d�sa>�6�S�RU�^ѫ���;�Hgη�>mt�Ԙ�)W�>U֝�Y��t����
��J���7ݐ�
b$��i�QИ��+|q�2��������C��C[o�Rކ�(�	2�	@�Q���&����5�N�hn��8A	�Ind�mQZ�:����,ygi��cbU�����
1t���cXb��1�}|�\�u]
�!�th�X�������^�u�.��K�h�+�a9m·g3.�������t����촆�����{t��Wk~v{jl{6p��m4@��g�5 i�e�	�&���	0)"!�w3��d����1��պ*L{z�%B?{����2�9ئ���c7�3��s6M{cV�%���W�}t��Asd/��g:M�M���"�Mќ�����6�q�[D-�2Ma��P�m��Hɦz��MpD|�و��iS���a6a��^W���~���RM�jM]����z��gԧI g�t{C���O~�K��ڽu�w�i�3:d�嬉�� {(;`S��L�FGcӔ��V���i�q��������w���&;����A��9�u`X
D��>iF�1�� �X�,ZW�4a���S�0����j��`����"�0�'5�Яx6�nV��Nq���  F��9D�X4���z.z�RA�m5�~|Y_��o�����Y�_FSZ���͚���R}��5U����ii���&qUc��������h��Ϭ����uD8oz���3�<�g�l�n�fW�:�1\�ǚiNkn�tF&�ŉ�ÎF>��	���[��e�<�A���Z�n�y��4��:Ω`�x؜h䶭�K�g�bՕi5M,��@�閃�A��jDTZ�R�lM^6�I��x�9bgg�'�1�L�3s����=wɁ���ӯ����y���ƺ��ku�-<7�-�\rx����p?��E��E�M�^���+<;�B�k��e���w���Im0%lP�s?0�4.��D^ESH�R��"�����?�	���>Ӡ��M��Ԭ�b�OL��2 � �=����3��}fЧ:L�\Ѹڌ��I$fnQ�)����[�;�¾�-��@N�BY�J� ޹]����cO>��V���ms�X[UgsEӍ������t��+5ըx�u��:0�1��^6��Yo�ǳ}-����T-7~�n�1n�S3�<���k̾��g�B�iΨ�f-EEK&�k�F/��ЧMbe��`�����5�V)k�̻4��?�9�`FVf#g˜z�O�������/��f�(i�������»�Q�k�+��W^U�3}�pd��X�8">B/֔����Iiz��� K���u�7�j:?�?�����=�����A�ru;c�8����W5��(ו�w��4/�� 6y��,x��Sc���Q\�o�~��>0YLnS��)�	
�D1�B�\�M�͈x�g��ƭ�����A���	�=?�V��O���r�M-k�A3UZMC#�ԅ�]h	���"$�Fs�Xx
�5�Җh9λK�H#�	�zhت���o��U���Q�����4�s�T�V����z������ә��ڵ8���������n�[�m���\�
G.Ĩ2�F1�Dql!���:�P���7�ەȄ32�F��5h�ۨ��1�Abl�d������M9��B�1z}�!��1��D�Tب���&�i���q`�Q��
�?i|�{�JS�db���p�2�5��ɗ�Iph
��6;,�$���s�` �+��G_�w��`D��jK���Y��Ҭ>��i߮%�}5
EUK8��~��E�xB��Gĝ���"�'��i���8 �Ѩ�NR���{*U-q���k�F�?��I��-!Q���)ԓ�4M<K��i�P���آ�an�N����f38�d����� ���R)h����}x�^-���3tu͊6��itP'�IK����w~��}޿CD����&��Ck����jU?{�i}���~ W*Lz޿v�ث�n���wMlLUC�E4��D�'�{ WICmĚ�O�p&�#Bi�e�FGL��Xt!���dz�7����z����o�YX�����K/;�]���ڨ�~�����}6��F?3T3��H�w�{�h�DiL�w��)������u��؛o�%eUV�u�ڳ[��iuG1!p���c`��
�������
T��i���5�·��x�l0�C,�a\yGC9�y�9��}�]���ƺ��~�K����_iåqw�	��'��lQ�r�+U�OPœ0̓T򟬥dz��+�KŚu�ц�����Gb�=�y�A���'̬�>�Y� S8f<�����`��D1haP31���k�x҈�����Ѐ{��!k���kB�6�j���f��;�5�v+��d�R2�X�Lس&+ݟ���Yg�Pn8�ƥ�����͚6Gc��?��N�Y���v�}��u���v�����Ks�����Oi}eE+�Oi�l]ۑX�JC|,�L� +���7�W��8<s u�M�f�m�3c���Z݀ѨMF]��XD!l�64@g�3<�%�����	 5:��J.l�-����,�H� �D��s�d�b��Ǆc��X�q^�͎Y:��4�ۗTk4Tf:�D�1�1Fh������J�(��`��F��,��idx%2I��>�xB޹_m�Z9����z�W���XS3s���r�����������Z�&�]��� kB�� �Yp�/NS����S�|Z��1S$����ء)<a��ԈmecK�]v�G�Cd'&Sjߑ�XDm�+��7�L��D���V��gr׽Aw��#AJ1t1�.����+�[ܐ&���T�� (�t`+�z�����ϙ挏vkSs:����~����[*�ɘ�I�h��s�QoCW�w�n���.�d�!
␬���kk� l>�XU<v��o+ԆU�^�	������ܮ��c�7�r���܄s˺Stk?�aC�љ\�R��RPk6��#�Elw�R�R��n��k�0e�� ���!�W|��H/ըM�\ᵑX��?�ĺE���^$dC��|6.�.�tA�_�ۖ���Ԍ�c�+Z���05�9�S�<V~����������2�)���xS��H�Sҹ�^�����>q��4W/�J�;��.\h�����F*�9й6�Rp�S��CgSa\iJE
u���`�k�-�N�'�K��-�>iԝ���D$�ޡ���"��~P��.�nb�y4@��Q.�5��4�����W��E��!����E�Ơ�Q|���7��`bT��C��;�6c&/����=hn��xT���f��=s�]�m�J�Ϥ�Q��X��a��~vH�x�%���UjM�~���'�׶z��`_:[�~Q�{�(���-�퐇��E�ψk5m��1-�am<7jҾEz�1^�3�Z
*@��d-�t	��(�)���Sf�u ^I�6F7���kó�R0��P̩ȅ?��1�����L]�빐����؄��>vwc���7m�6���"2<U�@Ǽn�TP� �gS�����8����~��G��/8?�5ya��ռ�M&�E�r����6�\w"�ĸ R�x�+陈E��'�쎼+�f���26;�3^���c���8���ѰE3XR�RP�F�4�I��P0�)&I^[E�/e�+��ͫWNh#���V�'�ma�5��Ơg���t��A�HK*W
�0�Z]o�`� ��.;Ŏ����1�`7<�)�M��;��C�ʠ��P6a�'�oж!{P^��H��juۺ��K��S/聇Q��U�V�'?���pV/<��n���ڿ�:4�MB�j�w��^A�ZPw�c�Z��C�'�d����O�K��P��	ΐ��v%@'�J{����k������=~�������/��okniɅ Yu8�u�"�4֮l>;	�&���wȾn�C�1�1���u�ܘ�{b�
��s5���z�����ڊ|FgS���ů���v�=�F��Jc��'f-" ����1�e��3�t	�&��^�i8�H-R���s��l��`O8���N~��
#�y�Μ;m�������>���tՁK4� �J��U�1`�w<C�3�J>3u�b��)>���ǹ�1	=^��a_k�6Ԡ������f�Wձ��{�S&����Y�(t�+X��PL���Y6ܞް�x�����2q)����;j�`�nX�X	�g�Z�y�pcsS�2�����D`x	�;�:��S7�����et03��Xʝ^���P-h��f��:;����?�W��W�W����ʺ�vh��j~nZw�r����Ο:�͵5�=Sͦ��i5j5�'f�v��kg'w�͎�n�eLh*��L������Z^]�ٺmvV���<�����쉓6BA���M7��eW�#����!3�1��76[�WQ�Bs^�W\�D=噬���X�	Ȏn������](�E�p�^~�Y��"�FC]y�>x�G̀"C�`9�s�隧;A�j�|6Z��B}�$����l �������h+�8_9��oߦ'�|J�>��.��2���Z-/���W\����Ɇ�g��&&�Ϡ�հ�m��3�3h&cn�m��_��В�_f�����`�2��tSgO���i���d�1�D�v�a2�`d�F�K5Ԭ(������K�s������X�֘�-�%4v�S�~�߲W�{���7�4��M-C�nM.QP�$E�8\5��7���[h�����GNd��ܷ��U�L[�aOS�)S�񁘝ۮb��=�K=���f}�S&���`��{����[�����
����3����P	�A����\��(E60��̧��偝C�+�`��ڃ<e6�0!t͇�x\���A'���ͮ����i��wJ ���O��C��RP��G;�9d'�	?���|bKq��bl�
�k��6p�����c/ l�Hhn���!v�FdH�����sY��X
>?�
&���h#B��0pp�$��u�L�yM՛*5:��Թ^˙��ږ����VFn�̔���_��d\�Q�ذÌ���C��V�Z9�=SM�s����}�%P9'�:�ґ#g��5*54ʗ�e?�ђ�0���0��"�qwLW���Z�����bB�A�������r4,��VF�c���������t�J)*h�,�����㻁�{��g�T}���f��,�4�(��b��rnZy�8�c�`T�2�����lt\?���*e���]O��4�s�ͦJZ��"�/��B1��ˏv>�	�+��9���gC�p~UW\y�>��t���v���,BBF&C��(`X|�q�(; 4eҀ�q�r?L��M�_��l��Ha����o���lʑL	؜)��GQ�p[�{�$u���OИ.X�}+WƵk�l[]��dѥӊ�����������p	�m�:��6L�a�DFX'B�AtLIp~�i�C�p<4T��mRB#ȽT���L�\���FC��cz��+�W��w�~NW_s��z�:�|V�sS��6�q'��%7�A���4���\4w�N9���RP��g�?l��˱=B
=��ٴ�4�"nG����5k�`41�����֑�h@cjC9\��F����cB�;~^��L\��t3�m��]F�cJc��Ŋ��Zkkbx��@;��S�Z��ƚ�9L"�+Y�\R~`�)P<�p�@ăd��i���w6J��,�8��j^ghS[����Xמ�������Ӈu��[ڹgI���EgN����\7\�.��r�ot[�G�P���s�ߒΊ�������:��n89�lM��f�-j~aQu\Wm���7Ԁ&j>�'��1��GN�[��:y�e�y83{���ſPcv�6�]�MSӳ�V��k��mN�(���V��u���5�57(M*�u�O���qO�>A�Cv4L�p4���}z���7_���Οq8/{󶝻���ۚ߱G�b��J���n�뽞�8[�s_�7�L�"A�>T�UkE���S����ux�EM�2��R-��i8)��mNO=sX�r^�N��cǎę�u�ǚ*���ܪ��x_iY'ΟL�͌H�(GN����(����v��Q\ZK��@Q±6�g���-T�1$S��:�7pӍ����o�ӳu7�T6>5p�6�ؔ<
s7[�C/h�����8���W�h�v*M�iG}X'E7��ZU�3�y@�Y;ih �|�#�v�ئ;q?� ��d��[�h=2�2���N�!:
�&���u�3Ks���깗��eW^�GB�ίhi~�)�s�Ӻ��۴}q!�{h~ae �����+rA���m�TQd3�hNӤ��A�?V����ɾ��g_�Fȷ��xR����9�#}��_�ˇ����ϽFU�}�s���냢�/ůMM�������[[	#�V�y=[L��y�p9��{[�0��dӬM�H(�w׼��A��;��&�HX���������}֒�Gc�C3���t�|�����'�(q��4��^�w9���`?�j��܀��i�Q�iaaN�?�~�������8#om��VkS�]s�n��:U?��5u�k����q���r-fM����;�k������c    IDAT;m<��c������KSՊ��O�����BM7�z���g�&@ޠ ��`����ׯ5�9k39�d�'m�W��Fc7�f��&��h�%u�=5����:u�tL�4��`M{/ݫ�{�$Iv��h��L��&\k&'^�� m���_��焷�8�l@ n ��Aj�`��H�TSi���<|X�|�9ml��l�:�rc}��uS�<�-�^�o����ײ�FPE�{9g���h�->r��PO9�����L(��ψS������1���j�.�]��>�n��}��֦�fu��7���;T/3\����Jm�C�;4�%�cy�L������8O�ȳ�nD��`�s���3�T�K/���o�3Y]Y�FgC{޳�o�V���7�U�e� c�/������jbn�%㺨DD{�-z  ~��A�pv�7@~.��g�w��R���V�i�h9��j5�?���@�����'�}��|s2,L�^����JJ��F%��ښ�/�飷]�+.٩�ZQ�>{J��}S�ڜ��Yg�@c��L�z��be�l�JJe��{`P��5x�r);�ڳ�Ӌ2��э�z2��QyhdgQ s�x) ���09�4e%���d7��m7�Ġ�0y	�yU�Q]�!�`�)%0bauԬW|]���=�xz�,�l0�Ģ��!��[T��ͱɀ��:8���Ҁ�eΈfЈA���aZV�/�������W^�`cC7�|����V�^q� ����S�W��qx����e�������T(�lC��E��ԍ�؇�uja�C>c7�	�5{ӣQ��`�9:�4�*c�g�����#�.��8��cS~p�����๛�F���Q�^�����6��l��=h$6{�#��4'll�%�[C�95�S��4�5�|�H�Pk�!eNTL��휼B�Tx�;��T]S�i�����Koj�:���5]8w\��q��r�=s��^�n�]�K��ɣ�L�\��	�,�fl��<� C��E�͗�P�gy��:ؤ��0r��'�g�ZNc!��n�I��:O���K���ǁ���+�w[�d��tS��#\��� ��B\���ڽ����������M#Ϭ�B����}Hs�wi��6��L�JƋ���P�6y�2h>
�s!�vd����n�m���L?@y<��BO�.K�JNbGKKKz��C:t���{]K{�������G���߻_���!8p��71�0z�5�4zĊ*�on���Sj��h��)�9~L��UL��kssS�zU��iM7�433���ڵw��w̫\��y�W�5�E;t�������DG_9�>���{��o���֜Q�?�z���D�7�>٬�U/��������ʅs�6������j�Y��҂�4�mZ�F�kl}sE�������}����E���+��/���z�������ۯ�������.u'����&#G�����>yV�ϟW��R�����iTA3����h���ڱ{��e�[CS��pq2֨�g�!�X6Z���_�1����'�����d���빒��f]�k���^m�Q0�>z�V)�T�)6��r��MmgB��Y4�ך,&a���b������Ç������UKM�c�޳[���~S���A_��b=3�Er�*S�_�cHB28�5ȫ�F��Qo�f�c��ӑ#GM�c/oo�����}��j���ACa�'���e�QK��0���d��d���p�ѫ՚n��q4�uj��zb�Ww�a:�܎%�Ã����_�W�O���Q�;w^K;,Y���ѝ�ݦ�BSliHh>�\�
��Y1����s�T��TC��-9����z˚;[9p.�����A�r��i(��Ҷm��r�Ɵ��?�D�ڔWcnN���/�ʫ�6]�"��O5�?0a�UA Ԣ��v��vT-�4"�d0Pcj� 6�6S{�h
۝�?+�*�`2w�{��ГO���5�,/ǽ�U��{>�{?�Ǎز@�H���D��s��u��M�:}�{���nK�
jT��p����Su�����r�7���(�haqA�|�i=����߾K�Ξ�^A�t����ޤ 4��e��P��C�z�
9zhV�B�n��}���/
k���L������܈�_/�_������z���m�gW�ܶ��>�1��Au&Cu��3����I(�?i�_N��;�W��2@9;;�	n���7� <J���`v7ʫZ���C/���ڹO����>�鎻nwm{���BmeFIH����GY4zB�Rna2Xcj'�Mt��W`����a6]!�3*|
����O�O>��`nnQSSM���E2��(��ߨ���fu�1��2,�sN^��=!��ŏ��Ɏ��� ՙ
B.j�0x�-�}��0��y�6�cG���7:��	�h�%]����c�[W_�O��yn�����n��I�q�'�1�7���)�-SK������"��N��?��~~�Cj�n�MR�*��_�{�����`~�adj_-���B���5���]X ��=�S��W�"�Q��(L�tC����Ab�~٣��U5.u|��VG]�mVG3�j��pU;�R�����@5Պ�l����Z˚�k� B���={��ޯ�\�]/�|N��9�q�����@�(�-pvS��(��r���a�<7ϛ=�r^*��n���3Rd~$U@T�d�lH(X�\L��fU�6�4�ȉSU��i����������pb=��hml�KS@�a��Z#>���������3�#3����ʅ3���'�X_�m��켛��8�p�0QeɃ���pBCӖ>ΞOF��4:}7�5�c��!��# Ɍ�g�������V���҅��5^_�-7_�O|���j�Iz�Qy8��¤ȋKpŃ����j���ó���1o�D�B�~�8{4R�\V{m�T&Z hs��5��B�G��%�D�a��q8��b�e�����*W��b�1.rc��P�p�뙚c*�)���ƲN�<a36^PMP�K�{��͆Vz����v}�9)���G�4S�����������3�8���7��554����������kjԦ��C��ȫGUe�t��1���.p~���*7���oݫ��������8t��|�l�^�*"t��v��4��B� ���\%6�������a�T/լ����}[�>�3���U���ާ[�KkݞZh��_9��~'�e�f�b3Z�̢��0O�j��@�+�6��b��H�rQ�]�SG^8�o��o��[����j..����w�W��S��,G�_�7U-��S_C~��sMD`�_V�Z��̔�_�n�8����tH8��za-N;=?7�G~���y�66�57_�W�z�ȫz���t�=�j������3.���h������bEo���Μ|[�O��������	���rA�����9r���}�^]r���"�,̫X�Q�PS{c�=K�Z>~B�g�c�?�QS*յ������D��mʕ�:sa� �� �)���=���|Mo��Ϟְ߶��� ��Ԋ���/.hq�-n_�ݿv���o?�++j�lS������z�O�o����8w�4X�z{.y���;������ˮu�b�FV��M�x�u{��ڛ]��mOm�@�ɵ�Ǫի��ݦ=��k��K�s�EZ�NG�K|��M,����O<����]������tQ6S�Q��@������}�`�� �>� �#�M����/�%vC��Rf}��\)��`�>��s�'Oz8��5�y�Ï�NO��au�[ʕfŁr������}\�ɳC����K&[\WhK��	\V��'�g&P�~�fN�8�j1e1bL��b�rY���3�θ��h�B��|To>��4�fS�f�dX9�q.Ry�(h��Mw��"�h��X��MS�u�ĸ�0\�Z��:��;u���腗_�U׼O�?��;sZ�;���N��;�������* ����y�)�П�+EMՊj��N�N�8��'�i��9O��ͱ��K��f�-h�ܒ���k�q�?�d��@����i��j��?���|��i�o�g��ӟ�u]y�UZY]���˫a̒D@�~W�ϟ����'�6/�)@�)�p��b��=j��kjzNS3���iJ�Tr>��vK�v�Щ�o���|�dL��e���鳿�yM���sZ�X7�̹433��q��i����z啗���������bE�jC��5�{N������ڵw�j3�-��3j����N�4��/�������-�Թn�wn9x��,a��w���5g�A5�q��Q{�=��u��W����b��%K����;��n�������f�ͩX��i$���Y�����G�7z�����w����S��[������ku��h�\2����]&u �GS���NG�*�`j�4�F@z��5m	QN�RU�|Mӵ������7���S<P�n��3_�������va��^
ֿ��IE�7P�`*�����i3��l^���)��l�T�:�r��g�> 2�kuu}�G?�/��kչ�%�L�jum݌$XtS�5�y�ͺ�ڋ=/] �2�ǹ�=*b߬!.�,�a�յ�67��6�;�V-{?���-������0��lRjԧu��c��?���������ܜ���>��Oh�v&r1յn0��2�u"�:��6=���3Z���%�Sm*��F�&l�"�x�sO�M�*��O����]��:��7�{Q���q�sޣ��KOSR�ݳ�7���u�>{N��+�<�H�TUmD97=���'���F���P������I���k�<�h W	���F{��`M;�9���w=鏫*��|��7l���y�U�b���;���tѾ��u:w���M����QI3�\s�y	MK�@�J5��_/�1�Ӵv�#up��n�)xх��g\˨�ҙG]4���)j,�..i�%��6\�2�����Z�p�2� &�H���2OO5}��⬮���4w�k��Fhz�y��ȵ�;{J/>{���G��Ҷ�E]~�՚[�iy�xb�a�ɰʦ���@�z`W?,����hCO������U���f7�B1�2�f��Ա�u���j�;#����ޠ�~�Nm�DcL��DT���*�4��l��F�j�v���9�K��hD���X&�9�R#��T�z�t��5h��fy��욫�+�t	4��4C�q%%���9��6U�<��`i�`����v�d�M����N���y�Am�9��ZG��Ds�w�_�����V'�W�Y�}9�B8�BC�QE(
PZ�|%W@�lH�����옛�o���C�x�5Σ��X���(��kG4f2�i}�����j]t�e���>3�����ؤ`��a ��ô� �9��^��^����M��_���Z��힆�K-��C��l�Ӷ�%M�ͫR���������L�-�N�������O�y���Tj4�����n��#:���Q���.[<c�f�����������Ar�gz秧s��s�`�9$��IQTXI���w����������[W>�����wVZ��(R�H�  r�4�� �{:�ܷﷱ�bQ�3������<��!���̒��M��L<�6�]m����Ŧ�tEq���ھU
t4ד����O~�䝫�dQ,�m���o� ��OBl��Q�Y�rnHmH^�ܻr���	��ʮe�	�~[�՗����#jW=V�P
r�@6/
���*q�9Jy��.'gO�b��=��6��o�Mf��z�����V��0f�Y]�E�V��l���
ӏ239���#R� �L��es�˪ϴ<'�lP����h�����L{_���xڰ9�H[���"47�G��{fG/Q*��6A]� ���GX.��� F��Bxy��GL?����$���t�j}V !Y;��0��n#v��Z����_����͛�x��Fc���������Y��THS1h����V��e�D���&5,���x��6w��<����b5G!��lժ�b�gU]��������5�3���ûih� �/�wJEe>$��Ao�Q���[�h�na90υ�G��o79��+�K:vm�Mw{����W��\�Oȥ�gy�/r�2+K�D,N8V�̩dF-3E���,n7V�Sent��MnQ6�yVWWUV��t�s�9u�Ν:I*��X�)϶=�x���)�eD>�6�t��Г��5d����B "2@�5f�����1q����-�l��(����%�(��T��~����*�%�[��țo���{��V.e�Y(�,�d�(
���F�%]Ȯb��f���#�j�݅�j�h�T����
���ʻOH�:�\�0���+���������q�F�^`qa�Zw�u�\<��A�z۫��B~�)����ٖ��x!�����S,̎X�S�OA.�*�a@gt�֊���[�Hw�Z�׮���P��0Z��\ΦSJav�����ȩ3�}-�{sm-��[�m ���j��׸����011ʝ�7X^�#�3<�&��RH�a��;Vn_��6��il��[ߠl��7;*3X糲2��?�׿aqf���u�ܻ�7�}�ͬ��E�����j"�r��5n^�ƌ�VՈ��:D���\(%dF��P�i�����u�h����0R�hJ%�.��n�|�,��_�Ήo�`s��F�jȒE���-��>,�/�XD�V��*�G��r������(��n\�%�8M6�v�}AgBoua�AY��S]�����衾��ϥ���� n�����?|ʅoN�
GՒ����so���]�D%��BC!�U�<"ł�IG��,�ͳ���
���Z��A\@v��ہ�����&�N9q����I�������ʹ�|��O������u��/�k�6%��u��ȝN��F��P�`0�����Z����t��BC�\��Q�،�֍֠�]+jtQ�EAT7Μ�!I�Â���?}ŝ�����t��;\ē)e{ψC�a����l\߮����
]Y�cD�Aj�j�w�r���� ��s�Ba��d�	�M�r�}�mV�hij�崪�R� �����`5ۙ�Y�?�Gf�)K���eh�&^�|>���V-��ryq(ɹ
����$����E\��JW����Y��/�O��]��v��eZl�B3�r��M���gʝ�7��o�cӾMl޵�ϭx ������lV@���Y�����fa~�x"���U�+�n�6F�U����u4��45�ij�Ip��(��Sw|Y��Ìޢg:�J(���$#,wmy��d,Ʃ�ap����/��j�+��|yr���H��������d�R�o�l���`T��JQ�OO��+S��Z�ʩ�(�xؕ�]z�j4�V��r�T��f9P�:��P&�؈�!t���K�x8z��{�H�VՋOԠ��[ذc:��H:K�c�ZN��g��ȿ/�N�M��H��J@=��������**\8Z&���S��^��l��#�7�(��Nq��1�3Ҩ���M���ؿ�Ɩ��R��R��Y%o)o��s�ؙ�ʒ�r���"���\���."��U���
伓CF�y6/�C-6����n߸Ili�b`�����`q�kŦ#�ZU�o����+T�����!��ul����e� 9⩄�����r�̈EC8Z��m3FΝ��ٳ�WCBZPǚ]���ܳv$X#6%�a��V.)�񒋳��-F]v�����������XF%s��n�U6�Z� Vup�,$W�8r�0��I*������[��n���)*NP��R�̘�V��x�l8@1S��(�E��	�F�=V��ǋ�W��fU�>��TX].5��N+��bu+m�r��%&��M&�הH���]C[g�n����q�HT0�O>��0he��WarQc��hT);�-���d�1�ٴ~�Rʺ"�{��Z#uMm���%�����o���L��Ĺ��p��7$B�*�l��w���}O3�")��+E���/��)%\%��B""��ϥT�C,�I:]���6��mck�Z?:�E�M���,f����@1V���<�yA�O��ܻ����%������d�Wf	c������Y�� �X�x$H&Q�z��7hUެ�����ںz =@¿�ֵ�3ZI�Dh	    IDATg�ĒUEV�oy��&V\&#�|����,����������\�z�CϽBKk�|���k$$_,ZYejb�G��X�}Dre�J%�V/
yY�kꌬf{E�ʪ%��"v)3�L��F����������J{�Z1��q�Y����������*Ӈ�E]� ���_�M� �,V�ʮ.��rc�:S��(��!y�j�D1&�Ҫ�Gr�%u�S�7���A�֬[��/�Bcs7o?df&DW�:�o�r������4�BJm*{{���&��xF�a�:���p���ϓ\������d�
*b �8Y&T��d#N�TA�%�Yi�\��=ϲ~�NY�#k���%dJ�٬r�7n_���ɩq�^�� Y����9��Yښ;��cU+,$� N�$�;D�p�Z����C��Y\Xd5 O<ɒT�e�f6au:�kj����Ξ>�9�(���B&��n�P��q��q�;F<U���;����o�Z%M��Xl"�$f�TF5��E5��,+�s$�1�)Y|���$j��ᠥ�����f��-�R@�5YZ���)8Yt��S�\QC�r�������޻��,sM��^Z�\�'�j�$+�&�)���w8$.���e�pc�8ihl�뫧�W��!�V�9,j�� +T����,�R���ӧ/2��1�vl���S�L?RU.������>�����e�R�j���J�Y4ģEn^�;#��jm��JR�'YZZ��G� �����BNlc&N��Z;{�k�T�XW+�Sy��<v��~�.}u����1��|���g��MdĹ�
�c�,q��un^����#
���/r�M�ήVj�~��C�/��u�-<�t��@S{��\�z=�Z�J�h�����o��_1?�X�z�g�u�v����X�fEf4��p�ՕE��\������Y���I�T�1
��a�PuX(
��ŏ�VO�����A����݆�iQàd��m!�ZQ�.�����ߨ�H2�T
�(�۷me׶���*�G��ŚW,��yo�B}}�*7�^&8��b.��"�Y�H�LbCz*B��
�ބ�������܎���������^b�4&����/?>����&
������W��.}[7/�I&2j�/�a��B:���;L�%� ����"A�'�<
��lw��X�8��h�h�������թ��d�r��w����?&����.-/����ReYP�U�b �M01>��{w���T�lq�)������K�GE+|�-j�ћM46�q׺��X1�>w�3.�B�l�?����1�������%++K qXmf�ڻ��M]�ަ)a�O!��T��9*}�V-���p��?|�l��D��M�&�z7�m�6����Bk{�-8�E�;U�T&���v�.G��O~ɣ�ջ��e͆����kt�{՟K�T���8β�L�p��MN�)�N:#�N({��x����[ћ������7����⬕э�a�����6�/���o?ayjV-��>v��Χvੵ+�Xl���	fea�3�N2��!�s3$�a�}��ɔ��V��\����a��ns�p����`æ�����]3#��TkkDQ7،L�ri
�F4<�i�,��b�z�;���J�l@'�?�D��g(�*�D� i��>���k�����H0��T����9��ݪ�ET7A�h:#�H�b:E,&YU���)$#�IeȤ�x�~Z::�:�sEe����dd6�A9����kܾr��Ҝ�|��k�3�3��)�:#�X��VGV�
�]�m7�s۰[�J��&b�Y��S})n����f��]��d[RK"�#���0N2�Q�M�ֈ:�r�X^���矲�xByw���:8��g��vF|�rq���J
�L����n�T"����0��HI�qF��k���S*I^J�հ�إ�b"22���D]3���Z�#2��};6�g�nRB�қՀ]E�W�o���N�)�J���MW�L&�r����e��tX�5I�1��2b��ΌEo��/+˅�d���s�?���*q1~�v?�<y���`�m��Ϋ�(�Y�b�:X+�4u���dI&���曵X�|��
����ɊP���ꠐa��rQ����{L)&�2k7��;�uXI��hK`�Qc�<��V�F�VB��>$[&���(d��N�lXb�0Y�66�=��֮n�(U$�%�K+�Rm`ˢ4W�Vv�^���1�85�D������3K���ڴ�CG�$0
ɷ��0(���JXK3��V�fI�ȧ�TJi4��R���d�6%4R��ť�Z��n��V���q��)uP���R�N~�FΞ ZR�.�f�������,�S�z�F�BĎ\^&0?�~�z�n2B%�2� ���3[1[=�.Z;��_Gc{&�M)�%I��65P��y�g?c��e���Op�V����$���^.Q���	"���N�]Ya~��t�b!�5�{Td�)Р��ن�SOsg?�C[�����+�Ig��ۢ�x�R����/>��;��)�YS��w��w�����<���7�a0�н�9eC�eɃ[��y����&"�u9��v�Fmi��
�W�e��VWB��btP���T4��7�v�^6��l���`��?e��UU	P�Xh��w~�c�Y�M�\�+�ܸv���G��S)�0jũ�Q�1�C��P�I��� ���d�t^�A�>1�04��������=r��4M�}�=����?'�2M!/� 4�2��cq�HfJx}Md3�|�5�^ǬIQI.�+Eq:$�![�(�S4&)*�ʴX0m�,nb��h���M{�v�z��۰z��Jb��x��D2�dt�k��p��u�ݻY(�ʫ$真g�}���f��6A�+��X���9��#���/�`~a�Xd�h$D^2aB�TN�'�ayIL��~ڻ{���������*�� Bd�Zk�s��Q>���+KU�F�9�4o���j_Ȟ67���5��e��(+��LO>`zj�ե
��3z��ZR�����Z�;����'���G]��BQ�E�y�.��_����F���k�M����޻G����*6P�Y!�S�<S�S�=x����s���[ȥ�H��U������s���J��:����=�}�.T�DY^��Vl'�h�e�7'/061����\9�̣	j]b�b3:y��s��RL�j+iI���/Y����=r����x��[�Wr�"nݺ���#d�Bh�*-�XV�.K�������L{� C�����V����v~��_s��Wd��(Y��:���{lٲ�L*��j�j�������}�xh�QH�Et�C�[+��Zb�A�ۺ��]�����VYXMQ���4v��52�q�5�6b�;Ԑ���U�����Y����f�6o��ko����r���]��\:�+/�%��Se�/K��&�I&�W6W�P0H,�$�Ւ˚��0;�q��i�Y���u�v�cu[I�bUT������	���u��Gc��(��;v�k�N�"e� �����j���_<w�����q�4،e���Tݖ,�e9�g	G����:O����:,.�m�t�顡�A��K��Ǉ�|��p,�;[x��oѻi�L�T"��n��l<ʝk׸t�����R�,�aqv	�F\O�ŰX�-v�.v����(MMm�u�R�Ф�br�g���|������gG�g_x�}O�Q�U�&�m��g�~�*���fn��OI3�P>��T��rN�y���X��ؽ��|����A��l��ѧ��YI���+:��ݧL�WQ0n.�T����Q`2��Nvo��*y\��*"n���O�U(�<�ȝ7�u�*�����iqRp#Y�HnY�H��Ŏ��@g�`syil�������|u�꩎ǓحVb�$���_2>rM� �|Y�y#o���J����������n^�ƽ�#ē1��OK�V���(��N�B>���^9j�8�Z�i�ꤡ�	�K�5�l5\������#��*B���6������㲫YG�{�\ONL(����7���TT��
��-��#���O��Au�W�z|�~��1��W-V�GH�U��DLh-F�D̦ɉ�T�ե�EWB_JV����I������Y5�(
�(R��W�l�>�B]'=������ry�ʠ�3W-����pX-�aH��)Y��Yu�e�Q�� �D���V�^�=���5�k``h��5�$r%�/�V�r�N�C!��u��)��)K��bc������!+�$5z��Z�U���r���\�T|�t<D:$�W�<*�%u��űc����Q}c��&�"1���^�0����"�c��=�x�D޹vϼ��zأB�b��@Yg$�ʐK&ȧ��X��xt�d"�l��k�XWe�*Y��n:�{p��c��*[�t�I�R6��f$�a1;c�޹Ktq�Xh�=;�p��rF+)�ˈ���v⛖�f�7K��eRd�1����
���X�B*���¢-`w�TN������^�V7��Iy��҃gU�ZM����+�p����j٠q�����l}�)����a�b������5a$o"���(s�'H��)�(�BJ%�������ճqxm]u�o�5�+���e�S
���㏙���)t���|�����(AT��K�cD!"��Dg��=$�X%��G)K!L�t��S��\���=����n�v�lN��2��T��h��rr��y�OG)����_c'sKQں���ѥj&��-ϘQ�^��ɌB�/�<bqz�������55Ru u �L�P�eUx\��b3QJFfg=6w#��z���u*[&Tv��^ñO~ǵ�'���p�o|�l�w�xjv��{h`i���0�p���4��
e�)g��d(��^��Y9��EV4f7��m��w����z-�XH���x����+&n�Pk6���;?��D�J%X�R�s�cL�cyj�T,D"��r9��T�f�a֋;M:�P�gNE�.���=ʹ��g��}�ۼo���x�\IK*-�F�tip���ܺ6B:���˫�z����hz�_~��N.�GW)+�D��G>����s��(gq�jԲ��ҩ�{ow3f��l6���ZW-+�K\�r��F��$s� �-�8��J������"-��l�{4�G���Ƿ�}U�Z�����|��Ek��@ ��S�v�<���J�t:�,�m
�KGG{M��4z�d�q���YZ	�$���D��,k6n���GG� ��Hg�L>��f��>��/�f�F:\��x�G?����	|�ɽ۷9~�3�./=5L!������ӫTD��U����ʹ��d�3�Y\Xe~!ģ�"�e�����x�M������*X/��1�&�a]/7������7l�`R��{���z�q͔1*s� ۫X�d4΃�ܹq��n����d�T�#�~�q���+Bd��B�b�������\�����J����lf-��9�>L$�$o2���}�y���<)�/��R�X��.3sܾq��[W�NP����ʂ��)�I�W��fCow)5~��6^|�<u^b��z�E��@U�����K��"!�H�Cx���{`���FŪ�Ӫ�VV<���1�`�|2�.��#�������P%EJ��թ��}k��?4HS[�U�b�V_u��u.������lߵ�k7α�h���rQ�E���g�~�_�,�f*�R�lH�<r��?q��Q(������ٹy�Z<�#�<�7���}�v'V������H�P8.9�
5�Zb�llW�¡�*�%іz�����C.;�l��ɲ45��[�048�h�^�m��ؽ;|��ߐ�1��]6��u�M�^���������29������r��8+�4�gc'�C���DW��4-,�/����*��d`������؜BL���9�2r�������)�6k���J�a���Z���3�S
�۷�|�c�V3$�b�ubq��ؾ��5��XCC[e}��D��%|un��p��I�u$j� �d�۵{;w�Q���tٵ�8�F\�4�ș����)8Ц�=��ױa��èt�h�筻�\�y����Ĳ%�b�38�tS��C�ņ���MÛ��D�~����d((:��-���[��",w�r���F*�4gN|�ȉ�ԙ�4h�jo����ؿsY2�8+�L�N���diDf��o��Ў�ӌ����������`�w[��6��W�g1Z,8��?�4���+���0ϕ�\�v�hd�I>{�1c�%�N�U��+���έ*G_:����n�[��*(Y]}�45�)���c!e����W���w�Ϸ@�\��̢8���ݹ�};�p�M�M��D1OI(�TT����sܾ:B"�\�D��hE�ҧ����K�Z�3Z��g#F�O)��`vtw2�����zuoJ�-������\UG���a�����Ժ�*��v�����Ӝ;�5ӏ'TF_?����\��-s�R��(��T�>�BQ�۰��Է����GK{;6�M�=�Vܞ�W?���;���Z��[�u�C/?�j�dP�Zj��Ǿ�ƕK�N[_硵��UO$����+��de���h�hM.�&�z�.&�:�����~z��in�+񭐖\� 4�h�F"AB�L�te*b��e5�[k����W*&�"n�"$�LЪ�I�v9D�%Ǥ��N��Φv�}M���E�a5Wxp��ņ(������,<~Dle�l2���C�� �R�|.V-����צ��f���J}K+�l����,&�e-�D�ތQo���ܹx���8�L��ͮCo���W�d�DB�4�-�I�$��&	���6k�Xx�R6J%�"�5�J}B��H��qֵ20���7�������\�ݭ�_��S�?�K�w��N�=�q����;<D�)�ǖa��1(orB�����Dsd����a��8��\$2U�W�%�UX�_����]l޽��x�HT��j��Z����z�0��ų-.(<��]�x���(���b��U��EB�Y!��ˤ	u�H�HE�V片�I���Q��U�'�vZg���x��z�n�Cs����XJ��jy%�߼y�s'����,������_`�d�6"��[�������KE"+ˌ߹��������T�IʻkT��|6�����u�~�|m��u�Ǳ�-V�ʅ�`"����O��u��d<+�ۻx�{?���B�2��jPԶ��9�W&	/>$��M>���$�$�����+P$EW�S���KC��v24����J4��J),*f����q�8{�<�&��φɦ#ttw�i�a0A��aje�h6���AoV�	�nʰ]�aq�.�������hrhK\'�z_5w'�Q*�����d��[Գ	��M[�z��o�0��Ym��q�ӏ�u�,��
H��������^JZ#N�Wx�%�w����\|D)CW�aԀEj@4it����P��r���+bU7X\x�Z�]����Ocoh" �r�'ұ����
����ٸ�)~�=
f�N���f��)�^8�ĝ���,P�>&i����րݬ%��0���j$FV� B�����\^��������w�%Z�h�B:+�J3�\
���鯾���$�^��x��Y�W�����T�d�R>>��J>ɕ��p��7d�A::hnp)5���ŷ_���)n\�����\n߾����eq9���|��l��`��� ��8����ز����g��F槦����5+�ԙRћi\���_~�-[7�v�9}��ΝU��B2FG[#f�,��u�w�6���٬2 ?����cG�P�!������REv�9@8����}Cq�|������w�>������N+��d�{֭���^WЗ�Z7�S��ӧ���%j�:^{n/^����A~���LN?�`6������[�渒�)�O ������w�#Y�P��f�S����1��)�B�me;]\�f����7�q��)8��b#���CϼLww���҉V���D��8�,g����e�z,TJ)jj�'���$���lm�D$��A%�o��1b�yؼu6嶺o�ɡH��.;Ν������@'y��|�W�|�r��D"Cc��V�ՋW�y�[�ϒ�.Q�)n���tw��8=G,����A�>�@�`uh,.������KSg�A�@�    IDAT}��u�a;��bՉ2�3n�=S��	�Po�{?�{��E W�C��J4��'�~��*�K�X�&�[���%�-<Q��fRZ͕kD,\��6:z��b��m���$�*�M�Ek��y���o�|�*�<�׮_`z|����M2Y���g@+%ϲ�Τ����'B�\>ɭ��(��1VRض�w�x�ΖFb�U�O���O�:<̋o|�cGO�ͩ�L�-��h	F�$�Țq6����ǚ[ټu'���:��O8}�KR�0ش8:�x������Q����������Ë�y��;8�{�o��U*�l�G.]��w��J�eF����diI�2Z-�Vo]�ؼm͝j8����dJ�S2�eöm������s:��������gnv�ޞF=��=[���X�C΄\�����C���+ys���+���S<��ee5J<�Cg������:������撥a�m���Y�����*#+
�"�j4l۵���v�]�rE䋪����s��	N|�G�(�-~����l��e��1�`T}��P��H�����[�鋯�uw�`(IJ�wg#-��m�l���k�p��9�����Zc��mk�o�M�@�d�F���f7���|��g��e��;ٽc�}m��n�C7U6�Vֿ�_�����U.#L/��(Up5u�ع���I[��:z����y,L>����?�R�8��γ/������(Dg����ų�>~�d,��m��D��C�٠U��B"���}�������D2e��X�����νnںZ�l󐌧I&�vE|6>��aF��S�d�H_m0�=%Ykбk�d>�Qk3�U�{�/��hbnn��gOrk���<v}���Zz:����RK��&>���������&��&��:��1��8�^z׮ap�Z��ZL�T�e����֥+��{kY�i�W_�ӄ�T�9�||��o�s��BkG3͍~,f�S6�{zj�PpUAmr"z�
Ȋ��PYT�Ë�����!Z;�U��n11�]G`>�O��O��y��Q������a�y�i�.L:�������g�]d���t�6��Ҥ,��Z�x�"wG���H$*� �
Z���	�Ů��	o��u�ؼy�Z�����l0�3���E	�2�(�b��\�E[�PJS�����p�l2+,��&EN�aPqCJU��&��Ȧ2*Z��{�hh�i�U�`$C� ��j=�A�!��fej����x��\V�Q�I�/ĩ��$��x��aDgw�a��o�{p=w�S�7���/߽q�����:}�������;�y�tQOZ�5�F�+��h���<��"��q��)*���$V�	��Sc��y,t!M�`�6b48h���7���c5�'���;�y��c�����1e���o��ӯ����!��N*8	��,��duf�LlJ	*�e*���%�J��@��sdk*�Ӿ���&[wo���!�H������$�X���EΝ>��ܬ�>�a���ɠ%���q�XS�2��X,M0R��xp�tx�Xh����TD�ich*2����ƌ�����;X�����]���2�<v���đO��NC*'�;_~�퇞#%�#������J�ũ9�+A��&L�#�	RS�Qɭb3UpZl�FW��p$��?�k��Z{�ߴ���Է�(�I�P�ew�X\��O~���)��J	� ���{Si15�U�Wxq���G�.>fuy���cJ�4B2�H7���B�Դa��JK����F<��l��4�즠1U�uBM,k-�e�q���Fo�N�eB�Rae=p�w2H�~�.��F�9���xŵ�KDY��`y�.������rɳW������VEĕ��&$��f,�L�,159���RJ0X<tm�Φ=/��4�3Z��詣�ƙ�d#��M��Ǜ?�M]�Tj�u����`��m�f�K,����2pKO��㸝�k}j����H:�g5�!*� ����������toڎ�֫�]�x�c��+�)&
�~�~��.y���^�O�oc��u&�]"�0I>�h,���I'�q�5��k����T�K��&3*z��<�X�vr%3Ŋ���!��&M��h�k5�f&K��¹c_���ub�e���|���������;��:�ڛj�l�#�叇�g��\u�6�S絡�dx����������d��6��nӶ�j����#���G8~�"�q�j?���g=�6����^!�J������CYr][�����Y�f ������_}AzeAm�ۚT]DK[��a��חɥc4�}�ǿ�?�%n��B�Ⱥ�a�	�~�>w���M�(i�l��û_``�F�Mr�������j��FKK� ��.�7l����;N���m��q�$��d��JbK�������C[��,�,(ݸb����o�g�>�_���D\��y���fx���Y��	�|ii���&n�<˵�'�RG��P���̡g_���GA�dq)?���8,�Ψ��û7����1��\��^6ٜ��{TP'аX��c�d$�l5K"D9G��zٰy��R�Cqۈ��̩���#�q����v�ŗy����]Qʊk4�<���23~�|l�z��Q�V۷m�f5���U����[	���Z��R(�1�j����t�5������Ԋ岤������\;}JY�&$��w��=����b0@ck��Q����������ُ�T���q�ˋجflfku�,��\Ye��Bi�̽�����Un���u�{����5:WȐ%�x���??ʝ{�|������q8�Xm>�I�>��@�R"5�ݯ���[�;s�xp���Z��vԱk�=}]�QΝ:�/~�SZ�������!�f9z��O�c|r�J��l^GE����C{��}���Ne�����|s��lLe��Z�z���u��TWO&���~�����5�Ծ���=LO{3��]�z/WG���>c��u������Ư��5�?EC};Q��"E�Zަv6m߯����(���}ܾ���46C7����P��R)f����s��Iv�\�{�Ě5�x]�)a�w)O|u�G?�ޝ[��^�b\���1�M�33�@*YFcn�ݲ��M{�[�Yّ��(�>q�V"|��Wʍ��K�AϦm�پk{�$v�R��:+s��G�O��s�Z^>��=ۇ0ՔqX�Lܽǧ}Hl5��l�=}<}�ytV�����k�f,����:l]���J��@ms;�n��m��?��'����݉���W��6��-j���g��~��_�ɦy��C�߷�֖:���mIՎ�f��v)B�7Ǿ���ڛ[4ɹ��ܝ�"���ܵw� F{;u-]����L2�o�����	�����o�ź�C�
)�Z�_F�s�ɱ;T�i5о�櫬h�hHK��^�Si_
/.XZ�ܥ�|s�k��Hh�Y�h��I��0�w��]��*:j`%���@W2��������&N2s��z��Zp��QM�-�ױk�f�v��p��Ȩ���_8�%�|��7]���[����%�����{o�ß���<Ɍt��h�V��ftvޖ�l����z�IEz>���p��%Epu����<ġ�����M�����}>��,<����;7���BkK}5�YSå�#\87��RP�ɬ���a���`Cg��ч�Vl�[�ܠav���F�D�����fJ�*��u�o�Į�{���nԐK�p�����֯馻��G��IĒD�~��015��B�H4E('�H?���2yF��ݍ�l����m;���׮��\*�xkz���T���#�gYzإ'�2f����4�����a�F�Y�s+(��aPA5�=���Z��i���ɉݮ'/�MY�4�� +3S�W��.��� �	�#��(�ٸ�Zq��* �Nd���
�`&�h�5bv�Y�a;[w?��d'����wn1v���Q�B�y�?c��H��dE�e2gqu�Hh�������Iʅf��%��T��a*q{k	FCʂ���O���Օ(�p�}Ͼ�΃/P28UV����:��W����=JɄ�*n�Ł������
a�L&�VP��.�M+�^fi�r9��\�D_��R1��"��bIe��"yQ�#���J!�	�j��q
&�WK`��9{���YU��}�N�}�yI�\��Z��ɫQC����p�Dh�����I��@�.���|���{ҝ%��4%=��Нt��E��&z��+����v�����	��4BO��9��;l~� a	:WL�"�ss,MN^�#45N1<Z�6������zO��Wʐ���C��aU�)�M��P۶�-{�}�̵>��I\�Z2�0�?��\$�(��W��?�1��RbK@Ol%���8+S��� �5)t�2v�Emk�&#�Z���*K��Y���З���M}�z�z��-�d
eVVě.ɤ6�F�p��e2�U�0�T���.u�,�o?���@./E������2�<�؝+�=�Aj�!�J��z;ݝM�ݹ���ģ	�L����{������#Y	E�w�.#�.36���j�R^��m[�����8�~��?�'F/_ 	
J���7��t���$]����������I�e���i�����S%�>����v�����۹���$�19��j8�bP��E*��[ٴ�y:7cw9)%�|���:B!%������[�R���*+w��w�w�4�Sc5 k���z����� ]�u�12�8�L�F�4�l<|<ǽ�SB9b	9�l~�y���6��zVBR�lB[�Pk5q��&��$]����k<�_dy5��ϿM1S!�����nRC���Nti��[�E_S`ۖ5���n�N�������ѢT����S�؂��V�@(��B
���5V�Z�������?e-�������ue��=�������5)����	����p�i�����m��7��R�X�ش��x��cD���v���x��x��w9~�"�}~�����*�uo�:��z�C�^gjj����\x���ZCSG?��ٴe�:���o��y����޺�չ	�������~��#�XY�ON�LeI%�$�5O+*��Fx�)�տ��\�v������L/�����������e���@T�������zn�8ˍ�3h�v/tD�����^�U@`��Z`�3ie��ԉc_r��W
���ӤT�����u}XM5t����⮨���Fn�|��f!����eŵ�!��A���`��0X��g����|��$�!&��*�^�^{��U��0=��o�:½��i�sb��0is4x�x�&5�{=�����p�6�h����I~⪗����BS[Oc� �;�a���6�tp􏇹x��H\)��v��Ȗ]ìD�ʉ��8�����dt��k{h��T�luu��'O(�e{[;.�C�@�ܷ*[j0TV�J���`Gct��a��W�4�S)��"�\X�S<�:N|s��W����p��y�n^�`vbw�Ig|�Ezz�U���M⭵+���3G�w��>3o���ݛ�s�r��l��{w�v��tu�04�����p�50�h��>9¥+w	�&��B֠.��{��S_o�׿����Q�{y}��?���m����ʇS_Ņ3�0�|�[/���aj����z���Ց�g����o�U.�Y�@2���lX�����_~��[�X	g�f�ic�w�0����������[ׯ*���na������]n&>��_��l6���z�C��Fo(����-� ]�����̍��%Ƒ-�����HGOG�~����[\b��,��W�:Z���5����6��|`"��_���#G��Iƕҙ��0Z-��2�vQb�Ib7�h������8������������>O�ω�c����|��qZ���30��<Ӿ0��1���I����^ol�����x������^ˎe[��)���
���2����r������}�s���.�d@��N��y?���`fr�SG�s�n+w��;6O8ل��MV�e�_�Hq�����������tWZA)�{W��Ì6���?~���4�V���Tƌ[��2<6(ݯYY�d��S^Z$�(�mm8�Vt�jZ���?���v�����&�tFg9fG6eu%�Ԧ.�o��}��uJ��55����K�X�/����	�'%TѠQ�e�&�H��HJ��z�u*��Y�G���I �N]���_��op�GAJNy���:�P���ׯ =�����j>��s<l��}�SPuә[X� C�p��ի�ٶ�QV��A/jU�tvN�Oq��	��#4Tд��U�2=v��U�ݹ-7���t�<�;z���My$�	�]J:[���vJ��Y����\Qo�����ޒ3��i�����;).I��v�>�H�'6�_Ɂ=�q8�tw�233))�~��3$�N����y��쑀A�Lֻ@�ʲ҆+�R^��[�uY�-��٫?c���$���FI]�װ�&�}�\���q�2�4��v��_����(A��ɞ}����������015+)��)ΐ
����7ډ+��e粪��u5ح�#���,��ӡ Q!��j䅞X<	��:��)��u���7
q��J1�pjIy���H�BWV��09Q,��h5,��R�,�'~����A9��fqD�Hu�V�b��uTה�v�Y��_�II���_|~���>L�Y�[B'�w�~�6�a����=��0;�N<�G�ѳ��+T�݂/"0�	��(�y&�Fqύ�0�Cpn�Dh^Ԟ0�9,�&i�T[
k�������O?f��eŪz� I%o�'�|���8y�k	.�����i.����[D=2�[U��M{���N����S##�15�Chi����2�z
�\��Y_�v��� ��x�>ftw��H��+��i+��o�`s1��H ��X8!�W�^�;2"��k6o��`B��Bb�-���K��3s,LN�������}���R�`7�3�d�ҐaT%�i��q@�<�����V��kY�a+%�U�ܬP&����N���?$���x����)oXǼ�@�jI�ev|��8ީQ"�C$�K$+�,G�r]SW!c<��*��25:!���3}$IÌ?���b�c���}Q�@�m4,��+�	�dIٞ_�c/���If�L�1�������D��IV�h�82,de�a1��(/���Rtj�$����3��2�ॳw��I7q����z>�g&3��V4��b����۷����<�b�g3>�c]����%MKM'��/��;W�i#92O^���Tvnۈ�禷����:�����`Ue���'k4h�F�stuvHx���񄞸�Nzq=�w��~=��2��&}���/��������PTZ#��33���T�5�&�P��HIՒ�a%7#���*Vծ`E]5�T�t^<�%��|�(Uf�E�XO{�=�Cɨ\Ŕ����-�)(.!�8�'o���[7%2]l,j�7���  Y1XS�������޺"�9��)�X4��J�rlnZ��3G�{�Is�14x�|2r-�5��X������k��&�畳��ȫ\�좠h>���&.�8F[�u�k��Yy����L02�e��C,G�#��Y.+W������4m\C^v*ᐛ�[�Ѱ��Y���9n\"9�a�ʍ��(����OBY9��V�P���cb6D��4*�����?����_��_���P��K��V���A\N�.����o��DYU]L, �>qqb�(�ELc4Ȟ���]��F�$5�.�8ݽ�\����1:�������сǷ$��˚*Wm����#���~�GL��W�+An^!������Ź����_QVSL��jr3�dZ�h���M�$t���C�Ϲ		h���)4���K������_|���:9^��C+�E�8�ҷP�2��Hǘ�k�t��a����߻&]x"��R�Ш�4��OfF@�3u��V���ʗG?a~z�UGiAUe��ز��o^F�]D��ō�������W\���$#S��CQ�s\X�6��^��u[vI5�Vk梈��=Oл$}]S�#�ܻ�����=�?{�k�Π�)�O�0�5�o��������#77���|��;�1�\�MF�ܿ��~    IDAT��شL'*�SP��S[ 8@ǿ���M;��͑ɇ�z���ɞ����&�z�Y6��/ /� ���֙/��Ie׶����`2������x�|�VV��qz����i&&'���axxXbէG�0Z�,)(4��VQ�jk�b���N���(��Νn�~y�ںj�:�i�-��Fs1�lߵO����E"�%23�͏q���D�s�_U��=M�*�'E7.����Ar"B�A'���~)���cd��y�NJ*�h����\�p���ey�P�и���?M]]:�s�/?;.;S��J��g�}���*yH{��_�wO��i%_}i�a���G��]��N_w?'O����
��	f槸p�"�������8����?y��	7s�0�� ��2�?�<�n!W��o�����.b�Y�����Ïˈ�H6ܿ#��e�3,,D���܋ORXT I���߽��M��,���>��_�:�?�4�~��O��������*k��
J��Ҵm��&�=n�ߚ����Q�u�� X Q�F��X�a�}	vjJ�������g��&,�50=DUi6[�V���v��<畗���������g^a��x�g�p�G�8͝�>��$;r1�W�YVǚ5k��*��G8��o兮V K
+�0h�0ST젧���_�u���ڴ��W8��q���UVW=rFb���R.���5��n�2<0�ÎN�<��{	ĬleTn��Ȣ�����JP&"����/��tʞ�-=�g^z��:}Mr��������uw����"5#U�b��L�eHb���FO^aᄂ���s��m�{g�/[H+�#����VOYE%kV�����EhF>��(���!�`MuaOKǽ���/4lB��q;�5�U	ƈ�֫0��\�x���>�%�5�_]FuE6������U<h��eQ�J���~Dv=�&��Z�=+�p*z'*k:If�F��E�[���b��I�������[�.�V�����x3e����er�,ع�t����ӟ���t��LN��y��)+��������޿��� ���F�M�kC��CV^9���P����B����U��A�%%�INY[�oduu>����d���;4�LZ��x��7�|2�2=3�O=��M[�y�>�N_��w���y<�>��'i�;�P��$T�����z
���v���ի���KϨ�I	+rTF��k�����
)c��0�����&Ha�>)zf��2��$VU�¬���#	���Go�bnb�����a|�c(�~̆$��乨�)a�Ƶ������b�uJ<��{��\�p���L�,
�
�x��g�LN��q�]w/3��N\�w&���
�u��F�$�TP�f&�bqn��L(�EMF��Qd��������O�]���?�`4�_P 3삚v�A��"�|5��YT���djt��}D��m��/`M�f6����`l�ٹif'F�b�����a��C�P^����6l&-���6�6�[P��!y��x�?����fb�MFI%M͏�H�b�AI9��ىi��;�wX�ŗ�����ݻ���'$������0;=�o~��g��n�{���Ѩ�Ѧ�:�X�36���-133- �w&�Ⱦ���q��C�X��Ʀ��ff�a�n�mn^��|�1���J�c/~���RW�������b+93Dhj��NF�d�l9"�+T�R��!�(��"���Q#���39�kl��i��<��o�SY��䌄>���Z.]&,:.3i��|�)�i�$���g<��3���T?~��5/au�IM7����dTI��� f������Ε�ۉ�))т�n��Kn�ͶL�o�K���DF�<b����t��>�n\�/�X�#�(��%h���zٴ�Y:n"� V��tW����޽E׃D}�d95Ԕg�nm{wo��_��/O#��Ph�^A��@"QFF�=��cH��kY
j�EM������c1���/^��`\l&E������_�`�)�k�����L��à��LY�lZ�nՐ��`͊z֯�(=N�%�ĕ�?s��-7HKOE�2�ƨ����{����0:�DDa#%��Ɲ�غs;�����-�woKՂ�V�]϶CO�6Y�ܼv�����4ԉ�n��,��(�1Օ�<�o?��f�����L�;�s���xY�I��g����Ԭ���~���=�S(LN*7�d��CcZ���[��]>�%7���1xk��}O�gx��)/���0�hQ>z���߻FAA7ԓ���*9JA����X
����pO+y��X�Z�v;Q�DN�eI^f�&ŕIQE-#S^�Lp��=�b��w�G^N	��ӿ��q���h��o�	��k?��݋<�{kW�-0>������0��H�[4cfz�����<��$��:�#��ݏ��YDo�0�o�blrRn��q9e|�;�^k����{�H�U$���o��k���/tw�eמM��-@��};Q������XtAv6��������I��P�8��d��ȋ������������O>��4�����:���M��%��,J	��b����M������'�Ȣg�R��hSؽ� �i���>�9�i�D}���i�~�����|y(�׼�W������QZ\,��b���2��%}�e����ko�����E"�o���bU�Vv�{���<~�3�O�0��x��غs����wnp��G�<3rc"������ߵ�¼4.�;ΉGe5�j5K\���-�2�(+�����ܾy�w��`T�P��w�U��u�v��~���������{��F���,.�ٳ/��o!�gbz�w�y��������s�z�� *U�����7 �z�F^�f�Ҥ�Bt�=)4����^�&���<jk�իi����l܁9���o����'X�P��H7�I�1Y�dZeg������<�ŕj���wn���4[�W�撕b �aar����.b7�$	1�������+��iY9����+9r�7�t��d�\0v|�����=�/>9΂g�ŅyL�i<��K�Y]N���|�ޛ�[xQl㶬�ڹc�����(��/���g�Q�Q���C�����8>���?�?or�~7���ԩ��y�Y�<�%%�_��m.�<O`qQ�ª�*x��r�R����(�,��i�l�{���R&Tq��b��*�ѣ�Sܹ�����^�����wJ�yGw?�ó�0av���f��?��lfVl��)��{8z�|V' u��3�z� Ȭ'$"�A/Y">83Ɖ�QW�OuI>�=�$G�xl��>��8MR���t��i������oqQ-�=EnN!n����q�FzG	%���U�V����kص�������^���u�Ǟ}��T��u\?s���v�ˋ�(Ƞ���#]�{f$�L6��uvrZA��J�ڕ�T���4���ŋ��p����>%I��J�v0���R����p������x /�\Y��ܷ��l�����&XSS@a��r B:����J0@g�3�^`bz�4���U�%\�"���]����9v�2�3A4�\��PY\8�2i޵�Bˢ[$����8��ݔ����4l���(���.`+��ٴq5j!�^M'����]��NB��1�M����s10���G>�d2����obKqR�z�3K\�v�����g�xD�CF'JG
���d� :�Mk0(u��ǿ����t:�vU�<��~��l�w�p�����UYXLj�޽��~�o-&�Zs�32ƾze��!I���6.\<OO_�C���$�.����)d�QW���j��׏�y���.(�c��uԕ�43�n�,�IF�S�)�޿�g��/���d::>Faq	[������Ν����7a~�+̩�mYh-�(v��ҳrY�f�L���� b�>�X�ϸ�KH�y�P)�B��@]®��5�vbY��Q���.1
j����M�����ukѫ��O<&tz�FG���i��]��77܅"�7�NkVW���@�K�rS�	E� ��|s��U9hd痡6�_d)�`���T׭#�0�ҵ���;�x>�`d��_#�r5���pON19"$��FH���̲RZ�Cn��U�Q��ը�8A��z�}44�!5MD�f����^k'CCsD��7�a�ƽU1?%��0�����	Iԭ�¶��X�,�0>��̀�ׅZ�`R��i�=M����Y'��*�F������-���������'��%�5S�e��dQ� ј�pO�p��Y<Cr���i[w�$�T%z�;S����aY ��3�<��ovURG���,'�y�f��bґnTaT,���A{�ٹ�j�A�I�:ǘ�`r�a�nV5����wos��I��ƈ��$i�z��0��ճ������P�}�&:��GŅ
v��V��jay9$1Ǣ�%�ɂ��R��φ����?<���<�Z:��`c�Av?�4!�N��ɓܻx�В��Fj~���$�1��~}�;<�"�%Ŧ"-�La�K����Ifzr����9dd��p�9 ��X\p�������Pj��r�Y�m/��*feG.FFF:-�[�y�~���"�/9��$��L�/��� z��hXD�\��l���r��y��b3�ڕ��;5�_[��m�8��Q>9�	�%��l&���j�`�Dr�$����d:l�g�3=�Ă'��� �J�{���r��=:��&��&�+��_xYjf�fyp�6�/�%������B+����GF����K������� ��z�� �X��{��_��˴���{�h��[��+_���߽�[Z�ߓ�������v�?��ha��Cf筋�#n*
R�_QBz��"B��@c}5?������BIQ:j��Ř��Gg� 񸚂|��ɢ�c�KWZ���(]�_�#:�D�PVnV*�O��ƹ�n�6���{h����<)aA�+\[SN<���?�!����U��IuEV�S/��`�������t;ׯƳ0�hSg2197GvV>eUܽ�*#�?'�p���'G/10��}�o��.�����Vr��(�<|9��m[�����_25�ɟ|�yV�e�M���K���|~�|ѧ��%�-++��d� ���k����	�a�V�j�4�7Eo��щ9��$�9�|�O����"����ӣ��G��������h:�����7�֭khl�$����Y㏿�g(�S�̘�ɤXL�+�o>o���3��γi[3�7���`�{�����$SS>Li%xᛤ�2>�A��K�CGW6��{�.2��.�Ѹ \�jm��{���,��>�e��,�N�ޛ�bv���\��iZW�ݢ���+�Ξ�e�R��'�m��%<s��J♓�IIy9:;9u���?N"�ĲBOY�Z^��ש^Q�G����1��S�}�.=�O�[�{�m�޾Bq���QS�CA��L��vY�v�<|�.f��];6�Dy�O0X4��K����V&'0e��Y�	H�H6�vSU�Ħ�����k��᭻���G�x�"�>�,��7������9�����Z�EKIau�%v�=��B8Fw� ��9,��1���ZB-�U���'�����Mhr",+,�-��ձa�N
*K	'D�aJ��9u�
ǿ8!eܽ}�<�zIhfk$[ٱ{?yyy���zf��K�dx��v��� �5d�LԖ�03�?��w�*�r�*BA��=X���8J�2���/��}��g�36$�0b�*f��<��ܻ3�g}!7���%2�
x��g�[Qć|ȍkhj��'wS_�˻��)=n��b��qKr�Ւ"��"i3:1J��k���k��_ƺu;X�z#?����,��,�zX�[X����COPVY�[���cg�Ŕƨ�����:HEA&��ɤZ�ҧ�H����cLy��/JH]Y^&.��p(����p8���d��uT���_𰵍��>:��FT��T�l����lvf��1Y,�݋=z�E�<K^�\PX�q;k��(^"�ecd���׾��$��
���9����p��eFƺ(-ϔ�dMrLv�UbI���1��,7���뷹y�!���N&)����լ��{����?�%s3n�T��0����Ԧ3;;J������W�X��kg��}�?�'	EP(��_���,�$<e7Y�1(5h���!7�10�!I���^�)����R��h�(?����*w.���#��{v�sW��ܸr���oa���1Fz:���dfa�����gt|��T��y+����#�hjj��f�?>�k?����
�[�喑�6�k�V2R���S�8~�4�._'at���tɄ�wI0�3���׮�)�R�9��z�{�:y.��C�W��䝥��|��W�2??��/� 3=�W^�:&��/�]������M342��#�2��̔���(+�䱽�d8l��'���KWQ��&�+��Z"�ae���ّr]vmZMn���W.�����k�,-��x���������j9�tvwJ�����Yaa��e�u撤s�ԦP^V���M8�6^���~�.�j��jV���yyiZo^$ꝡ�����y�?y��V�*T�$If���8m��DNN	7o��ĉӴw�07�D8�@mN���CepW��Ө_����U�,:��HR'˘���8;k�o\l�p꘏A	����f0F�h<,o��f0�,[�"&*��#)n8����oDW\�$p؝X-F���~Hhi�� KS����*�XU[DUy���ݺ*�č�8@��E�9�h)&Ҳ�	�t<����>l�|�+dfUr��n_:��h�����}���:y��,.1=4��`��(ǖ���1PS�#S�r�.�L�Ml��Q`͇(.*������t�G�e��Y��V������]���,P�y������{��H��-�x�)�V�twu0���TWa�$�e9�	r2���w~�{�/>~WF���V}�����3[�[�r���p��������蝹4l?�����H2�p�
5�3�����8+7l`���ą�YΓ��I�{���?;�{�����(�u~�&� ��5u�������"��  ���B�H#Ih�N��<�w�!��Ս��ڼ���J��o��}���I��+�y��ڕ$�O���q_�f�':�N��\���i�l�JPMv�#JOw�t�:���!��s�ܸ���Bbc�s���#'�ɇƞg�BaU�T��;s��Wnt/�4�fg��C�f��]�3��O_k3C�D���*��IO�PU�-��G�~@0�j�'��@�7I̲�dbaz���It�d\F���Hmc*��x��j�����f��r�+�ʨG\�m��d�d�3�	�|�0A?����$�n�ƅk\:}���>����).g���W��P�������63�H���~fg�$	P�Z�Z23\h`T%SUR�䨇��Yn�N�ҳc�a��?��q�^�$)��:�;=����1:8��˗h�|���{(�7���]���)Ξ�@Wg���{����H��!!L���$��M�Л,\�u�s���;�Ȣ/A��-|��Uo杷����[�H������<,c�>�ԱO��i�����6m�#=���¤� �p�����wn_�NEy��MF��Y\
�Pꙟ�166'}}+Wl�r�S�n�d���#z[�T��yVz*Wϟ����):��m�gh���0�?I8a~v�ҒI�{�?bf����ڳ���\	j�̌��1��JW�WVQWSʢgV�i�⿧P��ef
�{��(O��5�f���in� ����OW���_L�����!�4��ǟx�UϿ��?��������J�&��, 	��!'Ϟ��H�0� �т)(�ABlu��?8Do�0Vs�E��bh|lR�Z�L$����o�������296)�&ƒ[��7�����U�����@l��M�X���9��T=ݭ7%�h�=�~���b֬�f��0;����A��JN]x�/��+_�����y��/8u�6Cݣč�����_��������촵��fU��z���y�	������={�˞��//��s2���>�f=��)bUu+��RL    IDATKy��?���S4�r�S���c�'�Ө�kiX�L��CA��8�`�Q��D����+_�i�z�����|�gރJ�F�S���~�xvۻ���@�cۖ5e9)̶S�� +ӎA�����4��bm}��	r82ټe�,�3>�;hk�wHB
��@��YT��}��m�F�����s���f�gQ<����Cv�Y���N�x�7��<��.�j
p���������	`�p�ɋ�e>�t�!��$)�ʘ �%��9BG�0~_I�T\y�l�Jݺ�(��Hjia6'�_���c��1��:i�z���2XV�پsy��C>�z%F��������PǗ�EClm\Eq�����cd�����, �-XI(T��䒬�3�ࣰ��`D�ǟ��~��d#JS*w�?�*����{���������<�x�qJJsy��_34����j�@�Eɛ�������fS�����'C���Q+����Y�`�ڰ�3��dp��+ܹ��/~�&m�L�{�)��Ԭd��Cl޾���;Ι#���@�5�|�/��Li��QA<����ns�ėQ̩.I[�,ʑ����V)�	zv����)	�;��s�vr�������֍ן@kȢ�b��o��2d�l�����G>g~v��C,*@pF655��n��0��d8�xg��G�K#����_�3�
U��'�T��"K�h��m&�r�Z�����vi���B���c������T�WR��~��:G������,G:9E|�0UNN����$9v#+�r��X��X����O��_R�Zk���X,��̄T;�)r�-"���m���8}�4G��bhċۯ}��\��lݵ�u%���p��eT:%uI�ľ���r������������~Zo_gh�G��3s�IqY	D�,�gP+�fc���s���W���s_��~3�.��g?���ncl)��r-+��U�m\Gei���TFΞ<���%�Sowb��%'Dt~������U�_�
�A8��ĢK���xF: 0��@zu��4C#}��!֬]EZ����T=hUZVU7PTPM��An�z����=����	Ǖ$�i2re��)�:Q]�˯_{��.�2P�d���3��i71�~�遇���e����N�������%]��x��0*D�,�/ȟC#�F���������I��!kn
S:��H�d��.�
r���^���-�
=�TUu���T17�O|�I��(Gn��Ǆ�>Aff��(~��$E\Ƨ�����8S�G+b���Y�I|b�h�	gnZKQ���Ί�z6ml�`���#��s�8S?!���(�s\��d�x Kr���b�h�&��o�����|<��ߘ�g	WJ�7m'�37��rL�-Ł0uw�J]��d?2�\U�CSC5[��X���O�a��SƟ�\6����-)Lv��@(N<�Ln�j�U.~��Q�f�<��?�����>��[O��`9������R�zc�^&'&Xf����6�2k��S^��;3������]R�(\0��Ө�jr�s0�,$)UTϓ/�L�n��\����&]}n�k����K�&9��'0?%A(������gQ�t�����ɡ�{�q���д�Xle���מ!/��;�yM�i�
�Q�Ut18>�R8������5�5V�L��Qƽ�Xs*X��iY�v{#2�(z�'O>I�rc�l���e��ɀ/ehx@�H�hc��&m�ڲ\�"~FF�eW03?�A��=D�g�Ό��p�جV��aseˍmK�0��XrJ���3lܲ����������#5�T';��~aԴw���݊wa���V�s��X����Jl8S30�X� ��K������������fR[^�ÙFB���p�^-m��h��W�F"����Kܺr��������9������5NoG/�=�w��<OqE�U�2fX��NQ���x�Uzz[���J�P�tX�N<K^I]�̙���rJ�4��H�rwЃ9���UY�)�"���󠥕�g���ˢ'��O��.�{?-;~�S��O�KǙcg9�����cR�w�ZLz!%.������V�����@ dfn��N�RI$���F,��??G�p���\��ƙKm�V�|��u[8u�$WO#����1:Ry��(/�������N�y�/�p���HBt��)+�c~z��><B[[���'��KV����Q�%��	˾疭;X����>N\����IFf�r��կ���,~��7�}�a!TU(�Z���?������+�8�!��N�3�lh�d��U(�"��Q��$�8��S��OSWSL�݀�d -+�щ._�-�͑��EO���m$+���s��-|���SZ1�nAM&3���s_JcH�$Fv�G���w�1KA������W��/�d�}J�ٶ�^&��:8�(�����<J2(�K������4|Cc2����O{k7�0�h>Ȟǟ�������5�fB(��|�����
~��34����F����V�����Y������A=��]�Vа� �YIoo;���:��]ԮXAVf6�@����N'n��w���)Z[;�����J�8��Q���1b��������*~��7�$z��-����e��˼��`)����;)/N%'�D�U���$E}8LZ��ٰ����+Q
%�/H�7o<�[�Y��Xٰ���̥�p��=c,\|��-�����	�àӡ��󎌌>8'�H��m��ff�������TN��kOQ^����u��N5��?�ލ��;�;R���%�I�ˌ�3<6,��P��������?AWߘt�--E�8�y�ٗ��q�^���~�1����39ph?�?�InB?|�W��W�o�6�f%����a�Q]Y��� �|�=}�lnZGR܋�'�@AR�r�錘�6\)�,·����6�'&	%�H$�hҊز�0;�o}���I1
*qX���o����c�N��G�jM5{w7��y�(�"Y�?�G���U�0/Hx	A�\fzj��N}C=�.���,�O�j�r��{����y��F�øq�;�Ƭbjz���\n\�ɉ�'ٻw'C�ܿvY�M��IF���K~A��oŉc��q����7�1�߆1)��^x����{�7��(�Kg��E,��d"��3;�&cu��_����O��FRY9~���+�,km4ln����\����o}B4'�������@����-F�;ؿk;֯�0���s_r��9��S9�u�Fy.�1#!,)V�[�c޽�)%���q��`m�~���9{�s>�1��B6�9��'�9��E�z�`0�r$B��Z���9̨S�e�eR�\^���̅s83өnXM�V=s3��������p�%oH^��X2�jL3���tao �Z�A^Y=���
֌�K�����|���LO���x�'�Q�l��LeE��c�n�̀A�'� ?C�äard���}�+���
R�\h��`qnB�^�7�)6�c�Abx6�ޖ!�־@���!�=�çr�^�{F!��������3fF��92�+���O��k��c�c8�I$|S���@eI����p{=�կA�51=;'{ƞ�y���aq�8"ɢ���Ύ-;�ཷ9y��s�{	'�c�(Þ�O�4�(�?{�3�Ba��5�Y�q;v�cx����6�S���]�L��[tw��NwEU)JA8-�]r���H*�X�u�����Kߢ$�
��?����ȩ���xQeWQ��11��֯���^B���©�\8wQ�:�I�ɋY1
OuR"����l�� /���A�EԌbt�\���s2���&[c�
�^%#�AC��cjx�)��KQ��Q�z���&X��0�IP�P��ݽ���U��Ƈ\:w	�^/y��y~�1r\F�n�'��y�*��_|�!��}R,��vT�������F(��pQSY�ݛw�{�C�c��H(�Vc�(!�rH�X����ז��k��Υē���W`�������<_N��=r1/���ɢ�i#)v3���LM���yL@�b�'/��
����y��'��@�ϭ�Ť�WK�jBa������Rc�YV&1Yf:$,�A1�$)P&'aLV�'�I &W�ٛ��FK���	A|���Ȉ���񺽸4o�-� ��BJ��j���i �y���x����4Ӹ��-�udZ9��ǜ?u�҂Llf-:%�S̲�,�Z�Erc�0��ľ'�Ji�V���?���>v~�[�q���\:�%~�	���x�kߡx�:����36�D�C���,vq�y%)� 7Ο�~A�r�4�	�^���0^��тՔBR�RR���
�ÿ�+������/��~��Elkx�?��5s��w�x�wjL��w�fϓ�I$s��-	���H�5�]W��;�rl����Y���|�o14r+):	�ccґ(|Tn�@���.���0lL΅^��3����#�03�đ�`qr��_e~@��f�V�n�DDT
�ɤ����Ӊ^���Lt�fϦzvl\Ex�Mk�}�f���?�iN5�H
d�ɠעQ*����L�W\�ՑK{�-��%��>�4�8ę��8����#�谱y�.�nY��R��-�������0p���(��.�;OVI�I��N�<"�-��I)zvn6v�E���{�
���� {Z����S����w
��p�:O��/:tb;������(�(�ʥ�ں���3ޅƚ`��d�5��&u�|��\8k��������).dx|Lv)�ӓ,{�h�1V�W�g�$�p��8��rj7�!��2��SX�G��69�g'P�C�"fu�PZ]��v?�J��x$BI^E�FN|z�s U	{�7P��Hz�V�(Õ����s�ӿ~�Y��EE�r������ *eF����	2�lll���N��M0�Ɓ�/�и���Or����%Rr��������L�] `'���&vR�X$��DU�*nq���ɤ�$��ٓ�̞df�ɤ;vǖ�,��.�*,b�`Q�('ߛ}~8�:��E��>�s�k!S���~?UU%�mv��%&[�旞�ء*���(<$���{�ns��9�N	���
�}MP1��.���1���
qq	��ٍ��g����y����3��ż��;<nn�_?ҳsy��gD�M"]޻���IҲc8x����A��n{Llh �3*%%Y"�;;7�\�E|rv�-��.���F��ʙ���\����mb.�+Ryۃ��(n]=G� Z�#0<���]�Oas+(,�qR����ORt8o���̍v��E��-~����Mk��=�$�È�.�S_C~u9r����)t�\�t��{�9�"/��eA^�����{���YHL+��S/������/ �����##5���#���
�Ϯ��-F�Q���Awo'S�3"*���Bn�r�0�,,�fqi��y�"���T����"��M�-��g���o�3F��w���nIDץ�vxd�>���H��?~*.X��v{v�<��\`��� ��̔�KK�c��bc��L<l|�������V�KxOWL��#�^�w?a�o
�6�W��#���llz!����� >6����t6	�ߦ�Ϝ@��?L|b
+��x��$EGs�/o2��BYQ�U��<%@����N��6��JbLi���R��׳����ŕu�.<u��4Z[{�X��O��pz�s�������;��b�v9\����׾X�;�~ƕK��Y]ʳO�pi��*���A�!.>
����ʼx�K ���ILkV�!ɄF�@� m=�7p)�E�����<��\8}���V�bX��gA��ŗ>��݅���wh�h��S��QU�۱FL������>��I�E(�%�����(�󟚙����n^�H�Z��mU�tq��k��-aw� �#�t'O��2^~��g��a���˗/QSS�N7F�[lHڧ�d�*%OZ�u��M"hm���2O~z!�M\�%�+z�(�(���`q�ߴ�Mxyz��SS�:��p�DD'��vs:~z���	Q�P�'R��)����z8��Q���P�?s����=����V��N��<��N��F��`<)^��hІ�b1�����d1b�m��ۦ�C\"��/��W�r��m�����H�/��z{�Uq���ܽހq݂�ˋ�4)>����k?aWe>/�A�ʇ��{�Ǐ
^�ԗ��LgͰ���++KLO�1<ԋ}cC�͍k6�����u<����baņ�'���jvK��@�:>���bR'�1אZ�Z�w�%91]�-�xCV���_ԾV"B|��|���e��.��
V�����%q&F����ֆ2:9#`6�Y��������[���Y�IȯF�ʫ����e����Y�Y@MdB
Ǟ;�&:����dl���S��8~���>�P贒ӳ�{dayӺQ�ZG�zY\�E�����˷��5�d�r��%>��$=����`q�	K��7"�}�S[#�p��u6>�k#(,)b߁j��UtӃ*�h|d���jX���k�g$�����j`rfT�xb�[�}N�ݓ���m�EZ\�u'���|r�2=�+�Av�~���OL&;+��1���s�&�n7x�2 �@�F$�VV"=职��v�,��[Άy���d5�龴4\�����I�.��h�CY]_���C�Bfw�<��qيiՁ��H���L2:��n�Ʀܟ��l�"��v�n�����{�{��a��ML���M뽋�t�Ć�b\�fjb���$�2ұ{�0XMX�F�U�--��dO�&�܌\�h����<�#��.��M#4q���lT��H̟�x���OD�X�uEEp�@%�wg����M�o���ıcO���ʆe���������X��Y`]T���X���x�[\g`l�q��a	d���G�²�؄�*�	z�s�(b�z���v�����o	V)��2;��>���a�o����a�吆A�׌h��ٹ}76���
�2%�!��t�aZ�C7كue���X*K�%/F�������x���h�NL��o�"\���7��$��P�Sz3�O�B`x&��W�{z��r�/�*=]#\��$�3㸭|B���� $&���nf&�X�ae�� ?����k�1���7��{�72I�)�G�8��p�H}���|�Z���y4qI���W��>����^�&��\��c&�{0K�}/U�����aV�iiiF?;��HεE�v�����g��%��"n�ӟ���|��&cݔ"���+�`�r2��.��4�HtT�r�,m��Y��ۗe�Z��4^8���Pzm�^��5Xp��鉏�?
��Eݴ�]zp�^������n2�����25+E�|��;BHtx��{��Nt��ǉM� ,:���5��N�[�S�����y�'m�ܹ����*N��:���QZ]��ܪ�AK���k�Qn�}�r�$c���S��w��ǲ�J�6�����#�X[cU��nr��9��3I)i����=0���<��=�:�w۹~�:&��M������ˤe%r��c��{��b�K�&�P����IܾI�JIX��.������ӓ��BU�ۉ�lD?3�a^�y~���*r����q�^?�����A�j :6F�n޾.b��M�AU���Y��8p�y�T>8�6b´Ąr���_��8Ain5Uy$ą������$w��7����2�
�GXh�p������8P��Ξ�z6�\��̹��0ؼ9|�e*��s��e�޼��)����T++��no�֥�̍t��BEI)	J����}æM����E �?D"5!Ǧ�Ǐ�XX�n�7ŖN��Ɗ��%�}�X\*���?'/�����7x�܌K��'0��<LbB8�~�	��_ĺ�gKN,;�(+�����p���`!W��Ib_}%�*��s��ndMhH4��5&�Y^���WItL�o?�{������YZ���IRB�/����]l�5�~W��`0$�Is
1�,����
����o�=i��x��� BTl/+f���?��w-���d^";'���
�}��mv�'(    IDATKk'w�<`���W�FnA%��c�j��ҭVfu��f��B��щb���� ?@������v�!oK6M�r�����z�oe��b<1��+'9%���A�{�=�:������SAo#c#������Y��
[��kf~��%+m=�Ա����.np������ɴ.@����8��.s��Y��������r���70�'�H�$,$ oO7�i����'����Ac���I[����F'�fq����͆'��&!T���	���R�OO9c��Dh}ho���p2/��zJk��b��TmI��`_���o�`_]ei`[!����;�|r��g>^M��Nbln��ń]�ߌJ��5dr�����I� ��<fdRϒ���꠸���_�K��L����E77ǉ�ŏ�����wi�~�Ck9��n|���g?A!۔L"��Jrzq�1�2c6-3??MWg'v�&2�7.�?~*-i�������� �Ln�pPh�ZwL �����'gE�d�d��^y�=�
���'D|��	���X7;���N��緹x��b�R$-#��;wX^5��ףp8y���T����#n7��?���O(9U�����x�z�nZ.�ޮN~�!�[X_��q���@M4JU5��c0����!�u?`en���@��b���?��Ćk�ے.]!!�b�"y7�F�&�Pz)9�"���;$�=�����>9}EPWW7N�"����������o`��ıa@�`��(�*���1��)�KA� �WNy^��̌���JR|�xvJN��i�;:Y70ۭ�uuas�Do����_��n6r�N#zLno���Db-��r����i������?�ɉ����7g>�%9��tx�ZLK:Ɔ����L66-�T�t�ն����`{`Y��żI{G'��UfV�#SDPRu�����T��W'�D^
Ξ9��� f����a�f?�)��c5.�p�(Ȋ��8�`�&AJxp�gNDLl��%��%�M��f�㒞��nT�.⢴�V�O&��ɶ��Q+�O:������i�5�Fgp��!F�fy�7bYo�;4Mx��&&)���n��`ԍ����q�=��Ocw8����du�����lB.�ޮV��Gц�	S�9��0)��4?|�[o�M��4��0LTF	~1�;�4��)����y|���ML<�E��+G��br�K@�$��K�������O'95�y���A̖:�SSc�=�����$\����:|<�"Z����5���EB�N�1�bL���a���;�s����c��Q�����Ҳ垞����Bԯ��9a&3EMQ�/���8w�}B����#&>�`������$k�(�v��v{11<��G ��t��32ń���ވ��&)���d�x�QUKUy�{��7���o%�a��SMnRk3��@0��,��Q�����)��׎�nƦ�	
���������}�J���ba�����iF&g�]1��LD���66��M9�E%d�$�Λ���փ������ �w���3ED�U���AgK�H�<��Qԡ�8��b�ё~LFVۆ�,-/��v:�����/���YW-<��I�!�iT��7$��^��Q��@?%2�U\rέ�Л-Hw�
_A����x����/�#+��_�/i3��DuoJ�:a4�[L��@%���`��7�m�;�L�[��ȈH����hema�x.��˳�ܚMfr�I��&�-ݤ?n�l��LNZ*[�2���`üFDTcS���Q��(3+..7t�?o�W��=�V7���w��d�M4�q|�?��Rs��c�g'X�¼8NTT Y��|��������m�D��ό��fzZ*6�����CR�j��;8����T��
f`z����CWd�����O>a���$v���q𐈊�O����H��g�����bkIIZ��Q(�/�:f����.�������n�H�о�&n��qY���؋��ͧ�2�
�Gj~q�Р`��yn�?���.���5�)��c�fF��צ���a�u#�4]!:̛|�5�es�%���^�������Y1�G��Fhp��>����g[g/I>��n����
z3i���������;̏��\7����=GAy&=S<�߄e}��(��4���WFXD ���|I�>:؏ZL�Z�_p�X��H��C���E7�#2*���JQ�o�$61��~�G4�����˘VW%-2>�#/<KV^2�o4
)��3�G�H
�jw)ѩ�x�]�zL�K�4�gia���rs		�0���G��z�YZ�1/u�f��k�8\w��U7o�{m�VJwFa���(�)}t�����6͸-��j�VG�bw�_�KѲ�"�jR�"��
�W�bҏ���a�����/Lq��-Q�ц�a7��}����3<1MgW7�-���l�{���`>��<�o?��}�J�s/}���
N}�1��^f��$(Jʥ{S���ݻk��D�!��JeI�%9�,�l6�������.2�S�Y����ygu�fI�ɣ�>5�g�n6�[\C��1;0:�p���~�-[�����]]���#��C~�^�ʲ9w�����b�&&IC����K/�p�:���I�����8�(r�D2;?!�ݱ�I�<��p��7ɦË��"�s�[�̕G�����C��ȌN�l��b�~�<O���f]!04���b�2O�2��Kfq�o�"�gU��E�}�|�G��G����
�[�H�?������4����j�R��ܼ���1d���e��Q��y#��:��n�hWPY}���r�K���2�?_V�f��a��%'��ʇ���P;��QS��BnE�p���Ixx(������9N�Z-�v�]l��ikkC!�&7;�#��evnYD{G�͙ؾ�8[Jk������L�m��m��jj�H�H�`���oa�.�ʳx���\8�>���ׄ���aIGtD(�qф��EL�l�066������
J�QZ���&Wo���;�eSɖ���y��J��%ǪB�`P"_��tv�g��]@��6�/o_5{�/V��<�rRc������kka&ۊ2�v�I��rl���Ax�6����L)�.%`$hDW�n�?��A�@o�8-���͋��T��D���Hsk�o6���L��r����^�Ļ�p�:O�����ۉ��'����)~��!61���b�c������1=9č���Q��Y����ʢ������6s��u��}#�KKi�q�|p�����X��+y�u���061��?�`?O6-�T��0���;���*$wYY�Z-��PV&.]�.<���Y����˟'*0���n򰱍��~V�(�q�T`��Cx�I�uR$]FG��m��,.N���>v�7�A"2U-���Y7I�{q��LOv����������0�?�J9鉤��)�A��J�q�����+B�]��������$r�Zo��C!2�Э�b�$2���}T����V�^�+n�V�a�T�U���*�n�7І��#m��c�"�|��P�݂J���D�&Hlӽ\.�ޚ������Ξ~�}�� 26YPEO|�w�53���M�O��Ô��/�XM�򸱑��%P��GݾZ��#hm��̶L�����[��Jdzz��"�dRMC��*==�6���x	�!/�XH�/^�*:�n� �7uc��SUw���8�*��MTJo����ӧ�[O�b����f������jZC氒�AB��Ԅ@��fܽč+g��wٲ%���dU\_Zbrt���uӸ]V�+E�{غ���!.��ǹ��������z"�پ���'���G��
�}{H�Jdyy�Ҵ8��������������Qє�W���Ĳac�nǺa�у�tu����"%9�Cu�N��֍���	f�W�a!���b�R3�?x��������>�@�LPd�vTQV�#.*�͠Q?��P_y����r��y�3I�H�!��xy�E
L?7��!��e������g���7O��{'���L'.;	�$&��Ef���)�Υ�4�m�b���j	�9�_)4�\NQ^u;�Px�����4��Dq�?�M�9�ɻ��SRTHe�6BB�,,�XX�gfj��"a�A(�����I9�s��#A_]�y�1<ò̓��"�p�6�;*wRZ����f#�>���U����{��"��09f�O����x��''SY��@?�<���u�5�":��++�6e��oô����<�sLLϋ��*6�6���|�B���&3)�?��Ot�u#S�dWhx ;��x�`	��~|��_h�yY��kwV���J@�ˋs�u3������1:6�� ��d��
ǰ��\`pr��q=��Tj�?4���"�b��� ���DQ��`f̀�hà�Gr�JàS��f0�Î,��︝^ޢ3(��%���u;������[���`+JU0�kx)|H��k���V���Xm�{v�PV�.��Q� r3S���~�\�K��'R�e��[d�%���n�s`��m�x�?KK�Cz�|��~N�~x���\�R,(�W��]\���	��8���22����c�,l/$�����x9턫��^��m�xi�/D1�h0b���><%�f������?�g���|�'�k������`�n/Ȋ��{d?��<l��aq�P/!�>TWQ.}�=���<@���W�F�ĳ-,,$55CNg�f��u"�"эfF���浗�Ě��7��O9������ªp�l��u�s��bù�f[kw1kY�C����uzښ0�N1�߈����Eih�}Dq�[��n��ݎJ�&8@�:H"j���SʇKmO	j1)1cSˬ[�,����Ab~%_�����Z���K̰̏i0�ơ�#�T�ˌ����M+S���t��Fz����f��񩏅xT�b�d$66�=������<f�Y��.7��E�FF��7��*������R���>�our��5�K�H+ml��!�$���v�z:���8?BT����UD&iX3-�����i��e�"BII����M�F��$��m����ScS��B�N�%')���IN�n$.w;9��|�Y3Y����w�c^����0��[Ū]Fݡ�B�m���D�˖�x�=���O0�$�R�	ը��cjfO�'
�2���C��*��"X\Xf`t��7n3==��ϿD���{LG�m=S�O�K�_��}��7�cݴ�ʦL)�������N�1�ԄP�֕���JQ^~>
n]�ʕ����h�_|I��&�F(��gz|��Al\�������%'-'Gt^��͌�6�y�y��o�	��W����zҲ���T�P^ZN]m!7������0Y�	���"�~�+����?�Ƿ��Ǿ��:@��=TW�34�͓�6lN72�ݢ�W���QV���%�w��W`����g����ŭ� +#�[/�r�*��%ԑj
+�bv��UG��L����qy���`��
Gy��D|t�����F w9Ŷ���]tˤ�����-���jAJjZ26���Eaq5a�I"B��o�?�8�̢�ČJJ�HL�`~z���>�p���M����x���fb���.���g��F��2�� �W��R�x���Ƈ��?����"�¦�����F��q���`4j-ee��D������N�t64��h�R���k���"����(-�yBC�_��[F�څn����{JrS��^2��(�S�D_X��E��"L�QEi(u�ed��"W����`s��5�����4��䜭��r��c� �t6�U{1<�����B�+I��BQ���g�!""b����ڢ�4.��@{�C�س�6pn�y��.QI��OL}m1a��k2H~N����t�t��bvP^����4:����ʋ��9�.O��?{�z8wFE�!1�]>r
����o�@ss�����KG�Q����'�O��x�kbkR�����,��Y]ԉ������0J��x�����5>���E���=�r9}! ��>ϑ�Ǹ}��;��!� d��������?XƇ'?�����G��L� W*������X7,���MBj2�U(}|ٰm221Ec�c��}�Z,T�P]\B�����[DR�QK?�O�'�b/�����b2��P� �������|�xO:�����z�>2�rD_y}�Dl\��7�>���GwQ�χ�-�\#5)�Ԕ��I��!௤[O7�[�������{�>/�>o��GgY6n�54���EҖR
Kw�����~���źi��P?!��Ȗ�+Znݼ��p/�ˋ�(�}���_��4�����ajR���S)�$˃����361)���f�f��o�
U ��]n54c�BPX
��eK���tv������2�7��Q�m/'!3���aV�G�uYX�fKB$��p��h5[2�����\�Ǉ�hoF77+�����TVH����Μc�`b�*����x%���k$��a�9DJ���{xp��i�G0I�_O� *wԓ��#6�RlN�Sh@�4_"#EMY~�5���Vu����U���[$߄~eeA���0ݝOX][&0XM�ޣh�����$�LO��f�#������SJVv�O�p�<�~�j||U��NZv�x&�̌�,�<��+��ñ����'�/(���Z�¥>�au���^Z��355�C��g�?Ñ��9��Y�{�#�LVF�fq�F�VHfqu{���p���5Ӄ�"��N��j��R�Ӵ<��X/���֗_��(��>DLA�B�j�nQ���hz	�$����ؐ����q��m�6w38k��L|^%q�[HN�@�	z�\ɭ�W�{�f��P	���SάN/(��0��%�����pHC���h�bd���6lzb���@��o%3;C,�fg���|��̴�pp��*�)-�&����?afA�$��ƃ6V6=)ڱ��V���ջ��H�w��p�������`���8J3�§w��IzZ�
P!D�!�W��bh����	�Ż����{�`|x���	��G�z*���!#04�����J����t�v�����P?��尻*��� 1�ύ�����n]'!>��8�N+�9F�G�����ۇ�5u�lɓ�`\�p�Ξf�W�ѭ��M\q���F�n�RPTLiI�M����2g00o4��v�$��S���;b#�cY��v;RL�����l%�����KUP�rO[���biр�ˏ��h�&�t���<7�����þ�e���'�=��9�Gh����M��Q�e���C�����~m�Ĥ6q1�[&1����Q��hb~C�S���׾-l>;�~|׆m�_�~�pz����f��18W�Z�M\\0�`O�o�JBh ����gb��̔����P���N)깆��beq�q�\��Z��CN�𸐪�<��ήY����Etd2��=]]].�w�����XY1����!���x+������8F�@h6뉈��7X,��l��|f����c��:7�cdp��]8��0�m�|�;��uO/~�_�y���FxH0�Yn�?���(.�'[k�R\WǤi��M�:��A�[b�k�f�!0Г�Dj*+R)i�}��7�t�HO�%>6��<�Ǧ�����M�Y������?�g�8\D&��}���EΜ�����O������o+ct|���n�Ff�[0/��g�رZ��ԙO�p���A��R��яL|z:�:����[��j����h� �����d� Av���W�3ǿ��;mܻq�ts)�$8*��{�R�5��?�M_�C�+�Dū)��A,cjv��YDW��$&�SX��κR3R������̪a���%V�$F��T33,5[X�`�n)�)w&3�0-��<�u��4n��L�k�x��YsxRw�8ޒƉ�i#;)���!n�������bI{�_�������၀���*IMI���Mm<ni�{�%S�����:�]�.�Dd���[�Ƨ�OˣFᗔ0�vT�g��~��4޾D�DF������pRg�t�    IDAT�)�K���{�$>>�Ͽ����J�n�8tɽܻ���.��c9p�^�ZZzt\���҆��^�&~�p~���0;9�6^-I�x#�۪8x`����_��2NLl [2�x��!�������ޞ����m�_�`Gu1��JF'F��R1������C�T2�����Vv10�#(1_�%�Z�������-nK��_�q)
TZ��Eӆ���$���Ʊ�ތ8��3c�{�$�����o���-��M���e�|2�Ã�󗳲0������Q		Q҂���NR3�ٱ�0N%�]�GCS/&�/5����:8���I��>�>^8=d,��$�{�Ai�b:k��ܼ|���~�eQ��ʦ���h��*��	�'?����(+�bbl���uv��ǡGetc�F�6N�����mt:��"����,��8s����H}%I�-�bJ�
�������\��)�u�e��|���qn_�H}M5%y��O�����s��UVV�p�7IOO��='@$����on�ot���%�.�wR��!�H}A�B\.)^t�>$�_��@+c�O�K7\n9��|��������y=F����wr��i2�b�(�&2��e�ڊ\:�o��;૯�LfJ"�5~>~LML������(M��,�YQ���D$�jt`�ʄ&dvx���P���:e�;���	�[ŦN��a������/ǅ�7��o"B�<�����hU،�t�6s��Oq���%$��j�VB���<�����@)� �l���g�@L|:����n!|vZ䨢�8�엩�QÅ�wi��(�C�΍={��G+�s�����)*����Q�����E{Ki�RfN����ф�	���,���]2����$�P��ObT[������5�k6��n��֚Z�����ς�����ύ�a�C.�vB�:Ub3���!:��FJ��A�_/�4\gn��mE�<�{�x��gą��jbeQ'bn�n>>,H���nG&��)�s�~���i�z�c�.���)GgPE%������"�K
hm������K�˖e|����K�`*�1LOMp��IR�"Eme��	�%�,u���qXV��L&;5��W�262B\|<��5D�&����⢉��]�<}�O�\����W ��5�V�E���.���1���@�&:��m���a��{":�.3�v����[���{<x�HTD�xF�f'	ת�J�F�g����V��e���a�T�<|2�ݻOH)�aס����<&6�����(�
.�;��@7��eܞ�x���v��٘�R�r/Oq��̦MOJt !����|�arl���~�32��G)��i�
M�t����d�6"cS��s�^3����du�BDj.u���Q@hx7�?���ؐ�$���79#�qQ���F��#��`vf�F�6"
o�?V�[�x\VԚ �f���eo�!^8�9N����K�Y\5��[%(6[��+v�����Q=���߳0�,�A�P)���̌Tv32�����#=|���d'Gp��9�*7����I�^����������u6m����������e3##s�L_���N'9o��yb���cc�H�_ 7/^���k�r�W�&2��KlnI_-'';�ڝ5B%�@$x�V��r?2�����6��u���DL|1qQ���z���(���roJ��HJH�f�d|T�n�[��N��@vx
�L6;�+j���?��ޕ�8<��o�VzS^Q@YN��
344�ș�>�a3���MZfN�Mz��XZѱ�0��ĸp^~����n����{�	`Yw�V���H���PGƑ�����J�~���o��ҁ��OB(+˥,?�X�7��v�������i���ElS�b�jgjr��/;v�fG�lN�.^��+�ͯ��l��B��'#�O�&<��{v���aEzN�	�����[_j	�J)h���f�+�R]n�7��v(�qy�pHà��� 2�fP�3I�_�\Ifv>��I��+"&�����2=�,Ό��߂˽F�.iL'\��f&!2��D>x�M.�:ETh_�◉Պ��{c]|���FY^���+���Ggq���Zr��%qc�6[Q�5+����Ħ�137��� ]�7�n�S�����H4A^��{S��I���=| ^&�}�����H� F)[.�ts�t:���X<<�b\�$b���C�ݼ��w��H��;���;���ѱԭ[�?t OZ70�����~p�)/���ۉþ́��Y]��`Z`i����(��l�&�Cr��O�G͸dJ��F���ʕ��;�(b����
�?KK�B�0�Mr��Y��3������L��09m�icQ{+yt�:�s��L�cۘ#3;���,Jr�Ŷ�ĭK�q��iA:t� %EŨ��1�����j013�H��4K��2������s�_�>��Ff�z�+�Ӹ,�g���žf�������8�sØ���{�P���g_8ȍ�W���I�/�XY����l��������.�pZMb�<�7�H�(�qd���3���*%��Y�w[hjx�����!���VW�(��m�a�5:��aY��?ȃ��pBel:Ml��fzr��g��򔱭jO{���|�֗i|����++넫��f�w���Af��lxi��{���t2O1�kB��MO�p�2�鳼��!xk�1�U�=��*_�[�d&���p��Iz�_!;;���k�D��#z��Blu6ELD&nY��É��ea�$R�#?�������������Fbz�k�ͩ�O�-�`6M����)�%2.���2"�C����'��rS^��Ը(���Q��Q�+�.?�����������Y��åѸ���,�}]�Jݹ�j����s�n7��Gp*5��>��+�_���� Ik�7�U��)/�7~���?�MxL0���K߭[��p�	"H�IG�=�~�}]�l-��?�_D9g��D�s��p�ǣ����LL�2�7�SF��}lx�0�7�Rz	"���Wi�v��5=��!T�V3�f�m W	p�R,�R��6Pƻo��p��~tu������P���(n��/)ނR���Sy������P�m����X���2>�JNi[+�
�C�_S�\��}��|�P�ӭ	�߱_�8n�F�29����'����u�/m����0O�L���҅�b���9�j���_@��˽���`hl�������?�92�*�.A���ts��OD�M���k�h�س�V���n����q�4�7.��ൗ�s������wv��<�t�M���3�8x`/Y�Yx{{015νG�9q��P�P��%r�w0�����!�z>�������!*����L���z.(�UG���n�""c��/�_\��8[�)���A`��Ҽ��"1.�������,͍��G)+�#:2RDLG���mhx�E�E�/&�Dť�q�E{� f���Z}���dn^��ۏ0���nI�h���hN}�.�K���B�4����zkڐ@C;q�V�U��%��������4N���a�[+��?���Mݼ��	q�(y]voR�j�;�9R�p��5��=�I0m��ع���+�]��������_<��mI�x��^��&@����W	
	"H�& 8��J\���6�{Pyx���c�s��5��7�XZ��K���ϑ�������n���$A��� //�AG{���_`$�� %-�����NJZz��n�G kK�RP��HD�r�&��z���p��iL�+$!m>>�xx����'�|v�:6��٥u��F�)ھ�m��|�6��?D�wp�g~���s7h�AD� H�I��h�	������k{}[.�R��εw��q��DO�h���$�bA��$rΡ�ht�����v��#����~���|�_ (UKd#hLJ��8FEU)V���b7�_eaf���ZԲ���w�հ��������Y���,Ǐ���3T�6�P�Ĳ7��q��3�[~>���&֒ZN�����Y�P�079���T�"�YZB��#�hB������:C�ǌU'��˯����
�]��J��IF�����uuMh4&bI��pwp�]��H������	%����uj[���C"�J�s�Z�N����g���˅l��/�N]���X�"'��S@�[���<K�O�o.�<���zښ+Y�ǤS���lf�� [[>܅e<|���V�7v���	Ƨ���Y��C��r����"�=W����xN��l�ϓ��RY[F<$��fou��2�W��233����+hu&�v����l����Ź����ڛ������[�..���A$����i�*�8p�(��<{<Ï��G�w#h-6�.#��h�qҙ��X$����ObP��ݞG�L���E(��d<�wg����1�n���0���<ezb���0�f�	�(j꡾�����*�Q�$�g�b��ϯ\���>%������QH�,���\!\M����LF�ȹeR	Vs�Y��������sw�\gjz�YO,&���������<y�\��q%��9�;tE�>}��F��`����"��w~�!w> )S�4�@��h�A�v���h�������WD!��	G�MZT�������Z�����QZZ����a{{���u�W�`-B�(F�pSVUM��v��Q��|����'�Ȫ4��z�N}�z8�و^#٢��A]��"���F����`��#Gy�/cv��y�?��x�A���p���Q�Y�=V�~�x�m����0v���.'Cg0�K�X��g��u
�����A]>�U�A��'�àT:�ͥɦ�|Q-!	]yї"e��d�ZOcs%嵬�{ɦ����d<����B	�~��t�ǩ�9��Dq��|\B���wy0p��o�T$��.r��q<�%��w������V@mA�٭�	j�Nq��<yέ�>#��G>�@�(��+_��@��o��������o�����";fU���R��Y�zΣ�AZ���O��F)S��J�X��dll�'��Si<u��5zᩞ��c�U����C�b~��37=K&��tiS#�/���1�t���=7NQ���ϝ�l���d��i��_��[��9S��S�.�ı��mf�O�t�	S�T�w�t�362���4K�	{^���1�2Th3�\àoA����:y��S�Y���\�G1�����l�M�07L2��`3�]-BI��p�p+����_䕋����pOę��gie���]6v��.zO^���潧$R^<�&�ܺ~��"y���l����yA\�g'�Y�����14��Gy��a�E~8$衙X��%��y�s��FZ�bve�յ����~��7B��Y�ģ�(�.N]��w����!b�0�6�*�������jJJ,<���7>!�1C�KKKK�F��c�zEF�{��>sKT7����	:w��'aqbJ�\mq��I�7#w��2�C ,G�(���W�Z]$�i�l��[�H)���]��]�p�s��8��WQh��2��v�KX��}yv����?��H'N��QϿ���<z�B'�U�$bQ�޸N$����X2�ζ���vA�]Xgba�ݽ4%ͽԷ�RW+A`�|����<~@:���"]+��)/-F�H��;?��0E[s�m͔�m+�X_Lw{5W.�˷��/\8{��݇�)5,��0<<��ʒ��_x���U�"�۹rs���m,���[]�����ݭ�����bs���L}�DP�`���\z��Ȉ��\C��L[CuU�"�\]VHee!+S#���S��0�e���avQ���/}�h\ɣ��׃����f8��ߢ����@��\�R#��������q��w��F�ٓ���s��u���o_<S�7W��ee�)}���1H��7��oR]^�����^%�����^~�_��0�ɕKq��u��§7��w>d|nWi�O	����� %���7�\��[��3<%�vw1gΟ� ='�

�5�l�Cw>����PWv���R�U���eV��cҧDv��o�&��*�KT��T:=*����Ƨ�1��9���)(�ck7,��T2�{?{�t*�L&'��bw�x�������ߠ���T�χ�Edo�
��ÝM�ͬ�����l �	r�����'���RG.�$/KKD����W��\�����;�uT:�(��L�E��� A��x��6���#f$�(9��4:���%�EQ-���gq	����~���]���[y�Ŷ	x��][��ʒBr�4S�a������9EnY}�ϼ��~�˟�fya���3�L{w?:���Gܽ�@���������ɳ�h:P���-nݸ������'����o~�k�>q�w�67o�����
���`-�T_��b�7Z
I�u\�y�;w%��28��?�%:�6�������Q�%۳�H,J��.z�z�:�\�>'K���{�T0�������'�Vo�Y��w���ζ�K�K0덂7 ��}�)+�`h�9�۬lEI����(/��kmvb� �;kt���K&��?���`�G�xx�S2rVG9h�8�2Օ$2B�i1j((41?3���VuY|}>J��Ƌ'����N:�{��φ	z��S'ɫT|p�*�MxIf��X����
nAG�I:�H+)pU�����%HE|`Pp��TU���$����{�~�#Ԥ(���F}��B��|��M����������A��Ä�	������Uo�{���mVwđ�|�(�G�b���Lk�f�<�?���<��R���z������2�Ӧbb��|�b�R>Ν?��"g��-B;����QUZ�7�w)((&ʰ���ҧW�[�eie�յM�Ѥ�����>v��jȳbT�eXV.��>c�"�KCK��̹׾L���K��T�^Cy��چ������MtJIj1�內�������E�Ϝy��C���rLL�q���F�]���Q^YG��4�u	{v57o�c��=����8�6^x��ʺ2�%�[*�*�dO-�n�,++�r=2:Jg�!Z[�P�Ռ�<����W��#}'��\�:�ñ�	ַ�К��f/����EdG�F��g��O�AZeS������I%(����o��\�ǥƬ�o2;�Tc����h�R(���4�����@*�`bb���}�'���.ʙi������\�VٴYZ��d���׸z�S�R��A�����d$
��4�����ٳX�F$�a:���S�O�+)��$_{�E�h�6�+��@��?���C�-����O�|>Gț`���1����X\NmG�2U��T��a���+��l@��j��NC��#��6 ����)q��$�>��k����13��F�R&�������))���	G��{���K+��>������E�.�����45	�h&��Ώx�l��dђV��C}�?؆E�%�_G/O�T롭��|"̕K��ʇ��I�x�ͯ��_%���>����)Q6������)��Dm��1�8p���-x<nAm�)�J�}��q��~����(��<y���idm�ݼ<����\Z�L�r\)\(��YI�̣�*ȥ�ȕ:�t�((aǻG6���t��X��������̈́hm��@s��K��[�:?`��5\&-F��"����Z
�V�����"MN�I�ddf6�2���N�NC�AnߺÓ{���$	�ZG_{���&���^�gt����ZJil.���F�˄1����-�6V��5	�/�-�*��"'����0ã�̮� 3���&���?��1	J��ӯ�@˻?�)�R>/%e��6����NI���2��^ecr��"3�x�=]m�tR�ƀoo��?z�m��L�iL=M���,A[\]Y�`��rW02:���K�A�89|�M�5�l�'����LD7��{����G��t�<�Z"@(������`mv���Qf&��zil��`w���AM_G�(������ř1���l
S$czzV�}��9%-]}��7�����!�P�s�$ϟ�1pk ��
�\��ACO75�0Z��}�L����0I|m�!EC}���(4i��eJ��������مڨgv~����    IDATR�URՄ݅R*L�ꘘ�`vj��������
�~��;�H���$���=qP��ay~���cwv��U�i�}�jj*Pk4���{ %@ڿ���R!|�4Do�#S"zĤ����gq�˙����N������ u]G�+Ԣ�C
�WU������+�\�b�F1��9K�hl��:9�Vd����t�����2��o}�ћ��:����)��ͤ��.������	�������'?B��lT�Y9u$s
6�aFO��Is�i�J��
�E��'��#�!��P]�<Fy���u�r���7��}A1���=�͘4y�V%VC�+����<F��X0��b��ɓ4�6��������ywy>�@eC'Y�������¢*|A~��/����© W	����W����zd�4����33t��R���� ��������i�+h�������I�(//��`4������3�#p��!�V}DR*�;z9�ʛ��f6��ROO��B���al�&��-�V�5����YJ߉����Z�������3z{�Y^�f��M6ז(+*�k_~���"f&Gy<|���a����ꤡ������6��]ane�����q��Ȯ/F2��@s)�+���g?C�I
���Q(U�4����Jr	����1h������W��(�K�]��СW�)t	�X[�������!H���6>�~��>�K}s���[DSJ���d��*����;G�BH:_�_9Gai!�L�pX�������[�cky��M=�E{c#�H����_��Q/l�&����Z�+�b١К�ֿ��g�~.|��Y+y2�@:��j�!ShI&S�dyf�G(q�Z���� �|��L���Ampr態�V����i��� ������*�Ð����o�yE6�����7QI�)d�������h�~���ܸ+�zs����'<���?|GX�y5���x�M��"r9-���~Y�\��IU1GO��� W�����_Y[�7�rE&½k�]�����?�f2����d2	�n�[�l�����_��+�������"C#�<x<��V�p4Cb?E������X�$Ry��ppD,��R*������V�k<���\��=��0'����o� ��#�8�ن�eC�P������;w�Q�h�o����t4��Ș�Iųj|Q9��(���t�@E]+2�(O���>�@&�������l!�s��%RH��r:'GO^����x&C,�%&dE��lT���]�k���4�m̑��p�½��/B<&,��n	�aeza����B/����=f�7Pl=s����X\%������<gx�	�\t�f�r.�|���Z����471?� ���oV�{��Nn"�'�����O�~��AuM����%����2�����{�$խ�y�K���B�Wkl��J�|~���U�6�H����q�X%�U��I�v�D���I{��a�9@ǡf�$��Vgf1j������5�Gy69K0day���%bq��>Ù�_Cc���%�id�Ւ[>�<���t�ɇ�!UR(��"�Aϙ�^���Y(R�D&)�Es�t�����Q����S��5|�kQ�BL����L4�htr���T�v���gx�O��x4:���.vW��Z;z��n�(���޽!b�hUx
8{�$�x�kH�ź�:�\�Fo�+0�dL�����#��D�'���*�Y���1���ꬌ<��ƭ�l���@$��������h�NA/U*4����W���$ϲ>͉�'8|�O�����>�+s�U=�@u��Pp���-u�^*��4z�$�D��bV��M� ]g3j�~�����P9�8���Q��.�v���t"�Ne�,J�r��5B/h�
�M&±�b�JEMm-/�}��,�GR5�A��a���Z������V�����I,���8�P����L��ӄB1�?Ϩx$�������Imwc*,������fjj1i�T:>��un^�G2�Gm0"Ө8q�'N�w����I"�% �Ǒ�"����,��`p���"HH<I��-�*33K��m�J��Og�ipU�`t�⩬vm��%�%J�֏����$�L��\��m���G�۰�@���l~�f� l���L<y$b9[�k����q��V�{�Lβ�3xo���U"Q@a�YT��l�����'���\Fdu
�d�ZK@�f-�GD��m��ڤ���?�N>����I%��*�"����)qy�fe����*���a��q������r�,)a�C{��=b��}���8Zj�i���4�4��85F>@E�L""�t��@6�6��1���m'+�2<�Enk���k�
\|��f=D�L��Z���:ΚJ��@��298���z���e����gz���y�R�7��ңT汘L9��G�L<�bf~��V������&Ʀ�|~}se'�}�m� �Ȋ����,�P��Ae�!J�멨*Ǡ�1r�:c�/�On�;_{��}�+��*��%",���Γ �2��O�=���zq!�Jb=��2>�z��P�u�@�����Js��B��J<3��e�]����9�y5_�H{�	��~��N����$��1�p��g�$�>
=N:����`��P���]��b�B�M����d��QXX��YH����L��s��'��~�\l�kۘ_���Q(��F1���x� �GZ�A�gږ�Bv𸵴�SQ������(s���������x{w�ACsK#�e��6w�%�����"eUX\n�1t��@D�����9��l��؅Q'c��uF>���b;���� K�kQe�vy6>���_0�GW>d/���a$��Ɂ�^,�*�,�%P�=9�%t�B�O��rY*ˊ�p�K�7�Ew!�XT����XPF��W�g��2��P�3�,J�l/K��_� ��_��N-���2v�A��R\����W���ajz�#}�TT5��Gy0:���:�[a*;�P��-�,N����Տ/39:L*Di��EMkO/�ͭ��k4*0����c��<���M�5�q���|�ǵ+ﲺ0!ȖKs|�����?��1�%��
�+̮z�\���!�-�w�˸J��)���T����  ��rT����	��^JK8|��ՕE���?��8IQy!u�?ԃZ�#�!OE��Zbjt�s���ʅs,//���ʦ��� +��Sk���X*��
��؉&�ʔd
RR��jfr����I�{� �}�W\ʴ�b=�?�B���x"!����-����W��d��v�������P4Ȏ�ˎd�E�sQ�����DJFIi5up�Jؗ�%�n,E}�����{��
Q����.)���i4H�j&�'ڣ�� �Y��û<�{C(�}��u���"'.���,�$�V7Pȵht�ֶ�uw��ѧ���p��7��լm�O�H$���W���O������BA,+�.���a��*@Zu�el�/r��K���PX`��������V"R�X� �M�� ;O�k�������z�1��arU����@�H<���F�U���f���3��ev�&�|<(�]��f�����/Q� M
��3O���bo����((6���79����Gw�����l��-�������Í�dfmc�/}L�W�]��������~J )Cmvr��k�v��H�Nmfxh����H��(I���e���~��<��ȆZ��G?���$�����Y�d��%��[q[4����I�F�V��T6����J*�؏�X��c��sf����I쥰yjy�����C"#=S4ܿ#e�&�]2��r�qz�����K8�Ud���m&�ާ����];�N�]���kK�������d"ʻo����"���
M,/,p��'|r�ᄂ��A:k���N�}�Z4Z5�t�T2ġ�v6�����-==mD�~ݑ�%��.##3r����εɜt)R��F�%nM^Ż9CKC)�ŒM{���]-ʹ�V��mvs�����᭟_fq5D$�efz�pVG����^c��EŢ��S���'ܻ�@TV�76H�r�I����B���p�)*r0?�+���i����?���$��aP�����W�P��ݤ�T=2�x���]���<|���/�i�"#Sc2�D���{lI����X�����ǩ��Ι�P	<�ұ+�xw��%0S�{�(�)Q�bD"�/�ۣ)�6vŀ������{I�Ê�F��OQ\�D2�*�*��$�Q*�8�\��Cwn	�������?Im��:�J.'�NO&p9�M���@��M.Ũ���N�w��F���B��f��6BaD��Ñ�<y>���6z����C��ub���I|� �T3pw������aA]�ڬ���9�������͠ŨJ��=#ٴ�]8���*�dR�6��b1���JQQ!�P���f�?8���{^����������B�B��316.��/�B�%�Is��i��sҟl6͞w���B����*9��6f�BP�3���,(��J�/�.?&�~��q�����������0��^�SV!�p�a�Lɢ�1i�ܸz����	��ɫd\h�V��(�L�4��r��)
�f҂ЯU�Ľ�jP��ace���B����wY��h�[(�
~�7����w�&�z��'r�E����S�XGMc����*�J5ׯ��ڕ��biQ{������#=�E&EA�N���<�&��z��������w����8�%9�O{�A�$Ǟ1>�ē'��bXʚ(�j�^TBIe�u5�fT����o�ϓG��2�:����>����Q���!��}��$.����
d�+��bQT*U�$Rpx�՝=V�|<dwˏBcBc�bs�)�������5ԡ�(Iœ�R���t4�B�%��e0����H������Z�X����?�v>.I�r%ټ�&!��c�K(�����Q�dR�P�i�8��l��e���ZZX$� ��3߽���8*u��2	^�ͤ��2��R����9o]宇z:hin���C"�du�G$�b?ϧ7_���j;��+d\��f��Ɇ�h�.���2ZO��F���s�K]l�-�Z�9t�
�]���[���ҹ3,Ϗ���(�rN���HPҢ�Z
��Ih�L�m3�`����ƃgp��Q\V�,�僟���r��2U:JiC#��j�]���r�����6��x�7_C`x�a��R\RDE�Tޙ�/����A<�R<�2ҩ<r��H(���IVqB5��gh�9�?.g/G�SQU� ���ޥ���"�Ur��Z�'��HJ_�<n��J���4���[�Go֋����r<.ze����<�S|p���;��:N�>�ٳ稨�÷ae�'��+�!R��YJAq=%��LO.��'���dopڨ�꠬��ۍ�h&�0r�K��$w1[�44��Z�ٮ&P�,�@C3W�\�ݷ�A�T�L�HgS8�4������y6���Z�����$���?�������8�{��Y�!��QZ�"���{o�26�o��/�ƿ����G���f�=ݴ��������k�����TMFt�(�'��-��+��6�����\
D�|.G�����<��~Ddw�l\��1y�aЉ�YJ�WI�5�
d9�LR(�n��M���Sn_z���U�&���;��bT���XkT�9����2��T�]�~0��;�~{�@����m�lq�L�5V�+T���X�� '��6�Y8�}�چ&�;��)(/- �0x�&�OFD�����?�F}EZE
Y&���wx22�8���M�ȹ,l��3L-{Ţ�������ڈƳ�����y�'?a�/6]z���B���L<����b�I o����l�R⑞?�t�7S�q��eVz{y��C]�;���6{w�q��=�/l��������t�'���G�+Ԥdr���.�C������&v���Ç��P[
�2�dP(�" �q��eH�S���n�R�q2�|X~���Z�T�VS^]%:��r)w�����T������j�3�h
yN	9�p��r��Y���{�u*���`��N��"��A'�����*Oue�P�[k޹���Sl&��K��Pj�XlVR��蕒���3����Z����j/dm�K*#�`��rw�����<7>�$�#6�MX�E΋�/�3�9Sr�������H�C<y���٤�����d4��(��M��Z����Q�ӟ�##?Z�d.�`�B�H�sXmv��$*��D*�^�F-O356H�Y�������s�4z&{	gϾ��SI4,mw����IH�'��,����ٕ�ƛ�H7�Y������(?��;$�iې��x\�"��"������� �~dZ+GΜ���*�U�67�O$e��x�2/�&V��W�x��TJ�SQR�fḁ̊́�ޢ��EOK� ��6�Q$4U�`�(��Jgj���'���RZ�XX�r��s�>��P��ác/r��<*��p8��l���&�N���d���#t�����E�(�r�L��}�c֗'9�X��ci���t��?|O��1����\"�Z!�������ē<~>ǭ�'w�ؤ^�3_����T.�F�!+��Ń�6T�4?ɏ��EEIp�����Ҙ���8���5��%�KxC�
�~����4��q��'DB��o���C��$���m��NN�>�?�ʖo������!V��A���9�N�#�WMd��_^�����ܐ
������f��=̱S�R8�h��X�k�9E~נ�q�x'�\E6Mt�K~$���l��掏�M/>�tF��_�����E(�����VoDġ;wXYX����M�D�H����	��Tjm0jD?f,�O$��;���e��܅ìE��E��ﳱ�eem���[�;h-Vj�hhh�����D&%��(�e�ȵ
i!�A�V͵�?f�������.���O��|��t樕��&+W�\�D5�e�K�a{��rq�V-��� mV+�g��a1D��o2�����
�4���)<��HZ��ge�T:�r7o���!�Ѹ(.����k4������R�Y�t<�����%cbb�XdO���N�cţa��iTh4:6V���N
�i�D���Z���@{w���J�L,f+S�'��އ�v�hlfr�'_<E��cēI���eJw	i ��,R�E�A�	aP�YtX,&�&%�:���Ǭ�.�PWO&���]���i�|���.
K+P�t$�Q�x�~�e�۹���<����K�+r�
��m��aQ�#ak��8~���
�� O�QHK���J�������J���w	����dp�Nɉ����"��/31� ��������&ZZ۩���bף��Q�h5:n���G���*i�`0*9,e�N!/�A^�?��K�|<�*���e�Pw�L�ə'�����������������(�s��y#h,�TԷSY�DIE�����)��V�B����/?d��k��[c0b/*���I:;Q�S�2Q2)��q���iף���gR�����Y���,�^��W�X��	�Ɋ�����6:�:�o��5�T(��(uɒS�0j�bM��&�b)&��<*�L��lY��k>.]$�*��I/,'���X���qV)�H�L��,�AIZ�"W(�������L,��[�x��$�Z�BY�Mx���hm�E-��lt���� IjYV�E��T4��[��� ���T�S�ڏ�]J8����]�G���.�&w1ǿ�dN��XH}l�`��׮�0��SFW{�KOG����o|��B+�g~qV(q��������Ս�J��/?��ξ�Қ^�:��*(��A���~�-	�/x�Jj{�Q\ۀ�d����,���Oyt�ǘ)D�_��++K������(l�v��P,�{���k디����d�Z^�`d_FFa�ZzN�UK}u);�\��'�}/w���gds*K�=G��e���bSdP��\�4���!��#���e}M	�%*K�hR��	����R��b�45�p��yz#����H��u�gV�[ݦ����C�h�.�b��W����[��W����f��j�d�t�ML���|x���2�}�=Mme�5����/�9��?�`�S'���2�D��-����V��͡���    IDAT0f�d�;�[����QU\���c}~��~���L����a�[����ۍ�B��2ˍ_��"����:v6����	Oi	�x�d&KEU㓓\���uuu�dR��>O��	�4T7���)�2%�t��L�\�v�B��ͅ�|v��w�lb�|ҏ�ȅ��Fk/���W�ʍ$Sr�×�2��J6Nm�G��?���+�_�n6p��a:��E�?��s;��&����vv|LN�3>� r��mb�R�����\@O��]֦�r�<F��h2́����w�L�Ȥb�jj�����}����W�h�+�pG#���#J����d�i�VVY^�Y�hN�ܚ���=��J���(f�&M��TFts���s;�(5:&36��ޣ}��8"a�U9�J�B��{����]_��⑔�za��ʲx��E�׉��,�/�������̚Gy3���QP^O<���X*MJ�e��
]L?����m�k���V����������ċ��J)*�J�J@.�:�ȤUS��SUVHM����%f'�	���G���±!S�!��a+�����RJv�x<-.4F�Y\蒱%�nV���%p����tf�%E5�G\NJ邖#,>LZ�N3:��=�:OGX_[��xa���d��H�r�|������^����-���F����HA��].sS3ݸ&��Lf�� 6���Σ7J�$�lV(���T)��,0c6k�@����C	P��#�œ���L_�"�DKs
�Y2.Y�Jp�kD?iF�fY�$�	�f<�B�?B�QQR`gm�)�L�g��2?5&�p��:T:F����^����`8!�3��(-������\�O��D�Y����%.4���uX-V����h�f����R,'��|r�O�Qy*�9q����"O(}��8e%eL<�����hm.+�teU����1���]��,ܹu�g��p���/���i`j�>��@�x���{^��ST^#�Ǧ���0g	m]���=��R�ֶ_,�������6SO'��ddɑ�E�8���3�ٗ쌊u��\+S��y��r��YY�d,�,�F.>�Rwc5y�s�P�����\�1�R����_����~I�������fb��U�07�[��W.^<���wD���QDZ���שilg/#�N���`A-���a�
L���P�#ܻͳ���v+$ℼ;�8��?�}T:�D������w��9t�<����d:1|��Ҁ� -��}�����29⡰�Hv�ts��1�@�K]��P�qX���r,Z���ĳI����tz�����FIfr��F���p��y�L:/��y�\ Ҳy*������ט��&���5�����g��h'$-J�j�ҥ=!�WsX�Z��}f��m��n���\�C.��:�H8FVz���T��QR^%^�Je �VAN�<�C�ӇRA4F��+��y@���<p��\t�=�9JmS��Τ��$�#�"�А�!je�rI�H���˞o�t<�R�B�M�3N�JN�� 4٭�VRW�DiI)j��T*-~gRE�%r���7�2�pX��K�F��7_�����'�A���(
Y�,����X-::f�N�.R�h$�O`?���I�7	E��W+��Zojl; 2]����z�X}z�#A6��$�F��c��b O������#��n����nc��(-tP\��b5��h�y��133)T4i��4�W�e�� �-+-*���J%����_��r����~��ގ]�Z�Fow��#�a�����'�SQ)�)QզV*�E�h�J�F#��]1�Xp��؍r�)Sc{s���=6��X�_ejj��Ս/l��"�����AuE5V��2#*��29z��;7��G�Hg��H����.N��G�ֈ�F&A��`ө��2ă^J<6�z��D�p ���O�3=����X&ͅ²^��IIy�Xj�zb��|�ɂJ��?����ׅ=X�ס�p������T�F�Z�6����q�A^����2����'��' ج`J�VVS��Dck�5�d��u:�J&�xi�!ى�2J���|�����$ȨU�$w��k��0()�J�{�I�`:�߇A顑KA:#����G�b�B�:	��͉@�4�Ք�ᶘY�|ƃ;Wٞz�\����F��Z��)��1���EXsuy���-ߐ��$E.�2�L*Y�����9M4�#�ґ�g��|���8эmr���������N4-�l���>����מR^cĤ�bQf�l���ʊb|�]Q�jw	%�y6�w+���&���S3<����G�o=��]¶?@kkF���|���.�IHJ*�����U\�E��'��r��w���p��AKK�M����4*pf����r��Y[�
b4�`f~������Kᨩ��� &g9�ɬ��I"����n��K6�N
iߙW�0��%I���&��q���v�ו�:�=Ý�7�7c| A�8�	mI�B[���I:�J�\����R����?ةt��I�Smw�jME���� "8��Û߻�g>'^��pub�<�{�����k����840U�b��m\��}����0��̠9U���$<����0����Z��]^N++�ءC_�e�t�1�i�|�{�Z�/�v
n��wo����0+p�������'�+���0c_q)�����4���LGڃ#��t�����¹����%���g�з����f_^���v����}x�ċh��c�ï�hV�t�">>�F�0+����c�p왧���T�k8�0��?:�����d��OűG��Ez�\������R�n�fg����ƗW��������똚?�CG�AmjA�y�T������T;wWq���cg�
R����t��,���8�*4�.s�$I�E<��ݜ����R�p�˸p�w���s������#�0�<��F%\sp��5�o�T����#�J���ۜ�"��d��O�������đ��$�!�=�4|��;cRd��/XX�o�N���\3���2�KM��6��J�<���p��])hڽv�t)"����H��Q�2�g~��~F0���\>���>9��_|�r��agwS�榰43)r�Ͼ#�����l��4��T�,���~ ��������p�����ُQ�ُ�=���^��}��fBc,�C�=����Y\��]���
��I<q�Y\��ͭ���	��\�<���Iw8@���Z���,᝝��������h��p(�b�-BKsp]J{r��i�����Q.Wd�D�{`�Q��[�p����g�����23�S�z�j�b��e8�-EK����s�S5q%1�jm!���O5`qaIv�m�o�uH0Tq��
�}_V6$�z>���fswn�ƻo�����H�pu�w1՜�n������`Ё�ǰ��q�e)677�3r�㎝ĥ}��m��t����rZ~���f� ��PMIr�\n�|�����g����eƅ�q�PCu�2�W13��N���b8�BK},4k��5x�LM�������̾��/��������`0����o~s�Q���%<v��<�Z��R)`��oi�||	�y_d�yCG��������w�%�y#�T�z��;���ٷ_G����}�h���������A�����K��/^å�_#3\\����7W��2L6����8z�)
�E
�������ƵKWDA�Nn0�����q�ۧ�u�S��2��3%������ߡ^)<r�c�t�X+ܽ������O=�W��}�?o�sr	���}�U}�E�ZU�i�Z
MK��U�ѣ{�v�6���K<�)�67����M�#6�r����.4C�{�bR���u�ׅe'ط��|�z��8�nn��k�{]�s����?��BqC����=�(cva�a�Vg�&b��q,w�Q��Ӌ_���>Ġ�E��y����o��6���VwA8�fb�J.�S�w�>x�춇ȹ%x��w�	�M��F�B��i�,�f)凱����9}_uU��/]���.���B�}��ߕJ����l��E��B˸^��N�\C�X���̜-�� �C�FW���0�%��i�3T.����8��o�8p>5���N>����H�X&�(��Q����-K����+h����o0�sp�"�	�Ś2D��`q�ZJ�d"�]�ӄ�����3�Ņ���bƲ�����?��C�B8�%�I`D�-
�!�����Φ8RrἎ��.z�.�]h%��/a��a��Z�h"�Ml�)]�h�a��8���Kx�����7B�x��S����<�+��:��کaw��.�Q���ijZ�-x��7V�����[���~~�Q<��	.s��Q˳���%�)�K�R��3o��O~{��-i���2j#��X�u�?���^R`PjM?�ùTJ�-˂F Fg��<oa�E>���y<�:#���`�����Ҙ����G0���RUH�(�y	�e]v�����/�D�j��,;�#�>�S�~n����{2���e;��2��1�D�>��\(7����߬��p��t�JSX�{�T�zE�4-�9Cַ�Jzf�?����3��r���m�Y�?��wp�������..���Qf����;��������`��Ԍ�h�T�����i(��k9�t�y!��2s9��A$+$r�"�Y��N� P`�`>���������F1[���&��=%LUg�n�1��<������
��@0���O�K��sظ����ulܸ�j�O��{x��(�9����k����;�h�0��0�n�c}c���#8|�I��)��>5���������_�+d���������A]]�����~1�g�}�+��@��
Ǟ܏o=�����edqwm��<��i��eg$A�����6��>�B����鹣�5[�<{�aI*��_��W� � t�?qˏ?�A�
۵0����
�����k������w1;?�#��Ё�(�mxî�Z�������ܺ}�or@|����8���0K]�*4��e;b�l�^�;?�;l\�����+����Igp(ҋT�sqꊦ?�Mnm��w����m),f��"y������f��/�|.��te��]�;w7�&9�#�>)�kk����t���J7,�rX8|O��h�wۻ������F\���'�����vY���B���B�����޸�kW~�W�}�jY���� �~�3��ɐ+����'���#�yvZ[
�������s�Z]�u)���cϟDb�z�<pp�J0��.��7�a��UK��c�H��.I�X�u:%2^��`:5,�}n��Fv>��2��������m��/��ۗ�[HG��OU�N��(����f���yh�)�-YGv�z�mTK.f����c%w���Q�]��W�d��v�|{�@svL���  '�9��$�4?%,�O~�S�\�,��-ג��O>�,���&�0��#][_���ٹY��6v6�q��u�޾���=9���U�ea�)O���a�+"��|�U��g�0%qC����:^���9�Y`ԧ&��/ _*`x�k�'A1��}��!C\��3\x��+7E�j���{���o��n�]�׷Wax��S��'��مS��e:��Z���7o��d��y�>|��;�[����i����;?�3�Qq�!g�Nr&#4�y��ކ����J0Ҙ��"r���� �tD��!2� ��zv���w)������G{w_]�J�ql�q��d{�헢��!�b�b
X�)l{��7g�^���dg繋0�\r9I4�N_�Ȍ{6�1]�l���(Z�T���*{M}y���g��e�<g��HBҬ� 0���tC�*Ed��(N1ۜ���U+<�t(��쀕u�R"F�l�fc�#!
(���$�x��O뷮b�b�y���Cz��RC�y^���9��v��0�eypkw �����54�6f&J������������҆�x��h�����D�3��[8v�	<|�	L�,"�u���?
ᇉ��Ӹp�|��9�ww`aAx:���2��>ݐns���uY璅��y���c����_����=z�v��䧿�[�E�n����e,?�8O�-A���KAp���yﭷ��ի�J�|3�uq��'�ҷ�W]�8���*�2�>�i���ߟ��^D���ZŖ�f+�ɜJ����O.�X.㹓���������Cx��{��c�c�	qg�3��x==�[k+�7��/��#G���0E���Ԯ������K�6�e/(g�4v����T�Q�C+.J��G�kw�{3����$���X�*(�2���XviҌ@��vѪ��r�>���;-�}�m?��^|�mj�����,�ٝ�,Ң�_Δ�o����˝%�%
alpu�����W��9G�?G��9�\�ę�ocmmq!M$q��N��O<�45���;K��&-�#�iip]�[@� #A�f
\et��Ť��6���YN�EI�Iފ�A�!K"�,6����8����5Ae���"�~�e<���/ql�y�2�������c�!�"_v�y�aᨫ�r��mh9���ER�N�h�4�Mb �'I�ߞ>���/�%N�:]?�g+���F�w9v%��9�(�A�n����-�H!�a�B2�*���3�5��3{qf1�s��j�Q��e������֮�X%Ͼ�<N�8�$̈́T0h�2�g�:���������AG�GwI P͡�L�RA3�P�����OeƔ8��4���-����*�߾�\|�4F�-d������i��0��}��Oa��%qPN�6�_�w�0�a��tMGCvM7�jm
@��:�G��G�#CL�f�l�OL�Z�F�,J^���N�Q���d�������7���޴��G���=�&������$�~�F��⹏0�{hw�����V�� y��T(WJ(W�ԧ`J�4�j͚���2L��Z�9_��������s�Y�Ӑ���w��O�$�8�{��G����t�9>��n��X�h���^\ίNM7��CB��"��f޲,C:��3Xp��rbV��N�b��A�'�C�A�A�?�>����l����Ƒ0od�@&&�͢ '���8v��fa�J ������6�4��}Kh�r���g8w��ܾ�G��W_��OC��­[��` Y,�[F׋pg}��������#�Y �q�a�4���Ltw���Y��W��ھ=hy I0W���҅����>Ǖs?��G�����A�8`<��7��KR��jS�t��l�D������n�����>��ӝB?���������h��/�k7o �#h���c����O#���}ع���>��<�W���O>��Ρ����caiq^��h?�B�e8����iw����A��>s�G����{�!c"g�e��>�6�0UD�vg�3l]�]��o�8� o��{�X�B=���R�b��w�ᙷ�z�+e>��j�(���t�f�F��������as��E �)cvn/��9�
e)�XLp���o��_�����5��ҡ�x��s�W����F!�Q)b�\@<��k����s�����/3EX�;�(la��5<��1<r��z)n����g����_~թE�VqJÛ]�\q��?:��E�Z����C�8v���;-	��Ղ,!����+�q�<vZ�;l�KEq4̓��^Nv2S.>g[XTU��rE��.,��dp�"At{J171���&N����]�
=�F8���T��E�ș�?�S]�$A�4��&٥.���0�dL'&ꘟ���z��lmo
��{�pw�ϠS���lۆ�Di:��"��jL6J�2?��/����S
Z���o�9;��h(�d���lkgK$&��q����������b��Z���G;,��bjf��Cw`&D݆n��Vs���6n�⍟��V�rY���,��^@�ZAw��KX:���d�y    IDAT�87����ﶰ�vw�ޒ��v�rO>�4]`�*(T��y1�ѭ*�yh����8P�}YtB�^���������]�/L��S��˛7�'�G?��ؕb #@ܿ+c8��R-��	<��1u���,KN)�f�<K%�[�+��?��#X�-ǌ���۵d'
qf�>�)	��J�J^���H%�%�WJ�XX�\	so�����@��(�\DX_�@'�����p�e �:�Yl3�x��V%)lǆ��0z��j�y)�L�E�7B��:��VI��M�&�9���G}x��ցJ���G��	��bC�\�Yp��?��`�]�Y�4#Kʱ�7"+__B͎��rW�+0��cvi�������s{eޒ�D��5e���>F�6
�	۠{n�V�bks7n��>+�q��ٱÇ��Fs��N7��V[���	��<'�0�s�|���8��Dc=t W�^���"^��+X��Ï6M�^,L��/�`��Vq��Gx��2�&���l	�?�痾����9�{����b�:%r���0��F�@�Ox}p�]qs�8*z�{�q������P��)�	�Z���'�[}|��E\��9ڻ�m KP�mt�鞜�^o����p�GF���N7�vǇ�*���<�M��,4��~���O<��#���9�.}U��|/~�a��C�hu�d��n-�Pt��ק��F}��V�,\^�ڶ����!z���?�x~ݰ��[�xʴŊ��2F!I2�w�|�k�!�h��\�
���	�$�ƙ�4���k��(�]؆&q�,>��,eV�ɉ�X�'�S1Z��b-F�׈�$�lf���ζ�m�)M���P�N �/���!K�����v�;�G���+�f�$�K1I��䌡��9�'٨є���p����������g���D�`P�1��O��m!��0�ɱ��D�g�{2����G�$^,~!��I�3�N�=���ή"�%�n(?%x?�7��Zd��X?��c8J�ZY�F����A��A��bڑ#����N0�F�[��e���T���b�I�e��,�M���Xu=�}y����m�;r��s/>�g�;)$4g�I��弄87t-&8���jS�����C�a����+g�����U � �|&��w��M�q��N��׸��w��&��	���N_�I�=��q���w�!2�{IM]�F�+c����>3��1�=�� ��kk��)�EQ��;�$(eN��0hL����ܝ�����Y���r$���=sx��/�9�@��2	�p ��X.]�r^��$���F.�yʤY�� ��G8�w'��9��	\�"j��o���/��YI	���'p��CB����<9��U6Bɻ�4��;�b^+g�uLy&1���� ���X[�A݆.�S��e���\A+����`��;��$��);�C;�?�k�V����
"���H�`�	���1�܋G}��"Jy=�H�qp5��i����sXh�z{�]�~���������|����OΟ���0=��f�Ki���7�R�	hE�>��)-�J� �������ϟ�e�����b��OF� B�4�oq7���aw�k���x��������'���g��(��mow��`Y�I��E��A9H���Q�:u��_�����//#�"�2���FazZfV(�K�>�W1ˎF����۷p����w�X����U��$���Lͥ(O/c�Y�M�^_f�\����{�����x��_b��]aǟ|�;8��	d%GVKP�gY�h��ӵ*feܸv7�|.3:�NK:J��E��AwM���u3��m�<���>4&g�z"3����j;[��[�1\�D2��M�p� �?{��Mt�)�8�J��jɖ��^��7q��5l�ݒ�ˤ�g����c���/��I����)��=�ksh�ł-N�V�`�2���>+kC�N�Jn����ey�1xZ*3��\�����D����	�j�z;��Y������]����e�J�7��L�J	(	$���<�x(I�I�����V(�����o�������]'�(N-A����g~����o�#`>�K;�?�$���%����J��JԎ���N�2k����yK��`AasN�r0��4�*�1L)�|��U���.�Զ����`�9��p���JW��ǮU���\�1�R.a�^E�EV��ſ3���N?����)�0�K�N|�(��v�{��-q-#p*6����'Piԥ�������7��3X"1�@�\C�aȜZ�׆.��#s�d6�#�KX(U&QkL�?`WC����iQ��w1Y.��k?���p����:;�8�߽�:����1
�T�O)V�b�$���#Ƶ4��P)�P*���Y��P^����%x%coZs�tr������u�2,q�cQj�4D�a�wӅ�t� �*��d��?��	!Ť�}��礰������hwzR�ԙ9���T�$(�yyϼI�0�+Q)��n�"�o�p�`0���h�X�K���Nh��,f*�
�)F�/�d��ɮ;~Ga2Z����Q�8P.j�b�M>C�.�g�]�MV�}�3�o��W�{��}�-Dd���W~�g��݇��P�'����]�ԩn3\޾y�S��6e��9����	�J1�R��ֆ�N��I�H��J���7� �R	~�>>;^:2\[��ً���A��7ɟ�{�Y4x��}4��]j��.j����c׈�f:�hΣP*�4l}��HHE_L8
���'��%�y�4��~]��O��w��G��+/�L&I.�Y����
c��s�~����b�Q�����r���BF��U15a�Z��D�Q�OC7��vp�Q���[k����oq���~�M�[=���"-L��w���Nw$��sb#:����D�Ha� I|8EÀlz,3aE���@��QO\�I��}1ꚉ^��,]���.��b�F���W3�s,X����Iw�;�6��H��ʲ�9D Ac����d�&���!��B�$�4!���g��]СZ��J���<�JJ�<A_�8F]}v���B���(ׄJ�� ���0�/��`�$s�5s�	2<�$㘛h4�<��]&ߔ]&�tP,��gp���0�pϜ�ƞ�x�?���A�^e�-�lP��=�=�|�s`��"��1��6�:8s�ܶƤ���ʌ�I�j	�xvM�@�ݑ��wh�L١755��	��Tgp4�4eV�`�]K��@�trl��&h\�2 �s-�^��c9ֽ���\�)�>66����˒���(����8��a��s��s*~
|w�����BK=ɮ}Eib M��8c9�vmGhə?��rB~׀�0�`f9��_��w�A��&�@eav,�#��t,^Ƴ/Э|I������y�����&�	�t3����	A4��y�4�cvY�%�0�&�A2C?l�2�D��7W��0��(y�mNʸg�O�d:U;�중���#pe=C�n#��H��cJ�c��ј.$i�5�S2�=9���7�3���h !���D�FUT�\t��9����p��H�5�f�∊���|�R����sY#����=�UNS�v��m/�j�-��4�Ygg�6�̠C0x����O�PҞT�2��#��eW`PR;�}���ч�B��8��2g=X�$��`�Eյph�4��-|u�Sl��F��c����s�6���ꓳpK5�%qz��}�Hb�fBOԊy�W>�����6�|�nO|�1�|�D�!�C) ��cs��V$;uxIΝ?�[w�	;�K`Y��,����"[:)N~��G��2�40�O?�#���w�{�k$�H��܃�`��Q��t7/?F�U�,�����[����W�a{uMX(�
��=3�%�3��Oϣ�����T�Gڤ�"��?����w���~�������x��IdE^K��[�1:f�u��
�B���VW�r�:4g�}i�K�T��d�a�X���UZC��nO��L8/����{�~í����`n� ��xsK�t�(a K~���V���1v;�b"��r�׃�a�u	�����4�0.F������#�)�5q��Ӹ|�<��Pv�8�<f��q��g��W���J�H����\�B�F��0�,��p���%�m��-qh�	�!��r��E7t��C��4:`gec���vnA�����r������ţ����B�pY7�/�f�;A��
�Y��Ꝏt�	ʘ@בDA�А�-4	s��(FF�T9��R����F���^�/,y��+Ƒ A�>�i�p� Y�8$M��l��j��J�����V�&�gI�G&7d.��;����,A�OLa��m�,h��A���lS� A���
bENƗ�4N���D�c����fR���nU��N{�rE͙�.\v|��O���Q*����M(����9�������C����LI�po��(p~���b����4X����t��mIۚ����G���2�,0�����}���<�	���Х`��<�O�j�E��Cc.�DO���j�D*��gX�B@�)17e��`f��zU�c��rN#�.߁�r�;���|f'�4J��٦dw.��R7)GNa�ldp7Y�f��N�"����]�@� ��D���WC�H���d���	��4�B5�'2�$�� %���P`pq6���^���p��E�^�(�����$j̓����������E-C�*��<;g�Yx�����0��@J��)��9�#y��nG���||��G���ّ|!'�[�Vp��K�u�''�
����+ ��Г��B��Xr��m�6���MO��t�a��(Sa;�hڥ���	�k�B���	�w�,=�%��Q��7oހk["�mo��c��ٲ�IӐ�w�e�� ��uzvZȄ����%%ז�6�����0�����+�܏�G0��.et�tI��ڷ��{�����W��G�ڣw��B��{����̷~������ܑ�d�$���J7��'�8/#�4T�%��;TW%��z��'���'񑠌���|	咋N�G���c�JB@G��NZr�2jr���5Z蔗
�Ǝ��VKQWpfv���3����*�H�x�Ta��;"��rn(�����?�(�P�B��2޲CC2�sPT���r�/D�E� �x ��7
!�K�B�%ҍ�KG_��0��ȉ.�l6�2���'��[�B�`����~<��wp��1��0H��q���3iX���ט��T`g��-�t�+��B��L�����h9v��V.�t�3���U�V]SvO;Gg_��E��$x~Y�E�tbH(R�M�w�A���/�V��cr�R�ɜ�FM ���|�$>�y��̷I�Z����!�8%�������PA��TXRd�Z�>��d�Kd�l#���Lb�3�����e�Kp�g��7��:��ę_�����3�f��@�_L���Oaiu�_�UG�G1��3�P:�$�@�g0��c΋���q��I]sM��7G�$4�'Q@2�$F�T�e�:]�s��#e�I7� N�	�Y�]��|w4��Cr����n����>�����F��b���pA�:���Ρ�V�L�N�R?�n���\r��T�0.��#E#�:��\�%c"�#7C��;/;�-c�(%�$E��`���C'q#o�EUO�%�ͼ���`��n�G��˂,'������q�4�m�ZX:�#G�B������$���A��jq��z�,�G���R*"IC��t��Ɂ$ �5~0v&�2G�3ŝ@a¶9�n����%�H��gq���EfB
��g��]��C/�E��ϕ1P��\C�N=��,����<2��O�BI.������2J^zN�ka	��MI���~�.]M}2#&��<����P�T��F��T /�Q+c�Qw;o0 חK�K��v�C��1��V� {�c+����!����r?q<�d�B��7x��?�pm�]����^@V���J
"~O2�C�A��[�q�d��}0����S�-�9C��w�:8V^��,��j���
&�l�����o����>
f������\��Y��`������Skn�d5t�������
�7O���{]���my�,p��.؊�!��&(�6&U\x�#�|�����;yRd|6��d;��@΍�CI�N�D�lKqFs�[t#;v<X��H8tM�ba��`�`�6�b[�P�諅"F��x��}�h�hթ:
�$�y����$L>)jo��d-��I!*���r�qQ�bJ�@�����^�ք�:W�C�]�qvy��])�fL-~�(�.���u2���ी%8���,<lq�J�h���Q�e� ��+r�,�uS�f���	��d����	U.�7�xQ �M.�&P��v�����$M8Nty�h�CÄ�:vK%�&)�1	�D
-�ldҹ�ύ��Lgi��������tV�\�C�Ǟ{���{��{=d	�e9�e���Pʲq�"��NE�xd;���S���rCӭ@�Kb�BI���d�E�7�@�Ph�05
�hɮAwh���YL��h4d #N0��]��QZZ�B`�q��0�|.��b���R�f9��1'��
-%�����2����ؕ��M^�"�(I���L���Ȍ�/|}ض&�A��R�E�ZA�?��-��)��(����PV�`ʬo�F��͵��V��p�旸w�"� �^����Q���6��6ZH� �ł�;���U�;�;ńLI�&A c�0� `�^-I7���ϐz<�T���ÔI�`wc��󑳖�{c�N�x�d��g!�%�H�tJr�P������&(E%��&�t���fG@j�<�,�I��[��4C�?�=�*TY��}NS�{��ݸz���C�~ѵ#�S,Mf&�F��N.ʔ�,t����P)��	�TxV�~ ��1�$��ņ�V���G.�5��o�)����~������ϣ>È�ˁmZp4����vo$���Mg�W�+��r�-V��`��xFF�`���,�J$�i�taxʅ��0q$Rp)�M]|�$��)E9;�ҹNa�J%�2_��Lh|os�%D1���E*�N���<J�]v�c�y��^���8��
�g����m�L��T21ϑ"��a�.�{ �)vNLWH�p� ��3^i���|wU�a��J~�C,�ְ�z�?�.�;[H�#��?�cO����e���J��G�l>:��������c�+Ff#�l�t�0N�Q�;9����!\�q� )R�c�8u�e��wD/,�DeF���ɸ��k�w���2� M/p��9۔�Kv������w�H��,1�I+��n�lN��TR};�:�c�t�>���k�iQ���궬��`Β�M'�r��H��X ;��� ��A����|L�יM�{�M|���1�Y���i���hu2�?s`?�=u
�G����qv�?�ʡ;��qT��߱J�Y���J��.�|^�o*0(_qx��̲���r�����C�Y��U���n�,�#��:�t����sS���R|�b.4D`$	�Dv�Nj�*݀3���9�bj%î�uΪ���
q�4����rǥ*�@����A�wa�	&��QRV��%� ɩ�3=���=�nn��EW��X�sǡSr���vE�j�H��̠��A7�A;��%`����;��P*J�.\|�j801�G�=���ޔ��Fc��ə"w�C�?�!G��s�9�J�5��L0�;X�0��>GITH��-|vK��2J~2d�'�^d��n���7_#��ŕ����>���4:\P'pM�s%�c>x��9cB�5����Ю��ߜ]aP$H gq�\�H0(���>=�\[���}&���4�����    IDATy�AT��脑,1�� C[$�#�#`��g`c�!�()p5�Q,�X��,�97�Sm�Nf��B`^����f#�h{g~����0��3�����!+�X��0������P2�D�I@�&n����3p�,�򖘟��$#QNC�eXa2�@ gJ�(&�Ȣh�~��e����!��B����4����KDfL]��S�":x��h�-a��:\�n~ l�榇���FB��h0Xh�0�ZXZ�B��]�d��E���-2��5���F�.�dzcQ��й��$��,����\�3�-Q5�F2	�A4��x2)҄ٚR�
��������޼��w�ps3�L/a�|���D�d��y|D�2��B���s"dj�(�q�:0�QSA��P�s�3��I�����w�E!���\�˞I������d��N���3LE"k�L��XY��4/�n[0�MQ3-��0����M��� �]L�d��&G1A2��#�Ǝ9o=�|�b�b��D�C��T���DYH���ϧ���&��e�.�;���.�HV%�2�+ [/���,�|�%�w�A�#<t|Y����6z�^`Sꡒظ"�+��"��`A��/�K��|�\0���B9�(` �Eɔ;�y2�b��S�E@ș &S�A~ �Y� �o�l���'�;A��""����\�U ���X�I�p�\�&#A"�����"��YHv�h�����1O����H���~UlQ�R.11�om�����cI��v�*�y���,H8�Ƀʽ�Li�~y��#_��T�TsI4@>���&u�d5�`upK�[>�o��G�4���e.�F�q�Ι|�̪��=);������&�Z~���T���D��]XwJ�)ݖٙTI�(a4���$�d�,/f1�� ?�" H��;�Ē�1g�I ̾T��8��(ʈx^����ߗ��Д�w�b����dcyGA���;vPԾKA"i0h���+Q��
�=k�v2�-�4J�MޙH�h̠��>dh6�r�2���O��# ����oސNbcv��"����<�PG�X���:�%�$ϸNb�!�����_��ÁZ��܂r󤼗�o�}b���=�Le(&�pD�I���va��=��p6k<$$/���DDBLb�����8�/�t
�@�:�1=�X.77�e��J�3��e�J�(i�
�c7C��sU1�*��,3��X,�G�E[RT*58nqb����-O�t�HJ���Z�#�h������*�����)��6�0Bsa��Sh �;�S�D�:yo0Nr���}~6v_�,�5^W����)�
����(	5&E�������D>*������J��W��&'U�13��$�yO�}����u.��	?+]Ⱥ�D��FT�����KRx
P3&��9ӪB����Zr|r�!��(�<�e��m�'qQ�+Ǧ�u$b$"s�X9@2����26��䐒�F���w�����H�yJ/g���d��u���{�Iz��&��A�V�d���;��䄌��H�r9�)u�����M� >w���ǵ��*�u�q�ؠ�C��$�wy!\%C�*�I>�(U��*�
q#��ULc|�& O�D-�x��9�g���J`��`�Ȃ&|R��R-�ˠ� �/kqv����'	w�OI82�J�awo8��T��m��F��n��Ȉ�`#Y�a@��Y�=���	t�-P1��)]Ɉs�s�Dԃ���ACXF��Q0�F���b5���J������ꤨL�Amr�Ȑ��.pq0:�X�YȌ$g�
E��2���`�u��"�"�K���lª�9
|�!ePJV��%�)ʷ��������><���A��ak����d�i�� G B7H&T�eP�� }5�q�d$�.5�\�ꐵ��/���?�/W�:vC��`�Ԇ�����<MD��_�s+�*MĹ5�l@�\�����dS0�U�5��w҉bH-f��0�Se$�u���ߡ��dVǞ	?w�c"�=^<��T��)f�E�A2�,J���=�3�0�Aj�T��[X	���d!M*SK��Spl��ЃM�ȏLiIL��.��|��*��l+/��6q�)e�%'���I��)hݣ���F�[wv0�"�t˳�Onl�R~K���<u0�(.����@���T\�J��dv;/�;m�x��I��8�>�?�5a��OPB+t>S2��!�#?��#@�\$e�����_`g�k�6o�<=�����4L�<���#�CN�b�9�d�L�g7_�{U��Ʌ��ϑ� g>(�cW��{�UR�ɀ*����'^�"cX�)����5�.fT���AU ݘD x`F���J�+>��Y�t����l��6�{)����C�,�L��Ɍ���$X�� �]U�3�`s��t Ƴ%<�ҁ�,$9	�2|�0�M㙼���:+y2�:��\[@��@�z���ŋX_������ࡇ��S�W�_���ni�JyR��vZ%*Iz2�IL);9�Gn��I�X<�@�
�2�|�..�q��_������Λ������Ou#�dAm�Ƞ�tv3��ʓ�d��T�	��9贀��!�v�&�O�(=5�h�F�%�;��dlQ���#׊,P`��gT�Q��:�L��$�])���\0��݀�����+g	�"�B���R��q�XyJ�4n8�!����L��ܬt�s:�� 3E\��l}��`��p���é-`� W���V���'Ḛ�����]Z!#�x��ɴ"X�~�`��V�����:2+2���Q���:�#$l��V8���[�t0ċv��y����3d~�$�W-�(�c��WF��
R![�f�gbg����8QgW�)��
ԫb��R3Ű��,c�*���=�t�t����\�s�T�k2)KG4GR���`"�;4DR��j�}z�~�?���6�}�7�f���6Y5�|>gv�T��}��
�h<K�� ���a�%f4�)V?��$�~p��*��܏�K>C>!}�Ԓ�B-�2@�`Y���V��cg��0�)�Y��1bo������4����K�O�#OS���JA��Y�~ �:
�	�$)�B�#,����$�|�|>e*�.s���׶��D�n��-6d���*�Jq����̔�]&m��/���v��vzFӨ �ڔ�8⺬��{ӈ��,.u����,�9J$cq�����Dئ�T��j�I��I�ȡH��B���5�����n�zi����s�����_<���%T��*����xJF�Y�{(���4�wT�5���!�.���!cs�XWw�l���Qd-��$�ظ_'�1֫$�X���4x���8Ud�=�C��d\`C�w����	(sB�J�"���YõO���w���ۈ�����9�K�EGqr������9��t�a���L���Ɔ8�rLo4؅�BӸփs�%�r4�3��zd�dH�*䉒�2�J��,U������ۭ8�2K���P���۹�ݐ��[rߨ��W�d:͊� � m�b�4��>a}����4]�|��	
�N���zٌb)�8��G� y��w����a�Ej��u�;��s?�}T�[���<���ڨcfi��!3#�\"A{	�,@^����Bi��́s�$+�ɾ�}{����Sx��"/ƗW{�r}QZ�Fd�9��>�D��E��=���dy��A_� ���^����fP��.V�"��7��W2�,����C(SWsq�GGX%`�aIa^%C�.���	Y��8r%D�X�q� �umC$��S�8Jbspt�RQZ�d�Xqfm�Ι�!r���m���m�p��� ��(,t))'%),�ؕ�0�lL^�a��?A2(��0F���"�Ζ��ݯ�F��q�����3�"u�.�L�Wj,)���ő_c���s"sed6(�	g8h��Au�6)��"NY��2w��B�^.�&E�7-غ�������?
}֕w��E���0m���ya�{�.:�M�N��k�Q)�E�����[9������}�f�"��]B64�E�A�@����)	 �!�37�J�@�<�Tg� ����/�<��Q̛ȳe�s��xwDPQ�,��,򖖽P�4��g`�?�X�K���X�}��*�ݻ��Jh�.a{ǃiN _�Af��Gz���P��8�."��P6ɇ��^��D[w��._����g���L)\)YI�/�ו�Q����Ȯ��+(�vҘ�H������I���1QQ�EY�A�>�0vR]R$�����|���Ur�����g�;vE�'Zy%m���îSI!�r`(���3�ϱ#h���t�S�D���X�0�eJ�9�@iNL�l�|wo����
�UT�i��q7�\��6P,�#J(�S2b�i�/�e�ȅ�E��wPvml޻���7�(�lJ��0j3(כ0sE�%��8)���Q= ]:��sb�����i��yNXp�����ʞs�N��~wkIkժ#��Ѓ�Qo.�)7�0�k��,�I&E)(RA6�|��/�9,��*A�:_L���`�'"A1��TNC���Z��d�0Y�����8�(�x�$����lK�~/�;5,�݋j�!�����
�~�n^�L ���2��E�z9m,g$^w�!C�F��� �H9$�W��I)t�0ɒA��)�@�XaʭI,���3�����g�T�Z\��I���R�(BK��t)�kX�˳Ur6j��6�ɯqV�n��<���3���aQ*�m^�?����Wv�D��*W�sQ2���*�y�%���$�t*���2e��<�Y����C��ةSґQN"�"��%�+>?�O�'*�t����������}�����O.�,N�,�`���!FI����3�x�g�X~�WHڐ��mdQG )݁+sȗ��5|�����b��k�>I�_��I���� ��EЌIW��P���Mb��N��.F�[�G] ���5��O@��E��B�J���*N�4�@�X�:�� ��Vy_͇��EC�qG��Hj$Ђ>��:[H�9��sE��y�'��9��K�'c0(�3�f�Ǯ	��,���Ӎ��u������Nn��؀q�yZIY��K�-�u��q�y��&|�vW0�]C�m�xrp�H����cY�*�';τHx�G $�)�G䒬�dǡB�J��cI��^��1��w;r���4��9�������T'W^?!���I�"c ��lv�#Ƴ5����?�)�'�,�xl�QZH���?Der� �LlnvD�J�����抉�dJE��z���a�����c�l�S{���Ž���F�t��Tk�h� _*#�2$�҄��Sf$w�5	�G���z�-��ٹ�NgE�L�B�:�Ry�]1>��wʏG:Ƴrv՘�}�J-J<�c���6��C�s�%(���Ckc}�A2yG�Y��G�8I����X��8��;an�T�U�%�5�����X��d�Wc���)��2�&��uv71�nϑ�k��,bzvQ���?4M���3I@�Vކaȹ��g1=?���#3��$��:����0�.-����w�e!�w��8�[��P&�5q������J�y	F1��(-d׎KG=�J9NʼR�#���C�#�ʋ�2�N^��Rc�U�f�N��EK]qX�J���S����� QzQtF���l�k�ଆT��&27� <�ߙ̨���^@�X	 xD��@�5Y�9N4&%���2H�U �!����#c��!�(2.�L|�ߦ"�bC��4�����ӄ�	�3:��L+{�U`���z�7oC�]{�?�t�Fa�K[��(��8

;�l����EB��QvmhEL`Ď�8V�妬����:F��d�)?M?;�1����?�؞l�(�LJA(���B�l2;H]��!�7h�Yve���`baaj�Y$����HM�	BBV� ]�*�V��u�Z�J�Ѓ],�sܫ���Jז3	���,���n6��z���3;�Ľq��#r���zc��Cr4#�%H��2��`�?֌�/�`�@�����M�2$����4#�Z$�[�������+�*�Ȍ}���<��*
n"��Օ����}��<gAi=Qd	'�(Q�E�S
�*�qU�hHz�Y��c6$�[n�S���c?�B�0X"M�;���K,�1���RRǊ�{����t�1����G'2�M��.փ@���DB��A�5�{&s�D[!.������lb���iy�I���E�R��HbN�V�l�H/�y+�ώ�OF�D��j-D�6���T�?ӡ���h����H09��B��@]8��+Qoa��E�Q%u�:�
OF�>ƽ,�=z� ��d&4'��{	��,����]�.�Ri=4�m�h�z�����+-��7��G�p~r�z��XM��۵�����ذ�$���xn�4���x��>z�?�G�.��+��ou�0�c��$�M��ey����f��J�E�|�*��0�w6�V��/
(�gN�ǽ��p��STkԔO,�!�a��u$�f+:�R�M s-Y�fQO4uY�dW�,�b;�y?Y$i���i"��Ok��a�O>�r�C�qڹƌل^�+o��}k/�.I���
Ɏ�tmn�4� e��!�[4��5��Ϩ��~��}�c�7��Cd�+8yX�u��D�|=�z�V��C1 	�Rh�q�b4`TLWS�v��Q]��k���T���M�]=���Z�n?_&Q���[å��oQ6y_I!��;0��lj�O�YS�U��e5�7��S�87e�pEXT56�0M��)�T��j���Ұ���	�����F*t)����	f�s]'��k�mĕ��r=�\<_�<�%a��%F�
��7n]�r1£/>�;7vQ)���?�=�#n�"m_G־�Ɇ�xf�F�����,����!��4��ZMZ���1z����_��� ��U��� ~��AN�I�gqȢ�{�9&���5��;M�m��+&P�{6a�,rL�^"�@����L�/�mr%�E��w�ڿ�z��r��ft(4��{"e�i�`�Ԋg�����������j����L��Q�9u�?���)�q�X"�_�խػ�&4�C�bS�3�9�!m� ;a9�0�ji$P�����1���=�͒"��ijB`�4f�Li��nG�%!5���G��Q����o������F)n(.EuG�t�ik����r�뀫�A$]����W�����	�Nq��>c9;��qP�>Dm�M,��M�8�d�4��D)����F�FZ4������Z�3�}�����x%�S_��>�x�唱/�7���7~ө�/{��3y����0e[��
�`9z��o0<���)ܞ��i�}햼C�q5��*��"3��S�ql��aE�~ͺ��
�Ȉm�}�����b(<�;W�ھ� �9C�ƚ/�UXkhm96�X�N�5�v���˭5��a:W�!�F��d���cN���5�URxq��ۢ��$�Ӱ�$&b�8f�~OAc�g��l>���ث�^YB��$�ߗOǨWCԫ�Gxz��u_h�Q�E�Bvp�Wo�Zki2H����"�l�%����v���h�ƺx��� �A�?���7�AL������K���7�����G��?������_�Ϳ������w~����.�F�r�ᛣ^�('G�l�}�0]���-�gX���,'��ѕ�Vk"W�t&�(fJ��f��\Y�Z 6�;RH����"ڵ�:tx��VBN78���>�&�y%�a=�z1� �(F9L���~JzO��<T��S�E�5�½�G��/��3�B����F;�׶�E��qJ�.ue��6SM٨��-38�.��,f�kQ�4�`��*��k%��#T�!�����/O�*n}�k�r��I]E�(g���:ͫ#�8�,'�8L8���6c�����T�-��<D�����䖤npjˢ�F��(��x���Q
tĊ:ŏ�DH�	a�m�'y]#f3q���F×����G)�{�h6����X��J�]�3���    IDAT�A�	P�DA�d�';
�,��4�I��\#���Ta�[�Β��55����]{W�C��	�Ii}K4B҂�I��F�Q�?g3O��U��V���/��Ӯ`k+C��峧 @�8��s��:��.V^&]�()�g���D�8IA�IIzqv�|��{3�jc�jmTZ��:f˒@T���ڇ�	o�3�۵R����,�4!�]������Z)ӳ��b��>V�^3��x��*�mY�r�)������%�'��rl�m9�����Ƣ�qX$��6��jd��̪񪧽cLOc3>�6	Y��|:��҆�?n���Қ���F�U5����!0vxx��
'�/�eԳL�������Ŏh��MAԤǝ�A)<8�ѵ2گ�y�j����8?~��ǟ����^.�۲����f0��X��Y��M����S����b[Қٟk�#3�騻dA�2�D�[��$
�����N��x�>�D��I��\C�5E���Nߕ�d�UM��d�
�Y��d	=�k`� ��h���NP��lJ���� O���щ"5�~�ZZ�E����-�m:��Y�ji�@缥1;�䣵��k�^<�
�ﾏg|O�{{�*��\�c��:�Ӎ11�s!��
�-֊�(���3,z�5Y�|`���uD�=��:JQ��fK|�����*���cdN�|�W
��9X��*b�j`�5ff��{˾��^#�G]lf]�����:j&��/K���b�`ق��-a�w� U�Z��F;�;���A`ZXNLh��xt���%��>J��X3q� ��U�6��<{�l�!��csE���c�]e1�z�t:\�<�~;�79�w���b���j���h���lS�| "��MaIs搢�s�Й�V��}|��1�/��<���˵q�� ڹ���5Q��3��XF5��-���9�zH�.�k�{�f�-�AlIK�9'�����S��]���^�~�{W�u���ULl�7�zq�F��?��Q���. ��()k6���!kU�5����S^�x��ӡ6.�xv�'�_H�d�U����쿁�k�?��C �̶4�y�~�?�����7�kH�ɽ�QZ�Q��'���I��5u���q/�ā ]K�lFf)c;ʹ�/~�ϥ��\NH2Tvo�q��Y�=�G!t͠zN�Qt�no�u�Psa��I�/�.���s������9�_�p#�P߹��)�v�Y�I����W�PX�2��&�ڍ�vKS0*6�r�	rT&��F���S��Sl�3 �!ؾ���_�j]A@�"�F��� fSM M^D5�f0��h7Ct�>���3,N�g`
���Ƅ���A�����@Bƚq��b& �-ʩ�����Js�:3b�c���1��O���)z�y�a���w��v�p�TP��DGtt9²'0���V��Q����t6-����ˆ=��
���p���j�e>��r���ns�6������5˪�x�x#d�IOX_k�[T�^OD-5>Ѭ
ŝ�~�n$���g?�飏�� ��!ܹ���ME1w�T�x%P�:��w�y)G��px��&����`yI���5��f������P���Ϩa`e�Q���*�����������f�����_bSj�����!��^9VS�PUYs�J6]��s�!|��� �&a9<�z>��)j��,ys��p6��o�b鋅_��5ֲI�f��y{�Ĕ�z �AQ��6a�tx\0��� b�٨�դ�̹0�a͠�5.��F	�Ȑf��R�\��\ͩ�|@�PF�����Nv,���/�!"N<$�8E>�rt��|lԻ D����(�,�]!U�\�"����9/-��B�*N�<ļ7P�J��:��}����a3���[6A��q�� �E�墢�.�մo�ZRi�*J
��a)��QH+h1MJQ��:��
�\Ȣ����-�� 4n�=�\w� |��05���#,�G��_b�����NJ:�l2��']N& |X萾�&�>C���Y���q�7���A��c�D�%��&)b�����S�Ӿ	h�X͍�����9%�1�s�儉S4Z��d�K�Uqx톄���	��[[!�������«7Qm�`�ɰ�Mo�9�u5̨u:���~��,��鞼��z�T�α^�Q�2T;��;Xztx�D�������B�������ɀ�M7�3�$�!d��X��$��Eyi�G�����(��i�������kן��57��������l��$՗������t��!�:GٌX�S�����:�?���16������^sAc~�Ҥ��N����䁣,/�e�*ob]��=?E��&,&����?�b8D�Y��:¤�)5Qι�pIGS�^�{g�$
�U�b:����},'@>r:����D1i"���fd)���Ҵ�����Y�8�z�e�/3�kr�ʵ�k��pҔ� B5I�����=G��P��g�>��r\��+����O�2��Yj*A���3���'t�nЮ�#і	��Hխ$1�Mf|��Ž0�?VS��q����d�a��Ԁ�x.��]�9]RA�aB#4҇���W�}p��xگoW=<��#�UZYcY�*&%j#��61�mj�?&r��#�h�CY����|���C��7c�dB�Ҿ����4Â�>	h���=�lW����Ӧ0�GO|GmS�x���qj�f�!�QH���gȻ/�$35�̡d�o���ZkG�S��q����g�3F�6�g�i�I��F����{��h"'Z��\6�,)K�n0����||l9���|Bx�]t���Kv����i)� 5����^�����Im�&x�Koao����T�F/���o�+����2���{�M�*DLp���؁�DI:6��lX���\N�������>��sLG#�+אm��Fg~X8�I8)�b2q���>�vc���gS^"Z��9�`�hp2ȵ�J��p��̐�8?ǬO���Q_b�h�*Z{W9�ƌ9~kOg��LN�lL-+Z8�L�F���'��'�>�3�N2)x�
�r�G����K�(�!J~������[hn��`DV�B�|j�b��h��m��gͷ�������~��1M8i��1�.P�� d#j@e�zI:q�q�H��Q��b�g�Y<�b#���5Q;x����	�r������P4Bi͊���W^ip�S�\�BD� ����@���<{�3�l1%�/���wս/cQz�r?��[@��ԌK�`Ӥ�P�k�ו��L���B�ȱ.��LӴ��	&�#N�@>:B)�[�\n��?�
�h�	�*��)<AN��ߓv,��Y3��v�/>�6&O>��wfg)܍���0[���V����\�[��X{Xp�-'24�d��Y3�QKBT�.�������a�� j �\Gc�ٮ h�k����A6��Y\���p��b8��^��܁����w��HJ�=��'w����ʟ�w:h^��J��R�k;>�\�Á�N�ܴ�:^�U3�2wrS7��� �wx�+QY�`��<��'�_<�9'� ��W~��U$Y]C+��Q#o�[z���%r/���}�|��̱.�]�)'��L�/6���b�f���6sEA�pӈ�Ф�Q�~��&�ÿ�������?��wp~t�����W�һ_������~rImK:���"X���9n3bIB�L��X'،��m��b���
�ѭi���޴$���y��~����S�u��1h�@Z4/���3�'�>��c�c�!�(���)WP
I_˰��-	" 
5͛hh���T9���d�L �#�hOlu���nG"X�}v�h��9���6s�^�a�0k"L��ot/����)tN�|h���&���},�s�����2\�V�vQ���R8�tE������U�݈�� f�TV��h�Tf5��LY�3Z���pj(E<�� G���� �"�n�$����6K�D�h�j�}4��ĸ˜�#�Kqʃ��� ��-�Q���� 5'�Q�Ǽ'6�4b��T�+�+'�2�d�1h����Mp�q�:��$���$H�9z�O�}�@���n��"��P�� �Xұ���*�5��Ҝ9�`�������j���p �\�������]���9C��([��F��lf�����SHCk�Sm�t��c�=�����XN�Z�qs������� s�xs�+(�]R��O��l�x��9�!��Ź7a4�3�a<��)%-�1��������TV~�f����P��#�uП�4�T
s13��N�x��^9_�4�eV���9b1Jj�4��n(jm��d�cx~���ʛ	�2Q�\:g��F��CT� /���޿�.s���V+��T����u�}�k������¬w�����N�5�8o:/���lC�j�ic����x����DJ�߄uD�=T;Ê�g��g:I"�V|��$%���׉�1�k�
�U��pE�>�T2R�-猀����'�ax����Xmb��-�Q�u�;M�cV�1�!��nP^�j⥛p4D����f�w����k�f~�$��у�1꿔�A�`TA�u���M��fR�g��_��A~&�!�FV�
eT�[�\�"ӌF-���!���	f_|�'YIi�*J��6��S](͍��)K/c�e�ծI_���]���>��	fSDW�m�Bg�*�t�>�$�#����q���!|�(_��^Z&)BH`HxH�t6�4C�qY:N�9	�ז�'�r�^#Bm���7�uL�k\�v����=�t%��d��t�*pxv8퍛����N	�qbROy�A���Pϧ�L�@u;�o!��'[A&P��ᱢ���Y\^�\�P�j��[w�j��<@��������%����:7Qߺ��{q$�3<Y���ڙ���:-�/=����]l�����x;t&����}�Sy���;gl�\Z�%�\f��dj`��6�q��dLfN"�:���ܮ��L`�{X�w�ͤV���0Fu�
���0�,mR�L��z�`'�k�2n/p�.��8C����;7jJ��Zu�<��'���fC�^#�w�١~i+P����C�/��&&�T�p�5��3l��p�'* �����8m�y�.�<"%�ِecȌ����-��w��Ά�8}�	��lfC�am�� j��4�t��	�hM!p�MU�kbl�G�4ro���7��leleTq�X޴[)NO��ɇXNO�ݏ~I;�o�o���m�&������������o���=�x<�*�4�]�.��Ƣ��A�O0:���`�{j� ���u�;�=x���D�NַS,�C�Xu9��t^�J��������{�6�l;��J�+�d��������6����'��d�qߍ�&��@����Ѫ��J9����>�����4�~#��
Щt��&hj����u_l:h����ObF���������m�.Ƅ��8L���)��C�ѧX�α�W� ��:�7P�	�&ج���ɠ��b�5��F�w�}���p�͠����yv8}lP�t��=�/>�)V�����C�m���˿�M��`ͤg��(0���4��͜�D���q��FS��������&�d��.*���d3��o��R��m�CC�#L������O��o��~���w��ؿ����_�*�������M,�q��z�R�i�Vh5uX��0�Gz�P8<ﾔ�(5q\�Is�	D��f�ਘ,����`P���f-k^��x�vD|QB��)����Ο}�U�\S�Ph"��"�la]�1�̓�&�OA)p:��ɸsrc)W9iJ��9�G���F8k�'����FFғ�mčmQ��VdSO������KYg	5���/���qӄ1ԴJ��2ۓ�����Vިv�Q�Ҥ�D	蝜ؽ���J���6��6��ε���u��=�v'������P�$�%R�Ak�%m�CP�U������R�{�>���C3
#e"蠵���ńg��t�8��/�g��f���^9���tBz��4�G�l�D�5�7�p��S�6cx�2ބ�;�5P�N���Y��7���i��Uf�]�=m�I�Vg~��/>ó��e�%���ؔ��%��I�x��l�ئ�6H��fU�����G�c�� �*�QF)잭X��^<(Iev�N�K��6�g*��4��/'˼�!�4�b�d���f��{?Ĝ�-�v��(EUQ`k�L4�"��@R����D+!�df)�;���=LG����ut�UA�b�Y��f��#̏)����j6�+�i��o�&]o:��Sm�F��~��u�]���ց\���[�.�|�O��G�m�����>�nyA���Ю�,���d���U��j�]M��{89y���c�Vi�P���(�\�z]f�O���2��A�e8��S��q/l 9��HF����Lr�������<�cԫ5e�~q�gOz�ҫ�;�R�/�O�y'��vE1�m�Cڧ(Qu�]�M*����D����Pw(9ʚm;��k{�>ΦcM��ϻ���Y�M'h
�PhI�?���+����e��B���^��>8@gg�F�F�O?�>{�;X���(gWt�c/��M9����(`!.�[%f��%�Eǟ���9@v�dԮ"i���CB�oE��E��qҡ�"�Y+\d*#*&K3��	����X4b8�))�Ҩ��1]��pq�#�J�׋�l��(3����5z���B��Mctk�tX���7�k�:�SN�(��"Ӏ��^>&�S�'2g�}YM�،g�[ؽ~崆���4���0Ej�yP�L6n�I���-��61����-��ޏ��g?@~q�ru��7�h�p�W�)i���/�S���\'�l�l�*�z�#�x��ݧ@0�Wi���Ja�O�9k�'�|c��2V9c�]ar���(cњo���ɽ���l
�g�8�9V��� �]M�P�S�s�o�NE��S�>\Ql�W*K�i�C�L�}ӢG8M���O�˫�~Z�����\cԿ���5�h4�Q�~�uSgs'�������+Av�O����si�Y'z�����5x�%O�?�Z�6  �c�EAyT�	��������Gw����ƪy�k���b�1��N�	��az3�k:Wd��f:
tA��=S�.�O�$�E�	�T+e��/p��s,/���h6���w0���H�1���X�R�q����:�&ڄ`�q�14"tl>O��1<�]�ت'���/�@��'ȇ/P�a\A����W��V4	�k/���w3A��,S�/s�%���`'�����>�)֣��:�6Z�[���h�#_D�ڽ����2��L�������g�F=A�付?��DW�-��W�4QJ���R��nz]PDE��Ym��>lQ]�!�3tTM�I�Jbdi��[���1�w?P#��H[d�&j�L'��iHh�撴闘Y+=��:]�Aw.9�.����̐l�I6�v����gx����N4�jn�`���[r4g�8�W�N���=�g�SR�����oU��/�����zc�]t5,�!� �����9A=�
}�����n�!1)G�ʤC�֢�5j�������7���� a9Ɲ��V��ӏ���޷��Ь_���]D���N6s(��ؔШ�Wt_<���2aعss-%M��6��a�A
X�~�F�H�K��U�W4f|���_�j�Oh�@�hY�]OѪG8?}���O��fX�8�c8TQ� 1/�:C~�<�I��P�<)g@��,<3G��t6��t�5J��]���,�?���{J�����N��=�6�<�tm���īnL�Bp5E1O��
���,𳴆,�c:a�i�Dt0WMl�X�H��1�J��
x��:~��S.X~����JsWN{�	]ǌ*��0��X
*Q�W���@Z�V�3|�F �̱�� �b��
Y���,���8y��RR��칰����jX���fQ��zbS�IB&{�/>H� -�W�����P��v+�b���� l��Hz"j*�=E�c�<)q�>.T`k*��,�Ӹ�V{GY���*�����O��Y��    IDATg����&�*��
J%R�@)t(�0g���sA���[m�]���09~���\�,eVjH���:�^��
�sZ�T%�~�ާS��hf"�(��,���/�)	'm�Q4�W�^A-�0>}���3���+M@s��>��+�ʶI��bcCCR���"*\ ,Zev��'eU:4��w�MD��4���.F�.�>ǂ��#H�M2T������֨Y.$�<`�%%�P�������uEӹ9Z����އ��tr?Ko퉎;g���Ӊ���r4B-")����U^��|��d9�ы����\ˬ`W�	��8��hKa�"��Ōh6W�Y,��t��ϋ!'Np�2����SNx�.���"՚�ӛ�T�bi���ǒ"�<>O�<s��B����Z��̣�Uh���Qf^h4����B�&�}�_\���a2� c��z��j5�<%R�YlQ��k!�t�<�����t_"./����x�H=����o~��y���6(�*J�܊���fX�YX#K��p����2�����j�FPfqL����!j�����M��h�B�q<��ڴ�����,���J�˦_,�+������j�m������}����)���Жe'�#]����R����_�~�"��� �@3
�;��g/�8;�fc� Bm�nwW����ܐ~ �k��:i�������6��_��흚����
���{8��}�f�:W��t����.U���Dr��I��̆�)��w�,�٨�ݨ ��t6<��f/̐U����7��:9���it
�-I^��CZ媲aC�&�5��@�3iS{��笒����ZR������&u�e�s:A�aPQCk���ԇFM����&8@�.0�83.%TZb2
��0���x��Ob���Z��l,�Z]�~j#�&7�L^�ޜ�A�xt�*!�t���t������
!JS$���M����|�u�L�A�,�.E|Q��:��J��l���K����}���DIc66�(Lb�
JU�j�M�,�G�� � +RF�e���w4�S/���ܺ�|�A���6�Fk�j�r��
ȵ���i��via8��铇XR����h Ӕ��Ќ�XQ^�i�����6�h��'����D����ݫ(7n"�k��)�@�<�@`Mjp�ȇ�K���һo�p7��_'f�C�� @u�:������9f� W�T#�]'���*�����a�s~���٩�飻�<Ś�n%�����U"S7������1=��H��)7�.���:ТF����;�_���_3���n��|�����-ܥj��ޖSL�Ew956��s	-����~w�*�U-&��9�qcwwQ���8?:��+��i#�6̀NM���� Δ�G`d�m%�՛��z�*����x��b�U�P�G1�8Vi�spP2o�h�C����o7s)���1�
�!��Ϟ㫿�K���/�`w����.�NGh7p���޿� �WV��=�Zlײ8aA��j�F�E�����c\�x��|du9c�J��8Re��w� ��_,"^U��
5ӂW��W��(Y�!q/Q�F�j���Oq���
n���˯���؂�A3F����/�ݵzZ���\�Ú���� #q��f�b��˳��0���s�z]iuǕ�^E�����V��i��Ni���uDϰA��\�>H�z���"�$'��#N�p���&�x�IW�N���s�f�f@��!jl�枆�]"��J�J�n����}p�.���M��2TT��Q �%���0���)�Ϗe��Zl�Uv��^P�4�ڄ\�r3�:�֔�ץpܞ�B/��K���W����~���f��/���u����%�BrI[B6k�&}Nؖ�LO8�a֢�y�F�)�6�:��>j���U�<���?��� ׮��h��Rj�@����F��b��rP�V�h�E�\�`p�+�G�
gRҡ�JM�Z�V�����1��4��ݻ5�r��h�Y[y}l-�������4�W��.�=�b:�-��gMlʉ��h:R�l.k�r%��֍���
+@��7��kk_5�9v�w���^k�=�3d��.�1��a�� � ��E�럫����.v��D�ZAZ&Yf���������	��}�;װ$J�'��Z�lϚ��I��rz&�)�(�%t��|&}	��&˹;C6��,I�!�1�mr̿+33�i/i��N�9�������Z�.ٚ|�Q�ɸ��``�.N�U]����I��\���Nu
�R���d�y��x�6��9�&��f���'$���é]�= � ��Q����q"��A�a���߹�	���\�sLN�썠i����U�(�1�e5���RM��l��tɋ��F:��$�Y2���Ɠ���v���a�">'�� '�4%0�9���J/�拔0^k��r��fP8�������G��x�"�4D�SG�����G���p����Vka�ZP=�x�����<3�l�=y��h��� �.�����V�&�׽�Q5b��9�Ϗ��D�LT[t7N1��R[�����4,L��1�Ԗ1�)I�֛w���B��V����_��b5�H#��y�eko�r]�M�� ����H��+�A��X-+F�Z����h�6��0Y�2>��}�}֊A���>��=��"[�M���P��	�Qh�����Xc�\�����{��rp�V����?�d4T�?ؼ�B�4I\��&^Jj��<��p�F�1�b˩�ъfil�d�5�� 6��J�uEЀ��6ҐŁr\�橢gSŪӻʌ���=>5m�cL�aú�"嬊��xa�:ƚQU4lN��t@�^�#Dӧ������e�ө��g����٢��R4I�@(u]�f��{�w M�8��=�N�]d�V&���x�I�4A�|��VK��/&�����#F�);��E[5�u%�� ��y*cJ��4�9��
���t�rGw�m�Yŵ���U#\��������z����>zS:·f&�n�7r	7:�0���@�J��Z���w���v������I��Q��̯ak���s,�!v�n)s�J��*���a*&2�x�q�K�x���b�pG.����\s4M�b�1΁Q^�ңk�q��(�AI�L�,{�WXqQz�(a�-�VۘT��H>`W�^Q�t~������%B�y%��8�p��S����NSu�jݫq@� t�[���v�a.�	�Z[;[��ٕ�`0�h440�u:�}�kxC�+��2�\됆�%tv�ppuY5S��1:��#f1SB)ב�(AژqC^�h~�f���V��9Q�ʥ5�8}�L��wn^G�^�|2��O?�h0��_B�T��/^b8`Vg !��6�F;��Ȫh$e�9�i�>#W�hT���x��`����g#�Zhw���C�u����x�8��$�ѩ�]k�����xFLS/C9i#L��2�𤧰p+P6Cc�I2��O�R�N5�����+q��2SC�.t�,e��w�����5�[{H�ML��׬�9%4g9stZ��bQ�F�!��DE?5i��L�.�YW�w1�{fS�Ų�J�z�z5C�^�ax��ِ.���*�-�A��#�١�޻�E&ݓ���U�W���e�i
9�*�f�@N~��A�UE��N�8;=��b$m'�i�#1�1-�d9 �N�WӾ��̞q�C�T��3Dt����f=EXf�)zD���+M�q�ϦT>�2'Q訬�\M��-����C4u���]#�<���pz� �?~���;W�ȫX���YXw���fK�e��	�j�	~��TS��Hȣ�HM��X0�s���6n{�`P���s;<5�պ2ĒNj��f��1��
µ��kT#�����T�� Q?>RA��3R4�	�����!m�;_�y% w��k��UW��T0"���g'�ZW�ʚ��1��r5F/!�.lӜ�d��lM_Ԧ+ׯ�֨`3�a3?ÓO��g��{����=\y��2������Ȍ��D�c���J�x sa5���|)��)�t��*�IӋ�*��5�w�R@3�"��4�����Z#8;�)�F�M�M�Ht�4�I���ez��g�/�����;��,lG��&��h�\ŏ�>�ψQ�l/�A*��4�%�ے�8����7n��c6+�\��c6�g!�S��������ѳg8����R�8I �?t��q����S,���Y��|�dkw��U��	NFeD�=���e5���jS�|f˗וT��i�!�y���0Q'�I?�B���n;~Q�:ˈ�k��v#S�̌"���w.%R��N�bu^�Qm�P��5��?;�|<S3p���y��Vt_4�R�i�d/�N����B��k�o����KΝ��H��A�6#�f��
��R��1�LjJ�}�\F�V�\���LE	��"�d���V�:'�g�l�8y~��?SPtu�*�;w��X�Z(��(�&�DIY�$�jl�Q��!擅�m3W׌�	f,T�5�e� ����2�u���PX����5��?|ټY#�,G3
Z���f����5���H��jq���M��M-���/�n��<�in�:E�*3kQ��k�rm+OY��5:�O3���+�ʤ(������N�?N$�g���e�57NkN�ɔ�n�M$z�ٸ����)�(1��R�u�!e���l?�D��l^f��!�ג@�i̤�:K�pt6�Sf.I��+j�i@�*
P|U�YR���sOE���+�x!��5.�)g�Ǻ���G�D�9���a�cE�[n:�MR��������"�I4[WP�#�^���*o�9���"�a!��(#x*��@�s��SK-2i�t\ԉ�k���&[��#��2řM�:�6��_���\���A�����+�F�]xmS5�aTXF`��;N��_�X�[�ʽ���FRM�o2�[�R�i⪤s��p�$+��BWc;�B�	��%+�WZ�+�i�����`�z���ȕ��Z-];�.�@�g�i7�tUt���2&c�o�:��r������zT���M\��a��U��N��S��L��g1s���Fܫ���(�p��u�'}��]���56�h�؏�G�$�^���)����f� �fũ���t���	œor1�fn��e��
j�6��p��W��ز�1�$���qm1���jTF-�Q^�0Т���Tyct,�u����q<`���8/.ۍ��t^��4��^�=
<��j�=�W� ��yxcL��B8"/y)���(m�C_���^8�4��i�ԁ[2�B���K��f�����Ht��.3\�+l0������~��6a���@�&'<�E�� ;@C:�2gz:}�P�*������ a�a&Ѳ�f��X����9x�.Zf�"Z�R`�L����l��h�/� N�JI�_"�̅#���`��`A
��T��^M*lJa�5-*NԨ�A���6�(�e�cJ� �tBqomU(�5/��`]_6y�7w���k�u`��X�v0ҍ*G%��hVP.�1�1�1��1X��(�M����+�*!R\���5���*q������O`���5"̧=LN���I7�R�M��ڐ%74E�k���Fe�È�E��D�(�d�{JTW~�?�2�щ�hM��8Z�E��X\'�>kJQ皹ƫF��os����J�{��B�8�驙2�N7�q��,P�y�3�ԙ(9M��ݢth̫&P�S�EVc����j����x��pl:~��*9o���BKK+����P	%N��Vo��6��j��~���'�^�Q߿����h_�%�t��1�K���2���zLK>��n���6�D��0_p�#�L�Y��hi1��M����=�!�r�u�e����E��=Vę̡�e#o���22�w�l�̔I@���T��<��ҵО�.v|��>K�LXk�e��HM�����U�h洂��h
IGd�Z���)�䤧�Rl'��WFeL&#���O>~���������fh^Û������1V�]�!D�r{J%ڃج��*f+^��5������z�%u)	�s,鞪<Uj،�k4C��F�� +af�&��J+�e��T�e���'����$@�`1����f��b�@�4�;S������ ��1t�4�^�J���w�	إ����מCm�|i�h��Ob�3:R����u,��\X�N��%Я��)��:D��D�3#'��|�f+/���O��ը���!�;��X,*�@`�,�}�ܾsC������HY�=��3��-�31L6�ǣ�)ʔ���!�j*��WX8���p,�H+��5֌T���A�����szj����#!s��c8����	������/dT�'�1��++�kH����{A�����`�	����bSRhmS:b�(�1��Z�'?�0(�@e�0]ؚ�>`�z�����X�Ǣu��d#IGy?`F���h���`�z2X���܍C�&c$�Wn�Dg�Ҋf�	&�<
��S�)���&��3���}������p���P%�E��L�ʀ�-��%<�'�4��O�>��.RJc�bc�7X��S�lM6�y��AƇ�����a��=��I�:&ɂ�Լ��Dl��@.^�2u���d.�&[�	y�Q@�f��i��N���	��	��8��V�����wp��[8z~��OO0-�$��Ľ���������$Q��˽�j&��:���I���-Yq3�,�\cw����U���D^EJM��mQt�4� ֔��%�ӱ�D�����S�����A1[J.��E� �{0�l����~�0w3sٱ�^U&�ЪNM�_ɪ��C&1��2���YI���d�h�	�f������xJW��JfQN�%�����/���{(��Qz�w�k5��OF|�"3����^���/tI��X�t�D���vs���qѥ#�e����Z��Aҝ<Yl��NB�^rs�!�d1ǔ!]��X���K�.���*֋)MQ�;gN�k�h3J������7�r�ip8��i�Zt�*����*�!�enN�С�&Qe�<.����B���� ��C��I�<N ��h"B�'�}�����<��sv2w.�| �dF�>�vU�0�Q
�h��*L[�k�6mXx�Y��$.ݳ�ah�Pfڐ�Ĺ��WB��D9�`�Ȣ����T<�0ddbQ�j��oW�JWQL)��l kr٘�T��!_���Y���ҖdqU����t����v�IOq�0p���0W�!�+���+��2�������hr+Tj��ZF�h8��@��h�ET�v��Sd{�����^#�_hd��6ڭ�x�)�^>�n)N��S�{H�Xp*Xb�:Ԭ]L�FNp�B=�X44tr�X��(�u�z9k=s[��G��p���!�:MMo�ы��k��E
��8��t͠� ��O�>�(/�*�`��C��N3�a��K�	G�*�!�Q��7D�[1�w�Ģ�W�OH7��r�e�Q�Մ��SD1�y�D�!͗����ӡ�Q�4��tE�����*�{�6����?���!@mV���;_�;��X�8/qp�F�`�!�>��?l���I�Æ�]R�9cl����b�+�á��^F{*�S��ɀ':��-�@���w����n5	�)�5:�L��⒚�����,��TEj�x�Y\R[��
j{M��s������*�ka��*s��4<��0��|6��<힉F.��OT9������t<�H�#�l��H��͟l��	|5J�z���^�_����g��k��/��}��2�)#���ͯ��ߒ�9��h�S�U��r?�԰0|>��2�"�(��Q�cԝ"X32(CĽD�i�6�H��j�"0iX��A�DU�dߞ�\�x�*�j�K�c��1g��j�J�a�/��IQ,��L�s�u6i�I86<+:[�hM�\�إ���4Cѩ.�Jc��p����L����؄q�`S����a4�����4�H:���	̭�    IDAT����UT�T�0tPf�d�����#������Ǩn�`{��cF.�Т�1Mc������w���HU@�OmZA��d�����y�q���p�P��6��,�R���^A�v.h�#�.����y��  @߿-	����c��`2f���}.�4C}�U�RN���aT鷌ע�u�s���Mj������<,��(`ǰ<6������
K�t�O�2�
ng)�.�5u�Ǖ�A��-UL��������Rg��[#eLf	c����C|��GM���׏��\�}������C�y��@l_�9�;�W��p��y�L�%���2q��2��2����~�򓍹����P�²	(�;�s�giK�C�`9S��M^0b��[��|�=Нw�wI_,s��(V�p{U�zƼ����lb3(9��.��a>�J�6�|�l�
W�D5�M#,��U�c_�y�u!�Hj�`00����7E���8Ť؎��:ۇ��"<y�ǣ�/���3��͐��r��r��v��5����b��<N(Gt�v����ad����Mu���
F^�u��zXT	����L�L�`����3@ӌu��d��筴p4pы91,|L���G�׼�51�T��7���c��L��O�C���:�2�����=�g�9kL��j=�����B�Y�t:F���*������}�r�4���\��J}�/_5��ܝwG2�`�|2��E-�J�cq.Zd��?Eװ�w����_� ���v���8����͉��������HGJ��-S�
8ި56�L�6�դ��[*�k�t]V����P[�:cq��~
YX�N�^G�Vт�N�:G������h^��b^�8U7�����t1]��`V7^����zş�@	ʊ/��O&�ܬE�˱a����Ԟ�Kᴉc��cHt���{_���q~B��~I�i�AQ�/Gղ��Rt�(�A���X�Ns9Q��B�X��A�!�x��`)���PSfͲ��&�6��@W
�����Oe8RVPI�tN�,�JH�L�'D��u�2!�jQN�-�dI@AE���C�a��Ȫ&-�5���!�����h,d.Kb䋙r����t�L���<ǔT?,��硖V��?}��?��?����Fo�y��=@���+;���֤�ŕr?C.��*'*���"��*R+����l�k3#Ǝ7�.s]S�DC',�E��DȊ��pt6D��L̓�_7��*�ԓ�0l��H�����A�\�dST�
U6��6���P��-N��Q�eI���Y+֞=T�XYZ���}V�Tk�8!���=c��aq>�˥�>�A
�:AC�}����z-V��O?�����񵯾�o��o���X���z�ޯc�����n#jla�JAD�k�E���
�56�,H�$�Y(e̱x�|/�{��br-�����ɢ�4�r��s�!��D�8���^Q+dSB���'�Ttb���>��� ��\�j���K����SSA^K�˾N�)�B!�,Z}a���~���!Z��^GN\c�����3�0X��~5�,��ަI�z��ͽ���cx�)����������S9_�I���uL�U\{�W�����*�cJ�LG�]�seФ��V��F���s�S2�l�N��i�=��<��;�ق2��N?,4x�(���!�?�J3��1^co@M�D>#]h���t��d��d�PC����ȓV��g��i�S�ĬCJ>�-q*c���
ܺĺ�DйS��`\�9r��"����L�
m�h��}�jRJ�:#��	2l���J#0f�.-w�Ӣ�hjl���v��_�{��b��l���ʵ;�V��	P�p��B|�W����7�N����i�\?��-�++N�����1)��~
��{-�{��g�z�_D'e��)�@
N�ؔO��wu�ux�����8δ�N�+g3L9�B	��4�W�g!�(t�	�������O����Ro��9����Yc�LZL���7�r� #�PdPGH�XSw�E��$���wHY�Yo=3KsU�3�3� \��D�Z�G?�)>����O�W���Q��w���[71'��5Z��t��g�I��?��2�'����j+'�t���
�İ��5�,
�>��� eT*�:UIs}6���5n)�<~/������Ǥ�r���Y�AZij2
0���8d�X%e5�4vsy�_��D2�-9��r�x��n*�
��k��Ў���k�}��T�:I���\�|N�8��ipF��o�ue����ѿ�c<�L#6��<J�+���W����|	E�~����s7u��V�F3 �~�8�K����dN�Vߚ��5��v���և=	��3�l%%�?�V!����Wc=Ԏg��d}���:%�a�^��\�a��hl"KS&��G�RR�y�Ef3:�3��$��p�����u��E�c����j�0-�ު 
"=q�a_�GhW�(/h �7��f�SpKzY�ږ�Üƅܔy�Ph�ȗ��T	�'��|�*m��	z�gNtl��I���"�Z�����)t����3H��@k�B��(�q���FQ:�֢��mS2���HH2m�E(7R�is���M����5��3�hw�GO����KkAg�b�,��v[�nA~��eu��r��p��i����b�(�E�E�׃�S@;���.zgg_�	&�O���
��,�����{����:<�:1��0��x5��F[�8CT]#���uh9g3��i.@�>۸4(a5�9J�����*S���(Ɣ�ASWC!u?n�c�����1����ra���E�3��t�?�?'��#�W��F9K+��_c�wŊ�\Jі�m2���鯢%�����[\m�]�a���7n�/!.]1��r�'5�T����;,,מ58���ZC&���蓻���?¼{&����������w�{���/��7a�FX�CP�΃U�w*�dPn���\�ؠ2@>!�#}�}�F�kaF&�KZ����@��5g8j lr Z׮�C1�5�,����45< X+����Y�r��!"01��Q�x
�c H�P�#�Ş�l�K (�Z�Z��n'���b�n�o�.�n�k(ܙ׀�� F��!�48��{��@(kY �qG�'���8z����o"�s�y��O>��<���^��_�K�Zob�����[*�\��pd����۲�o�B�Z��ӎ��%jy�eQ(>�B_��д�?�5*��^����*L�L���`�"�4�k6},|H���dL��
~_�߬U$�+�9�:sN����7ev.z]b$/���B��$�V��'j�Zz�v�[�4YZ�A��ͦ��v1md�V�טL'N�?8�h4B��	�����?����6�	JY��o��uк�&��n"'5��`{{�4 ����x�	��:-��Y�ך-�#����O��&ЁS0�m�^�I��4�Z��I�Z��<�xO�9J���;��r�6�&�Δl��$d!��
,��8�b<�-iR`BM_�����06H�0�W(�Yc�H�qz�?��̥���WN��(�<�)
�9qoP��T�����?����i
��U�u9�8!0�N�����̃��9�N��H��L��?�=����õk71P�Bڳ/�����_�6�a���o���*gԅ�o�zpm���+F}�y>qJV�a�o�8R!����@�<�)���9�&o�O��ޅ��Ǩ$��l#�(�XY#H�7�djU�wʿu��:��^^�p�(+־N��
Pt���*6����{KdF^77g6z<;C��dU�I��X�4��X����9�ﰽXzd�kl�iZ�K��:��J��"ώ�����{ߡ�6�y��>���ڸ��;�:-�&#Tj	u�-�Y�
��Bk��g��]`%��1�:p`��b�����Jhe͠�F��l�b-�Z�R�bk��g�O�ʔ�ǜ��d�,��`�t��0҂S�F�5��3}|q�� �M��+s6���,҅�>�<6��a���dپ6� ��9�0�ձvv��Cm���b�{AЊ�L�m�43�Vצ�/�7�I�^�v_���}1x������?��B�ԯ����W�h��\l��!�BLs�Op�K�r�����.^Pf���aM��q.�SPZOkM��Zܦ���u���^w>�b���Ѣ�ش�L�
�Z�!�e�P�3�)X��9Q�1N�q��	.h�lLL2���%�M���Bn�����[�Ӊ
�����ڔ7��Mƚ��}&�>��!v	�vb���O��f� ��*�����ˉF䉮�1�q�@�c��c#�"Z	�e��ʹ�|1�:j�gI'ERE����B6)z׮���0��/�4,0=G��o��ܨ�nSrXBiM��VD:�^ț�l4�hn�R��3ݔq�5>��ԡi��V�\�,p�D�6�K͒�-�j�]��dם݉}����^��42�!��'H�H�Zٻ򔼫UI��8�-����U.˲�^�w5+N�0I9t��������sν ��9��i ����s>�t2��ke,np�K�����Z��T�p�9u1�Ml<y��'OQ/5󉍹C[�ܓ���109���	�6M��I�/�t�s8��fFG!�����J� ��K����3��8���S?
�I��aM�{�X�?�!/s>j��w�!E����`]�־��HS섘�0�<?�u��K���@B�#��k7Q�}�:���4C�N���Ӝr����ݙ>K��N�ɉ����s��0�w�j���H�N�%�&�Ι*t��&��W���-�}�
P���;3�d�_ii��o���mSOJ6�N�#@�=|ܯ� �����f��(��	��.��鉤�4��7Z�x}�D�y:�*{�.Is������D,�<)Rx;�Sd=�P���R:��qA�p4�|A;� f��n-��9���H�tBS�==s'�:,t�۷~��v���)<��6�By&�}��T�S3@��a6tQ�,9�����V�>�5�7�`(B�����EE8{���.Fg�A�7_2_�٘l�;jsOMT�b񤠹|<3	���j1$�:F��2U0�$���Ĉ�Q
b	�X�3Cȝ�*��t&֤i�Ȧ�g8�~=�45�q��r�z�)�]R"�rQD#@�Oz#��H]cSoݏ�t}�˙�¸�ߦ��:�w�X�;`�h=��]%�0�i��
��Q�{��n����#�u�b�y�6�7�9�h�Q�X��c{�6��.��1���f���n�4�����P)0=6�ׯDQ8����P羣Sf<� ����OJ�x��j��J��?�������ω�hjF�q�~v;����	tz�Gz��C@�8J)���<�|~�\�Q�E�RHIM�@��$4�{�Z�YuN_I�f�)@6���T;>��k4b�����!�'�'�_���Ϣ��W��N�7�x���nPD_��]*:�8�6�m�K`�C�&�j�]��������Xb� ��*u��")��I̾�]��it<~�NL�DG��	B�����d�p�D`�k��;�7�7R�%���$B5�,���s�١��m��ꌓ0M;���'I��y�t�����D=.Ms��`͖�5������{��+��K��>�����u���̩�ݭ</��#a�o)�_�G5��ե���/�Zz?s�}�Us�=���9�(��:�.|��V���L�v��i9�`����ݸ��;w�k4�<͂�a��%��)�u$�)LOO Ds�Qw�JQ_�,i�xszf�r���㝩z2�����e�fZ�����Pu���S>>�@������Hm:��Y�tZ�a�v�?�}^N�x�fPN3����ӥ�),'�Gq��=aY;)=X@1gaS�1<?|�2�g�����ɚ��j�C�!��Vt&q�+H�]�Ϩv�tA��
cM*�:�2Y��M���O���.��f�0�g��K�Ȕ�j�0uj��9��4q:���|^��qb�d(|3m��{�����R��ԌHhc�Y�j�(�`�}b�ĆZ�ʄ&ʬM���5��c�CƊ����+u�}��4	�M�Y=?8�w� � k���-=�8)���Ԉ���ߥ+;�r�e������-?��";�#�|��$c�ݡIU@<�ig�ٖm����lƩ?���Zǋtf�Ԁ���#MPЏv�X.h�R���3sL��xL�B���d���m@$���	:�ʍꄶ� DE/N�"]D@DH�8�=����:�g9$ř]�v�n��N�-�n^d�z� R$�M&���:��A�S]�����9������k78�-F݁�.H��ȟO���U	ٚ���$ԶbҢ�Ԇ��!��b4����?g8|10�H2�9�^��:�h�m��H6�@<�P*�j�B��%����LT����ҝ9��J��-\�NC��N�&4NQd���?R�W�%���Ԑ��ZG;�z"-����1�pD����FR��������[���xi��� �dѡ/;��5��]HJ�\Kp9Bkpi�x����+�|u��� ��Z���0�!�1>חU�î7���)��߇��,/�V��b��Dsy��©o�Z∧��O����E��_jާ!�2m��q��B	"�����n���J�$��(�d��8�؀���h44!녦/�!�(i�|�'_̕���ĩ?�q½����
�H�8ib�ůk7TL�EY�	���E�3����-F]�\ϓ{�E��J���t�τ<'�|Rtꢥ6�}�d�srޓ�U�|v�ZUt���������ר<���O��v��(�h�~C�ނC03��P��!,�"(���Q3��Q�b|ƒ�������>gC��v�|�i`q@���B~>7��EQ{��#���@���v'y�lܢ�TD'yX4B]ڠ����S�c�� �E�g��OU�-��`sH�}�!�Jn��N�����X�\�λu|�CЗ�)��g9�3J������ŏ��ᰠ�����qi����xz�s�=�����a?� u�,�"x���70��X+�5��f2���h���$q���2UUW���*���PB$�@(q�Ű���nU�5�GZ�P�VM�H���hL� �ǔ�b#,���ǲ��`�z�zW�PG|�d�@��.�1ҋ�(�Ј�D��U��ջ-tږLJ�*Op��"7*���u.�L�h��H!t�УY��Y��C�&�Ui��z��_'Y�#�I�3�]�tu���`�)��P�y�w �HZ�S˴��7?�9��A$���Ձ��$�h�^{G�{;�����i�k��D6�;�(�3ހ�H�S�I˒X$*?�5�	���PR�W0N�v�,!/:��o�j[�CR�ȹ�b�R�G��t*OP�& tэƢ�gS#�FX��"(+;�qh�{���=�3Mm�Y���\̗j���9CK�j)�;{_�D�&^urR7�5o�'UO[}��XqXҗI7fATK/����y�{Q�����_a��}����9�&�ڃ���.\E$�E�i!�IJ$ �/����Ӹ��"e7�~�xϙ�xݕ����d>;�f#|�2�dH�RXG��RS���1<i5W��0%="%�XY&rB��I��.LǗ��� �B�v2|�Kv�.��B7�*e����aM.g>	��A%וR.:|7~��N 8Nz �d���W8�����n@���	��E��U���6����Mۖ:�h� 7��KO�б��H<�\��ƾ��wd���F�?_������E�"H��ܬ	CQq���Y���I�O�f6�:g]�I�sW{ޣ�E��Z�9���&����\ֱl��n��������\$0��26�<Ը������^�����P����&�d>�3���U�Z�n�V��zz�j�K�u�}'��(e�@K�у8�E�Fr��9�?�_C��ވ�@1O������j�
�`�Yh�OĤSgA�$Rk .06^r����8Z\w��������§jD؉��
�\���L	D?$ai��    IDAT��:*M�T�����;	t�8.+A�<��"V��u`58������&B�R3�J��"�.P|�b�/�]�X� e��VLG@/G��t]�׎FGs��%�}�E��8��or�A.�P0$.S�"b�#�͎��@ ���gX]�G�VB��u�Z2��Q-T$���yDs�@(�x_?�>?:^�nC�g����C��37�Pc�F�g%̀š�W��.��F��\r����K�,�^��pڨ�")n>�r�{j8�N�\���
�ۡnȔʥJ�#�N��9�k}��n���X(�ܥ;�{w`� ��]F��+�����`�Z �o��05�!+��s�{�D�zE|�GB"�8)����X�v�Q.��J��B��i3}�{E�jv�MjNd[Q[�T�?��ق(�^�%b��i�L���$j��O:���B#�����ݰ���*M�ω"�RlB:��*�nݦh�E�RO�z���G.AB�Q*1�� M�!�T�_B� ��zQMN&x8��>�ˈ���H/=w�˿�M�N^hB��ce"���$���N	`T$�E�&߇�`���Z�� K��qbZ�����_}���=���.�@�l?�?�C�00�:��I��h;�����,�$?H�Qմ���V]։�g�&�l�I���� 'h�g�S�mI��W&3D��)�y��x�6��qK�gH���//榥� 0�F;l	u��&�����3�$Ȗ�#�x7-AI�}��G ���Z,q%��p�����Х��Զ�5r'J���G���#.�^l�m���%���LPQX�73��D���|�:�����	��ß��?�1����O�9^}�'x����_��k�l���3�<4g��1=Hӭ��F&�X� 6w�qtR'f�6Ǆ.ݱIq��(�D����A���G8��Z��Ҩ
���S�ⲃZ��J�,���&����H $7�^޻,�	�6ESCgPV�"L ����>�tUeC`�BSb��*�Pf$!�o,	B)�du9����+tA��{ܙI��z�^f�j��@0�E)�+AM�Sz��FTx�愑~*qR�w�yc�g�oc}�!�|����P/�Kc�F(�11��6��z����$���^�Sי�	'	[�^��+���9���ґ�D�|��3��b�����`GP�w��ys�L��a�L��H�-�]�n
0��p�ۜ�,4�� �.� �8��� ��	:K)�c95c�F��%�P��!�d���Z!P�($N���֌^X'3�g���3B�H��t�i�shn
�j3��#���B�sCOdٷ��fB���]i���F�x� ����Qx�&0q�
b�<*̋�$1<��P'Q��3.�j�B��9��\R��W�^���A�f��t�=l��M�g���ie�H@���#��V���@�e�=��Tc�4sUM���#_ℐ�?���:k�o�R@T��K����c�y�#Q���L���՜����㞒��䪪	�Lr� ��;����Ȩ\J�P�e�0�J-k�C�t�e����蠚�%p���k�����iT`���T�^~�M�!��#�T��jNF"�P��mUE�»J�k����B�m&���(�.��e�*"�Ae��6!��iʳ�:��j�%�)�>s�LI�j�3�TsB�F��ޑ�n�\�ܛ:a�(�6�&��QT>�w!�\N ͠ �.��j����O����^��s�a���ܺVAt2\ݱ�{y�H0��׀1�o���S`�q�i ��!J�W�B�Yb�!hZx55/�_sDK���*�gYl*�碣.B�!�`E�@���P/@��|]7����+4
������\ܲY%�R�N����R�4t�A�)�jӉy8s:(�&�t�q���hZX|ЙN\>)F2�Ls���#0���8"�
�˄n`���
��Vq�c�ˑE;�8�hQOjt���)V��k�P��D��u��z�A�6S��֞���H|��Bnv.Z���)7���]+'�ն$��Q�c�ϬZZ���<d5���&�	G#"�}֦[.t�tq+�i֋��ب[�M��ch	�!t9���fQ��:dx6��r����Iy�c�6|��YY_�*H��T(�2�c���Ѽ��"�!E�Zk���Ud��|o}�$��0jGǘ���ކ�*%��/�Ar�2#gH���dH����P	�$a�,n�P���礁ȰT®�H�F��/$H�d���t-):Y0���^6�\�t��M��!/UN9����ёϋ�"���BXq�wn����5%f���sZJ�o��#n���p"�:	�V(��?aA��P!ঞ/:R��>��	��\Z��e3A�����@(�+�J����f0��[��xss_���c؇k@�
�ϖf���!:p�ɗHN"�@��0:�vh7�r��Qq.�g�TKhZUD�����`�dP
�(�f]����r�rq
ED�	���L���8h��k�&��"̰͖�J�	_ �H4�Y!͎C+�$]�T��;
����k��Z�"�ၾ4����A$*Y�UqxT��QA�/|&�YX.P�yqހŮ����|�����uy��;g��	���	;�CI�S����A~�\7�(?kO6�پ4��"���9w���n���_{	����g�{�B$3���g����#��!7aU����&ͤHՓ�w�҄�E*���IE���Z�T�>(�R���!Ѹ"�I�Bժ
���G�iUD��L���;D��C�l��!��#�h�f�э�AKs��zU���A�U+�V<@4�����''DD�x��bq}�Ff()�#��J��]'�_��㔉g�E�7
p̳�%�-�)�̚ջ_�heJD �l$ղ˽)Y3j���0��W)��Ь*�G$B�����3l=�_i��u�m,�c�e�K�܉��ȥ7Ȏ�I!?<�Xs�RQS\)͆h�8��	���w�����@6�N�y&ţa�kU9a�!uƙ02��r���	a�`��-��qڣ�h22��*Ʉs���3��7�uI_dCCF�:"v��7��T0)z�l~{��f1*͹4dFB2]�J�-��r2A��8�>��p5�*�!�����em��Q@2��ZX�blH�F�J�7"�Ҍ<1Q�� 
!	�z���׿�­��."�m¢�6������+H�P�ڈg��J��a�4����R��R����_u�m�xZ�8�~��m4���u%��w*�ЦE��@,���ޗ�x{��a��?N��tm����E'>H�vO�6rVI3H�j�H�n�y�lTCH�҈G"b@S.3:��MDH����5�����!��e�C����jFÿ��{��)�k���S�5��O)��=�u�X)P.g/��׺����D_*���|�чX��ڵ�4�j8�A�o�/��F��D~0�t2�p����7�AN�Y�Fh0�em�F;�����P�	B8�4����r�v����8�AJ]��fͦ.Yw@�� ��X� V�'�:=�	�4��<kDH]��5�%��|DN���c��c��\��2�v���_��p�0u�.}�ԧ����hf�2�,OkW�=^Xc�����C�v���tԋ�������v��I��,&���f��juFj���"V"E|8J���@m�%��Ȧ��NlNy&��DM�!S~-}�8�J���"bs2�(�v[�o���DH3�p����+2\������>4i��	���8�PwA��4�`#H��R�%v�u�r�\򗓞�~����L��=~V	u7��8��(��RdL��"&�	�zq�%H��K䤊��9�<}�v� ~�O�!��"��Rw�Cr��}#��3���6�B�$��gr���ʬ���U�i�l�@N�d:�1�3��4RX8)���`"Qtj$]����%�	�q.Au>u�{�YT��&:����'��K�M%����m�z�Π�ʔ.����%�"������Q���DP�M]�η�ޭ6V�N�~�� �����4Xy&2YU�Wѽ8D�A3*�e��q$�Q���0w�Kl���c�X��g�Erx��0��z>%NhP#�����hYu4I��y� ��"��_f�R�R]	4(��D#�K�ެ�O��ǃ���VK��X���!4JY&MUct:��͠����總ȹA�ef��`_I�Զ�=�}6�OE�Wy0Cq}�^�'��F�J���T�nŮ�����͠��FW&qJ��VZ�Y�� �����s��Hs���&%�(��8l����9<��);���_�ѫ����Qi��9��SW�L ��?F�v�N��l2���aF ϖ7P�5�JE	S��E�\F�X�׌!�f�D��P{W�1ח�����
n޼#�&�T'�
�R���f��������j~q'e3�.��eP�hT����������[/�Z<@,f��)\8;��<�<U[��[,{����s+8*��f�$Po٨�a��0nri��d�5��S�9��<�h+Z���Շ�Mɷi�߾!��͢� 3���P�Z�O�c���<�������l.�tj��WNO`n��X�\�\v��F��t�9�$///c�@h�SS2]���`&׏H�O�+�i�
�hԊhw�ro��ʕ�{����}Dc	A�%6'�����hW��=;�K��a{���K�EQ.�0H#��.~E�,`QG��o��3Sø8;��� 1�<�l L+��G�5<^X�I��f��%)8���S ��� %umG_^j,�$��G�rN˨Y�y)�~�t6IH����&� ͠�3jB'%q��v��D�H�R�}xv�6݁�����*J����h�A0�E�bc<�:����,�}}��5�z5�SF۪�Ε9h,�kժг)Հ����Ĥ����V�T�a,B�TB4A&�F�(����Y���(j$��9qV���z������)��G��ad2qBKZ��?���G�v�t��C��Eg5l��pt|��RY���C8�Gx60b��S����[u����Q�E��u�4��DF]���s�_�A�3�Uk%�筒��4IFè��W�c�kh '{=t�ax2����T�(,ۋx:��P0,=K��F�`J������.R�"�H��w�D����i�񠳫���m_"���ਘ�P�7���A�Q��4[�x�FFdb|\��X�K��I0�cGY���罣QTj�e��-���^`d�&sa�y�x�F�����%��=��"��Pw����'ެ���c�ˆQM~�Hy�/&KJ�t�N�����*�aH]���2��pb0�Ba���ꗘ�y�JI��4B�D,:0�鋯����D�ןC*@8��2C L�.��� �Kv6�P=�E��ʂ7W5�T:���tjM�*���9�Pޡ��p߉!k@��8�}�g��Ԩ:��s���@��FbX�z����y$(ó�4QƊ0S�5����V�*.Z'���k?�K�A�Z��O� ���G\s����E�=d�a2�Jp�%'��لq6���?�-���'�����	R��6�
VP-�Z3���0Y(e�R�#�}l@�窙rܚD��,.�.���9.h��`C�#��x� ��`�*$q��̴wc�e�:�t��|��tQk�L�ްв�M���In�N�A�fx���+����j���D��&͑^�ڨ:K�@�ǿ&�;4ZË�0��DD�AN�ăX."lڝ���Qq(Fn�~�@qm[O�bs�1Z�]�UIn;���l���,�A��4�#�0B1q���k@ےw��#!Վ���.i~��U�ӥ��\HY�3 �ϊ�.	?�UPrY��^���'����g�Ti �e�S�iƔ��|
��o�k
���tGAM�-��!�QR
]�Z�J�P����:�ѿ�9��s���)�r����~�<PT;(cz�,/��>"I�ɟ�JP����(_�,T�\o���M��1�M�t��[��5�����.�t���">p�������f�	zą�k����#��'�^�$W?6�iq2A[�����<iza[5y'�8�o$�����aɞz}�y��K.�2��l��~	H����SR��4\5��AI�R�\��CD>d�q��E�NF�y����s�b��Jť!�)���-����ԐWm�t�&��|U�4
E�[��	��3Gp�}G$߭�2C�Ò���!�x�o��ˤ$��M���/�+l����V�HtC�P��������G$�p�\>��p�\>�SS~ll���_%����m����;9n�����{����i4��� ��p�}��es�r��t��ln�I�B:�B~��J��J���^�z�x �������-t��L(S�KC`��|�dm�o�g����q�\�RO�cwgClq��K��E��R��[��9�����Q�5�HH�W��k�Lp�[�d��!���Kq?�x2���mDܦ��r����}�(L:#=�A�Q���]�=���<v��8��g����OPڭ"9y���b>K��L1l���\�}�2������o��?"��՗_����$���b��c{�پ)u�5Y�᱉x+{%O�ʕi�x������%�rY��ci��B�V�����P�����[�7Pmz�ńzhj�|)6����G}�6Q*���� ~燗0�ai����c{�@�����ΜB~؏�����+�0Y���Kl��	�;NiVί�̦[�cd"��r�^W� ��4=>�gk28=J�Y�e�̆�C��f��N듑6�b�֗��V`���V��F�b��h��OO��̫dGHf�L'�zaP���(&�pR����G����䄼�lNN��{ πك�h�ղ����W��SSӘ�����6�7��$�TL��c���U��rbrgf����*��KhuI�j`���4R�LC�-8Y��U��ed�̩)����M���0W�tB�zO�`c��j�T��*�2q"���zM���nԩR��-�z>�!T�<��x'E2ݡ�^�.IM�eF�H$�k?B��u"!6�1Ԏp���xv�s��������Iab�*2����qm����q��&F��5M<z����u̜����q�'(��Y�����3<�G#�f��q��á0�F��R��Yǳ%v4��!�b�;�
�lBA��H$<��iaayGŚ�|t�f�'� 'G��!O6�v���0�6�\<���L��;{��=c���~��1q�^_;���.J�3��?��C�^��%
��+NKEC,&�!u�����s3��jR3Dm���p�M2#�����6+�"]'���K�ˢ�w���s<��K��e�¨3��d3�4� <A6�Y�R�6|F�f]�I���ԳҰ�I����*3f��������xf�302��CJ��c��s�Ds�m`c�8i�NƠ��|N�Os$iRO���ă�瓗�Ϡ�Ғ��M=��8cF�Q��*��T:(���v�#yu5��ǣ���o咪�L��
j�#�,K���K:n�B�V����G�G�6��� _1�Y��Z�����{e2��vӦ�[ݞ�D4��O�hH��	�!E��N�jS�`������/�G���n4���|D�x��#���O�.�N��TG�ǃ��{�
^���5oڕi>�0l�ȟ�k���}��F)��p|RG�LѯO\RI�cΡ-��̬Q�H��:	�Eǥȁ�܍%���B�Uۤm+����n��א�'6�j�*��6*"�iz0Fv��Nխ�<]���c�
;�u����ַ!��q�\�7= #�Cn��f@�=R!�3Wt��2���rh�*��J�ea-_ZQ��N���/7��D�upR��"K�ɣ��D�F#V�` �L�F'��)V--�t�ꚰ(�Y���h�ތS�6�9MMa|,�X���=�j-llV��z,!'��J�O-4����I��6p.z��]����^�s��p��:<X��N�H�2�eo鈈�k��M��V�QS���aL�$Q>*���3,�    IDAT���_�]\���A�Q�~�F�"=z���x�)pM4u�a�ɼ;Q���
�w�sj}���&a��B#a~VǪ!O�a��Z��щq��rx���B��L�Ol�Kt���I�z���(��p\V*r�C (@׿f���(��E��es�v9��ZfO�Oqf�S�#H%H����A�
����ۋ��)�Pe�I�MDc1�0��5�p���;�U��jB���םfP�[�ۄ�II�k#T'�����~UJ.pG�_��@m�`N&�O�cc���#���Q��@�nq�$l_�ɋH��"6�g�����
F�(X\X���g8w�^~y�r��!�͎�不��/��P�Y��T��:�lV�b�-fH2��������>����u�?w��q�8��@�4P8d��G0��־�<\ǳ�#�ڴ����gMm�Ќ p�5�=�u�����E̞N`k��k_^���3��˃�3g������t+�6>��v��I�ж9��}�j���`�'�{�	�i����K`C�3�s�_�9|1��'�K����vڈ�B8}j�Z	O�����S�v������L��K�q����� 3v	��H����GWG�իgqf6�������9��λ87;���#q����!>��+C�D������2I:����Q����E l`k���?���m\�t��6�T���zh2SVc�H���;[XX;F����H�H�s��h���#`x�@Va��o�s�<�_��{ϰ��%.�d6��U��I|�W�a��-���
����zc��t�y2�d������
-5+��:KP�t���9�X�6�tJe��B�.|z<K�u�lIG��T2S<�E|h�-+)�b��� ��k���%�K��n�k�10�B�QB��]��?��ӯ �C0�C"AЮ"f6q��8���!3���|s��G�Λg�ˆqR��<z�[[[b�D�2�lR&���q��ߟ�`�B�<���.Z����Q��d��D֑��� ���x8����]X�C<��P�I	�ǜ�h��ݭ�^;A<����^�2�F�X^��o��fR)LONbp8+fDKk�X^�F�K����Ή���� ҽZ�C]c�|(9�4T�	D(�Bk�^dA��`������|8݋�$�;�#J��(��${Zq&�D�p�;_}���?A�xCs��@��&g^E�Z��h:���<�B�.^�|��k˛�4�T6��~�*lo��.#�׏�t;X�_�Yt�/�s��Ȥ�����j�c-}&J`ccO��Τq��8��1(���P�Tʇ�Cϖ��}PDSlX�06�2u�eEBU�C`��d���`�ό�V)b}y�Kk(�G0<0&�SS2�\�:���h����`u��:<C��f]�8]
�)�5�c����r�,�Jq~W���b*Q0N��e=E����?}�JÏ���G�� �|�H3X���{��L_~=1t2�̇൫��$�a���xBX[YG�^����`^�ի��P�	&	�@�1m�Ȓ"�9�#ߟ�s�\B�X�A�V��j��[�UR�L��v�a5)�`mjJdF�-b'g�QOl�YsqC�-i�^�E���`!2*B�k�TY��n�Mk��D"PZ�
���p5�*��|Rg2(Qb� EP�]�*TW~)}^�!(P�z².�����6�7n 賑O��y,��/�F/�B ��	#�؞���*!�%c�KҴ�g=b��;@8���n�+��!�ì�NVC8�A:����	
%f�eĹTÐY(}�ժ��/�|�GG8<.#MK�JM�؄8M�89dN0�`�����10;���iL�&1��f��$�����,,obk��� Z]6����|6򉉐S8�:�^���A頚����$=�4DM(d|�V:g�hJ�[�����%��p������&Հ�|Z�U����bg��(5`X�0�,<�/��/���o�`3��"?>..�Ԩ�85ه`8���g��;D>�E_���r����mT[�I�{y�wZh5Jj!o�d��x����h�:��P\��v�^=˒)�ŋ��p��:�N���LeU���"�u��Z��U��j��H��}�rv�H@�h�,|�
��<X���6M��l����3֠CG9����
�� .�J3v�6��̂Gh\�t��g��'ټ�4She��u*}I��j��p��ΥQ>�ǃkb��gh/|��y$��z鱋2�$���i�,D���B*���6�WW$�a��(FF�h����<���6<�Si�b4���2L��ig/]��s�}Q
=i'��E�����z���ĩ3Y<~v���2��m�0�N��[�U�:�v�!��%�gZ�����?���5�}(Xx����x~L��Ʃ3���Q,.m���%JM�I4�'<�'Q�Hba���RY��r *��C��		��*x�Kt	i�nv��KҼD�v�@X	���E��H(����Z5������=jG8^�G�`K(��`]3���9ćg�B6���ȧB��x�b�|���� O�_��&������s���pzv��\ó�2<f �1\�<#� �TG�a�+Eќad����� ��X�DD&�tӣu=��IQ踑d��&Kmt�A��M9D���T�	�U�tj�zao�>��q�����ƕ+�1=9-�ȝ�}�{�P��?�����$����[��`{���Q�y'WWJЧ��_�%R�Y�-,��xH��63���E��͡ڰ�s���s ���:�h|�i#����3�Zu<��5�6���.*��<=����.ocw�*����ً�H ����~|��s��K���������1�ٟ���(����+�/��ϑ�O����_�R�j����@��:�� �U�1Chw}88:A�VA2C$�(!�QG@d&�_m#�r=���C� J�&=mq�$ ֥W\��^����N��k3x��~ܾ�?��_a ;����=��a��6�.�c~�!��8����Jae��_~�D �P���QXh���w��:�zU'�!��� :��4�]K�W��	�1�D#g�jQW�мx
ޥn����n[v�V]'��R�0��ޖf������&���2:�=@�H#2x�3/#40�P&�X"����T�����
��2�a��2��~���ȥ��q�6�K5�;	����'���kHƓ�����tA���j55�`����=|�����M\z�*�&��� l�1����yp��>�6�h�4���)�%�y[ܓ�6f�6���&�曓�4mܿ=���i�8�a�o:����^��LH>�����dJp#�\���.ռ���q��=�����A�_B�s�G�q2�]8U�y-n�P�E?/@���l�Ծ�S�0�i4K���S<��Z�@��y����0y��g��H*���$��&F��%�(bo{�j��^�+o����
~��o15}?��+�ܰp��]�������:�h�e:�	�M&�d�L�X�Iݙ�Ea�"HMe��ZK2�mO��U�K��
|K}��O���� ���U�\ө�\�8(&o������*2�Fe������$Ξ?-�GOV��_D�6�3�0��%#J\K�o�q�Ɇ�˴I�����h���Fr�Ӵh#:�%�'� �J��ur�$��B~?��P98§| ��V�����.z��`��[�FShy=��bt���c���;3��$��;�
�428�ɉ���X��<��޾0I�O&��Cr�t:�� ?�F"f�\n`um;;{���d�H�C05�tj�fcHe"8<,����ށgZX]�m�h�Ȧ���=ЉP��8uj �l�r�'�h�4�J$��%�N]X�`k��R�*�������̕ڹN�:q�ut�u]+�+�_G @�?W;��@�VR^�i%{$~F���u�O��uc���=����G �XQ�D���\և�N#����lon#�J���3B=<*biy�y�x|�R׀ݮ#�Z=��p�^�����?YC�}b��C۪�G�"Q�v�ヸpa
���ϯ�P!͎�����m�j�i�A�i�vao��>ҙ8^�z��F`t:�^"��C.? "ߕ�Cܼ5��*R0�q�S{e
|��l�v�=g��i��#�Bk�$!E�P�
'Ӆe5�XtE�"_�	����HD��8��M�"3��it�8����S��=Fugh�	��c��$a�q�������e3H�3hՎџ��f0:ڇ�b	|��:~���artX��ƭ�K��dI�O.�l"�ɡ"A̓�w��qjf�t�o���U��yJcz��X~��.�`b��"� ����g88��O�!
/��)��LE�î�x����f��;ѵژ���g�X]YA,����8N��crf]�ۯn���5�#�0<Y9�)�������J�<�r�Et�n02%r��D:����=��ԣ{+]˜�RE�8gç��P
�4Q�&�ϋ6����v��&��Q3���{ױ1w��eѫȒ	���x	��M�ol\�ޜ���� Ю�ڵ;��;��׮��Kh�
z�hԼ��(T�(Y@0�Ջ�0��i[��_�N/F�2(ּ�~k���%��+W03�B�g ��eI�;���	`q�����::=���z<�ð�,<�֫e$⌚8A����\��;oa$���۫���i`Z]�z�T�^:�w޹"��ϗ�����T�� ,�jج�]���@0d�Z-	=���msz�=I�!��A���.���d�� �V��T�q�eG�"�l6�����՚_�������|���Q�^������p���ҡL�i��P����Ͼ���YD�)�!b��۟�-4п�����+/����XY8�?��X����?������,n�ļ�U-��I�z�f�.�^1	!�K �6b�8U<A����g[L�fP��M�'y�H��L�e2H�rC���X��5�H}�][��� �~�"�?����ς�Ξ����}#CԜ8*����>�����f���s�o���[X]?����ڞ���Z��*�%#H�pw��k����"�$HD��!
�~��e0�#�n1#�g'��9���1 �Z� ��Q�B���:�A�����l-�Ga�)N����P��mOV��]Df�2R#30��A4d`z4��5��g����|��ﾃ���"V�����]���8}�����	�ɀ�*�-���5��n�c2ǐ&R	$2}2maQˆ�*�� б�ɗ��I��xf��j� l_X&�4� C��,��h�n�k�UW�O���?~+����
G'����L�I�!��������s��{�bt8�������:�� :�6�,�H#��Z֑�Ό��`k{;{88*�C�?�fÀ?�Ӷ��R��w����Gv"%N�D
&q2U��W�6D�LWO��k��N�П�c����q��>��#��B�?-����*l#�`�)�_~��a ���&௢?�ş�W/���g���uuN͜���&66��ů?�a�����?B6��W_��I��l>�<��c(O�h����T( ���^Рc�7�J�X�Q4��z���E'�L�D�l���`�6b �Ed2@��bx{���`x(��5-S�o����sO0��ų����SƳ����9uv.�C�c����a0:�c*E��	�C`�^)"ߗ����"�4��d�qH�K��$z�ͦFD�9F�����$��%�.��l8�%#C>�HFR�g�<)�ޗ������n4�"lZ���0�Ø8���Цv����4f3Y���������������}�)\�~w����/���^��z7�~(t�A'?6%r�TXj���_G�E�$�8<>�������rH��N�k�FI@8�E0��.IP�Q
d҃�L�ji����<��|7n����F�0{f�TN����M,-,�g�q��iL���Q��~,Q�?��f�S]�F�t<���M�ş��#�ؐ�*Ȧ�ψ��0���C�������k\����]_���F� ��4>0��a������'h���#�,=r̉|�hm��c���n����!���U����	�w�0uj��yT+4�ed3#��z��2���Ĝ����h��N���Y�����O0��f33���Qw�����3��`�]���>V�vд�%��cChj~!�c��!�9�hT�Dk}������N������=��D�a���2eju��>���zdq�QX�,f/3��5�!^\���z�=)���~.N�H��<qh�)2��J$}��6
3�S�fd�3������\�D�[�1����n��5C2��H���M�&^{uJ&V����|��_}��#��^��,-�⫯�Y�JȈvr(�t�'#�B��H$�s��/�u{��.�dafb�� "&��T��!���q4{n?<ƍۋh���yB�ET �U2������x:�H'����E\�0���Cܿ����Ң���Ĥ�F��>l��W�F��G$1,�)�Q�Qk�,#4H��;�/m�,�	C�9`R�}�4�$���B��U�]j�"�H�ODl:J��w�PR	<=i�V��r��G�m/�n���+>o�^;����Gx�4}9����U�|�����7��`nk�������j�"�ݽ��gg����Ƴ�m���᭗/c|(.�gDg�9�!�xpT��p~K���\�4�\��0�ۋ���8,F>�{!|��
�w�0|I����S�.�H#:B]g�d���Q��� �W���G�J|B*�A��"�-���e|��Y��|�˛��!j<�S]c8�
6�b� ���5Bil����l11��H{��������G+��� '�N>I�=�k���L6�C��CE�j\ZU�R�(J{[X�s��o���Sֹr ���yd�/!�E$�'(���/��*�0�V��a����Oބ���g��g�Ϧ������G����<JMҩ>\���Ԙ_h�L�A/�08����^Ý{|�&Ο��h?+�zVS��F�v�d��j��.�ֶaІ��E�T�x�*�=y�	�Q>YF6��w^�������S|��O��8s�,�}y�TkX�Z���fg���o"���Ƶx��#��E����&匦OY���`.hK ���x�O$�פv9���U���]���y�J@8h�/�]��R����L��D��f���� :�6��ag��K3��ѡi�p
ѩ��=�2�gN$ѭ� ����w�N��7��888��~�c���)��g_c{}W�/^��������V�ZM�dW����arjT�*�fS'q\(���Xm6�9���.����HvۃN��PЏR����bk��x�m�X��& MW���&���-�ru?��(�][�g�]G>�?��{8>l��O>�w�
��o��Q��W^{�{�����/��?2�I������l\�Ed�&��O����cmy{'�:��dyPk��� h���t�� �D?#|��
���f�Q#�Жg�bԵo7�9��H� <ha��}iW���.F�==�'�ֱ�]Dr�C�ʍ!?8� f"x���������{�����}������C�-�❷���WfPo����qP%%�Ś�D���Pgg���P,�pTn�naa}G%*	ɾɥ036,4y���`
��f��nbe�ڹ,zvH�	MF�ѧ�[2���X\����*�x}_|�_]���/]��������/�R���=�����q\(��˗�?:���'�~�1��,lL֞hNL�D;O�qnz?��$<-�rk[�X>(ci�^o�0�A�.%�͐65'����2Ab&��@p�hz$|�w�I��H8*.��t�T��~��9�����	��.��CNu���1��$e	�Sx�d��|	�����������>^ye���M|��L�;�����|v���U*��J0Hd�<'���n	�N@kgw_�J�TL��y�q"S��e:G`�4cL�j����|A:f��Q��    IDAT�O�6/�^��x��.^��ٳM��Ï096�7^�"�5M��s����z=/�^<��g���^�ùE��ސ8���;���U�Y�����[�XG�����x1;� �� �E��/�v������>�k!��=�Lt�m���s�m���f�ϢuT��/�����y��D������؅7��:���G(�`>�������su�b7o\C*���o\B��ŵ�7�ze_����ɮL`ɒ��{�ND裉fF�T���ޱ���#��đ�%�{��F�g�6Q(���{� ��z���}����Kg8:5�]4*똝���)��ϯc�o�qQ�f6��ͤ���P<�����|\}����o�|��J]�����U Y�d�x:"����O�dڵw\B�Օے]�{�W!��d��yK����]pL�ڄ�$��yn�(+`ʺ8��bl`��*>�ůp���A��-N�����I�0>{	�H=�#C�g#B��wf���p��5l��#���w�D*�'�\���*~�w���H�~����}��@�����%��
˂ }0J���
R��e��E��f�6	�u��b�0?�IT��l���&,ʩ�@�QA� ��2fgFp�t뛇����D_&�H�f^��mu091���A��?x��r��lL��~��� '�sI�4�!M�/ԍ�coFi��p�!����|mЭ[#��>�d��Π��2�_�T��F�QjG���lׅ2@"�F�����L�W��絭���c��h��3� D��DQ��>�\���\.��\>u��>G[[�b @䜁F����[ўs���T,݀D�
���9�x�����Vf��x��ZN����qW�<��g��[���/�(%�l�����Gv��[�D��d�2�˕5�K���Cp|d���6\ZdW�'[�]Iջ���G��$r��?u��r�T-c7�����O0�����e._�Its�����?��F�D*KGw;�3<�˽�ܽ�@��fqkV�l�)���-�tF����"��t����=W�>0�������d��c��!2�P]�4Q-�	��p�m�&xyK���F���%��_���)��j�,�&��j�C��i��n;g��>8FO����_��۴�6���������~���+>~�O>?�חf���%~ɫՠ=,�������b�mR\lu�)�Gή ��J>�����g�J�4*5m�dŋ��Tq�̉�ͥ�d<��xm?��s�J1����g��۷����+�B�<�G�g�\�Ź���d)q��n����çk\�������)���I��[�3��m&�^�l��(ӎ:|�,K��C�B[�܁b��\��O�"Ͽ�{�aP�A�숿^r�a�ZK����k�L߿��ӛ��f$S�nؼ��v�2��a�~=\�P�3����{\��n�?��s����U���'��[�_����j��_��N���r]JY�#*$tP�.K�%c`�P���X=zi̤"�ʲ`(P��S�X��͒�Ws��*y�ι�����*M�Z2e`���lo����ݜ{g����˟�V�|��I:�:���/[X�D�|�K���߳��~~���?���E�"Wq��=s�S��!�a'�[�D�I2FQ7�V�(Pu����i�CQ���jo^�$!��I��Y6�2�!L;6-��X�UQ�����R1���$�/�Pޚ'>��JR`U�����	�M؋�y�Ϗ���Z�3���s�/��%�ho'�U�O�3C�C�n����/r��$fO�ne�v��NM0����<W�g$?���3��x���v��r��n��d4���vn�̄]�G�\�����&���\(Xaq�s�e������b���{�	59���ϳ�e�������~���_�]o��.CC\�t��h\sʿ��c�|��~ ���Z@��}I��F�&��O?<@��I:Y&�3؊�Y�1���4�LV:����r�Z���,a,؝v�Ŕ�)l2V�r�^ZY����r�R�b���M����t�-� ��]�팍��jz����}��� �5L��U�#��9qp��{;��J��KY���3}��12;�n��rz�+�Q����S[Q�k�i��q
�1O��$W5������i��}���?*xO�V6q
¾��D���͖]�������1�D+�
�^�_�53�X���ק�9���?|�������ڕ�\����Q������)����$�iZ�|��Q*E.�!��auIlC./9U^�(�K��o�ݣ}�kV� �K�3^.F����\�P��(	��n��p��R2@r�ЁP[�=R7�N�EU~è+�B����!϶Z���f�B�=���Yy~�Z.*/�b���l��T������v�� ސ�j%��]�����c�ţ'Ԋث�ȿ�%��ç�R���5^��W�؎ݭAF������D���Ո�*<�T6�vB�n޵���^���q.��B���J���k�I�e����2D����4�-Zr/�s����c��#����e6768���^��bqi�޾nF��x��)�s˸<>>��	�(\��XFȔU�3�R]�qX�8�o&쓳?��f��h�X:�p/����u=�]��R]�*��zYƙm8�F,��:��l� �}���)勄=���)G3<�vUm���4fb��n�K���]Gi%o�a��ik	㰔�Nԅk.���aǮ
�����쥩��t���gs,�m��G��oim
�N�M ,&
�,OH�͒�_\� �fϞ��F��4�$�[Y	�	�03ae%������j��(j�J�Mɻ��X�p��0~����o������;�Ó�����>_�s�Oc�8���K�d�P	���tؕA@ R�9p[��Z�sp�(#=��I��J�Y��،e��!�`2�<W��*��/}��,��Q�1��u�c}i����>�ᦧ��|4��o���UW��H#�{[�;��4R�:h�l�!��TI���]�]n]������8��D���o�%���G������i�#}�L�&�P5���w�R�3Ri�'^o�j٦n��QЎWY��KԷD&�2H��Z���)ճ�JOu��]�%��D��V�{�J~����M���ACP��W"LO͑�dصs�Ξ6��#,�Fɖ�T�N�Pһ��H���oT���d���d�� bX^�Yf�Z���"6�#�x���6�+ݵ*��o�wM��Z�V��?�
Q�N��ό�b`��w2Z43�tJ^0�[�N7���ep��7_����gt�u����1�⋯��ū�u�g���S�,l��H�Z��f'��y͸H��jr����*�(��핢VXe��)aKa5� [��VW3e����CY|�ol:DiNSR`%����&cC-|��^����"[ڷ��#=�}nf��<y�����!?}tV���}����,FՁ��b�k����"O�Z���%�K�J&���j�bp)�߯�ΤV������7�j��	��R�f:|Cn�/X�j�}?bk�BK[�Zqb��6�e�o`��1�0(o�������8�p��bu�t����_�s��5�L��?�������_�2}��IN�s�o��r��+K��	0�]�g>��աvy�b�����ꓶ����qZ��;#���Ɖ4i9��6�*5�tJ��"�M����wI�]�tz��V/��|?��<��/_)B�С��6�MnS+H�o3�\�q���o��܁0��=����&�f+����Jn���"s1�@g+�F[I$S,,��O�3�j�5�=u��x�MV�JP���rd�h�7��,���dA�[���d�$�*��4m-�>/��%^ݽ��T�&���Om�ݻi=���ׯH�C��8r Ƚw���Wtw����qy���m^L�����_~�g�9��|_���b�J&��Z���M/W��e�5���d���ŠgR��1:خ�iBx��if�Y^KP�̧�EZ�.'	�W�D&��26�d��|��[�5����ܹ��ϝ��<�7���2��F��dni����R?3���g��4��ۼZޢ�l$[�.;Q��Q�n)Ე�=����!
Y��Ģ�O��lwk �"�5��ེh��n��ȖS�B�M�e��B+X$ �j�W���u;�ue��e��V^�Mt���sʱU��U�v���-C�|!�����R��O�ȡNEu��5�<zō�f��],���jaE��;�uS���]�>�������z��e����'��g� �����Y���{b���������Q̌���?����rc�G��9ØŒ[������LU���\�ΐ�_�b��x�o������/�v׵�,W/_��ǿ�%��o/�$�1X^Y���r�x?_���� HB�Yђ�Q�N��4xͼs|�j�2n���M<���å�ڕ'�&�3���Wޢ�HF]���p�����!�rm�"�R���}ugX횙�a�����/�,���$�'t��2:8̫�%�7Ӵ��߶��;HKWn��|:Bk���F���YZ)�xr�;w028Į�!��7���ԟ���]����p1��9W.}O&U�����O?gt���W^���#Ξ<©���?�Q��r.��),N?����;4�w�y�b�[�$�R'�]�>���b���ӏ�������;DbIv����]��G��_�����;ɋy���K�<�Ξ>Io���.>aj)��۬9͢dW�f�v(�Ҍ�����^jY^հ���f6J|��M
���L>�9��+���"�=�ou��Q�E]�n�"ʂԬ���L����ب���G<�u���{T��n���B���$�Z����]��u�j
�kP2�8�=�n><��O�|V�p^N�r��C�>ʁ�<{������8)d�`�`�D�D"J�b���c�;il������ĢIN�9Jg{�����霔*�����%�<�Z�<������2*Ö�T˅�L)e����G:XY�r��5].��Y,/^df~�#ǎr��.<�bjz�h,�{�cx4̭;kL�oa�{)���\Ȉ�$�@k%���V��P�D�%V�S�lF�)�B�Љ�+�O%�J�E,�Z',à]3��V��r�M���i�P��������s<�z��7���5����� �@ݻ���?FVD^��a��R��6c�tu6��szf���%��u����>)��g5�'5[ပ_|�������#��U��}��0>1����>���Miʢ:ݾy���u��%m|� c�],,y69��P��,�jY8��f'�l��`�s�����EJ%3��������"7o�����'��*ܺ���a����᝺0x�d����*��̮��K+d
X��k��.7F���f�Re+a�jn�U�O��F�/5�Z.E+� ��xV}K/�(�Z�"6�z�]]TP}�?���C>������a0���1הe������a���0���J( 
W����3�b���y�A�i���5�?��@��ä�n=�"S�R��f�sAO�Cka42Q�A�J�PcmC�}f2颊:�]-
��,o����ي��3d�ue�R���uJ�F�V����M��)��w��`va�'�Ohmm`��1ұ�t��Fss��V��5q������SKlD��e��]�~���w�K���Bl[j�$Sy
5��b\K2|���-MV=�[W�Y|���T����,��.��!�	�������Z�b���+.��'��j�ԉ������_��������O�'�����l�a�So�b��>.^~���U���'�����m!���P!W���T�FVT�
mM~%V�*�t�"�n�Y��#��U�5t�䪟���s/Q�m)�sl���ȡ��?,?�>�,��n�n޼���,G�ܹ�<}���ib�
�p3�J�|>����r�J)AS��#��Z[^giy��Q�P�aگa^%X*b�>�k��v�����N��O~'%�
���\��|[:Z5�]Zdk�5ϟR�haS5�Y���arw�4tG� ��.�~7�R���vΝczf��Ϧ������A�=z��{w9x`����e7?\{��̪Z�L�<�-^:�t�Iu�l�lr%�dx~2���r�����GG���&���I�n�X�j-�dj�{Og��SВo)�T�=�b���K9��P�q��G����p��#F�����Its��W/)eJ�����z}���_��s����ga1Ʌ�T��(��_�GNɊeS��彷��ʱ�aec��X��x�\ɊY;��9���gi=���:�5`�aP���e���V�=�j�S�fN�����#��ċ;WX}|���T���Nu��M�6r k/�P�r�ޞF>x��l,���u�r��>%�ݻ�P��v��x�~��/f0�B�*������V=4�;#���K�dN���[P��g|�]#}x��F��A/�6,�V��\��Ds
)�n�(��v��gC�Y��mZl|��A*��lo'�ݯ�`O����?���#�w�����׬lf���o�&R�<t������t��ݧ`���q8�p�mU̕,&#����kW��[��k1��l�Һq��Y�N��S��WڰX�Dix�q���TpH�d%��$���ȱg�bd����_<f��#*���^P�-+a�&po#��=4����*6�Flb��Ȧ��!��P�r>o�+�E��I}H$W�K������G9wt���w�85���{�.2�?i���3x�-\�~�م5z��y��̥"��Ӛ��T�j��K�l�ʍ'lF2��M��gS����qڥW0B)�Ɓ�~��=�{�Ə���zt�>vhB�*���u:|���<�|ɋ�m���ی�����y�$�śs�L~����U�u�\:3�=&>8��&��R���a��73�T��n��']|�l���%R���؝
%y﫸|�p�]��RY��e%S����W+�OàdN{�;��J��^z��{����fv��rJ�~y�G�h��
��?Bk[�|�Db�Y�v�f֬llH�H}k��~�R��v�>#OW_{ڈlE�~��UU6lN?JSt��w��^]���>>��l���~�D�69l�vɗ�|y��f�E9��R�h��`�R#a���G�q��</���{B'G���9�\�EW� ]��<y9[�����#=��ӧ��zs��Oְ�UA.�8-�b��n2>��G���P�"��e�����|{U��F�F��c���)eO\	�@��.^��Lks�0.I��2Vʿ�f�ZH���M>9�8������u��'wtt�����apu5B� '���v�ii&�&_Hc&��vb��C<�ene���};p�,ĄB�����,�|��~�=|�?033EFH�V흝����)��j���J�����.�]�����R�\������=ɬ���_����B�Ĳ��i5��(ĶYɥ9�w��Aw�-�zz���OO�v���?2����~��P/�%�,��app�3gv07_�Ɲ��=1awt/�2YX�
Q�>���N����D�X�O�Xވ�p{tQ&�T�ݩ����d �vR�E��H�*���:U�ӂT+�BN�����`3�D��׮�����7fT�e���@'ݻ��4���Պ���D-EJ�u��$��@��0��+���$%Tm�v���̖V���߇�nfuyS/�6�cU+��5+�{z~�WSӸ=.�ߥE��딌����(9������K���ɰ���5#��ܒi�&�vs�x��6y�����88����:��?��o��;y�|����eR���44y��h���4�p&�dQg���\=�k�]~
9CU[r��3=�����L&��l�(yQQ�$K*5�¬.���I%�&f9�,P,�e�L�T���#Q���oy���6Q��P�UKc�q�Z�X4K�|ȩ��.�����;S_ �Z$έ{q:]��탤bS3�� �n�DK���`�p����Z��.�f�j�}�z�|����0�;Z�EbD#1�.�#Zp�<8<A�f7YZٮW���H��OP�h����^k�#��Tͻ��)����    IDAT�Fw�`�D?��=��䔺�N�:L4Qajz�d|������ff1«����\ N9�1GQ gv���ﶒ��0�t�`;Ub-V����n�AP��t��V��V�y#k���G��;�ZU�S�àX�k��f�6�ԲU+�p�^ ,@ӿ��&�{	a*Uؿw�'�y��%s��۽�����?^"��r��^FF:5|��W���N�C��p�tj�et��d�B�*R���v���m6���3�ga�h?�]���0�,{%���fx�|��ӫ؝!-�i�\*����+RH,3�◟ ���/�+��DsEߟ����m&���=ܸ�ɧOix�ŧ�a�z�pi���8N��PϤ0V�~��lf��v?��p~��\2����3���o��O��\2�ԫ��P|�u�֛�7�-�
L�z�Pp��,�k�v�ׇ��%6������
k��qL5Q�H�{+C��t��p��Bb�����>8@[[=�&��T"���71
Y��~�v�kw�y�|�l��_�֐�3�G,�Α+�G��K�wt`w5r��3�������w�K�8;E2����(̣�WS���KI�x,bX�sL}��ȧ���|����T���N35��G��[ķ71W-����c������6�u�ɧ������_�b#��f�)	W3��*RQ��n0���G�Fզ��n���d���y�YS��嚣���!_���	4�v�T�P(��z��X�d�V�P6U�5�ZJ���~b����u�>n�+�G�A�	�c��D}M�d�Y�
G21�LPµe���\�z�D"ͻ�����[�|��HΠf�+���ݺ��u�^������C�~�����g�so�e3s��5֗1��*8�`�_��?R5���_�K�B�E��JX^2z� =��M����^�>\�Ƶ�$�y>��������]����G���'��p�˗oQ+�nj����m��_f�`�@2>�53>���R��l�ԑ!J��Sv��\�ĝ��a�������YCz@�r"VC�1��SJص�V&�{%�$��ݩ�@*W䝩�qX��ꢘK1��!K�)o�_|I5��I��bw�5���CC���\�f�@��&�S��5�(u:�����v�����#����4�ֿY�ݣ{�=�BK�l��!x��bU~�����r�*e����c���y�ZM�n�Cdi.�x���.O&�Kk%Y�l� �Q�lRL����a�>=Ɵ����5��ȥ�
�9�oN��tf�b�O9|��d�I�����$�H��_xJ����D_�\*��,!�s|����Z1[���ݬnE�~瑪����,̰��E� ��d���aP.f�^�QZ���N��3�_[[YD�]
7Xx��թ�l�<$5����F�{zy�z�Dܠm�*���­���U'��$�Ԇ~G�@�֬8�x��[�0b�okk�H�Y^X!�L�3r�|n�v��� �'C���3Q(�X�2s��S�7�Ԫ���1�������q��U�
��$��e+��S�:s�Y%�S-��JG�طk�M�����3����v����`k3���n����Tm����c��hePds���0���a^�$�p}��ɫ�M%Ӊ��n&��3����Nb�%���v����Z�?��<��=|��^UMV�b��ňgJlE��;,p�];9���zzIr3�\-E�E��K&�Ђ�ְ���y~�"��nQ�nc���1ԧ���M�xq�Mt�0�\�M[�Ժh1��DV4_�s	���-�fÐ��R#��Mkc+�@X�Ă(��#}�n���yf)H�TU�g{W�KQ�\�ʦ@����Ys$�I���=u{W����dY�����	)�L2�e^��F6��R�ݓ�	��x�V,�����@G�K���DL�1mx69���D2[�|؇��X�s��;T�ӵ&�t2ʣF�fi(F9{|��v?�|kզ�D�ĵ�OYۊ��եw�TJ�<*⌒�+%S�j�]/�&驕;�(Nf�R���v�"�(⵺�5cJx|���|GvC2���m`tѻ�8�;vR����O{k.K	K9����VN)��bwbu�V��B��aJ��؊�I]�ggdhj���ҾV�ׁ�cW�Y:Sda1��²�B�b���Vښ�
��{� O*�#�4x9�J�lQ��TwHTCr�f��rp��Ԍ4����5����g�ɤK$���5��O&ty"ߕ��%LVɍ�g!Ů���4�dr���m}Z4�a�a�a��0��g�7HŐ��N� �Lܼ�����i�I&���W�&��v�H9�V3+�W��J^���7b�Oà��E���C1np��oy(�`l�Y�#&*� ��n�F�	�R��2�BC������`����v/�Mr�W�K���������~6V����C�"P*���6�k���,�_<W%L�jn��=��+u���z?vl?!�>eq~V��2��x��>^N%y=������D��R�{�e9�,I͙����'��|0I�����ʉc�<�7ëg���`���W3L�-����=�w��ָ}��f�%;)`!J�U������4mȇUɟf�y��o����FD�bA-�%������ך�HfPD	����aP��Z�a��6Q��$���^�J�ۃ�����l��tc1�8x����p�U�8���U��g��Vu�����=V���!��oU�?�=C,��l�����>L.o��glln�w�0G0��%+�+�e��,��So��7��_��D���.$-�U�f���e9�ʑ};8�� w�N���;
�����T'��_}���*��}�����;,/�P�&y��	N��ʵ�=Y�lq醫,`�]��R1Js���o��g���M�A<[���&wO���	��|�n?�7Z�p봟�B!�ݱ�֬\ԍ�ȷ:(�j�u�kilm�͙i6&��_��VX�a�\UIz�$��L��	��cx�;�5�)e�q�24�M������D����*33s�V&����Zx1�H�bRx1�a����>��������
���GN���=ܼ7ǥ˷擏�����+�6�	��j��5����\����lT-��ȁ�u�B���q[-��k��6��';��O���ڕ�/�Aw��/4����X�(s��3}X%�|p�4ǎu��w�<����m�bvj�nQ�{b[w5���:�Ky�A���kB���\ɸ�\�s�A�8d��7��?J	�T��+��DWh�Q�6R�@UL�Z����b+�apE���փH6�\4�0z�ΝG0����7�Z����P_+�^*%+3�K�~=������-�ֈ���>U$���ɽ��x���lmn��ű�*t�vp�ݳĒ&.�x�B��P� !��N;�'��.�] !�}@4S����D�b�qP��*�[�kf��b#��玲w�/�tG/}�t��q�@7��ܾ�������ꝙz�ybO:��P�?���6Us S�E����L9���H'o���hx���m��p2�����饿�_K����G �@���p��t��0h�v�V;΄���SM�+=�]�r)f�=`q��IS�؜VA�b
4��M�g7������%�����z;}�&<N�HJ/�F��˖/�CYrb������Z����Y����i�ʘ����(��i�� �p�A����T��K�"�+��a%e�Hf+�
��͊��Q;�f�PN�2x��(���/o���T;��>nk����gb�_չ{��Z�fa�PhU,a�$�x�-��<W�P���0"��N:b5O�Q��᝴��X�Y��F��In�}�v�_����BM�M׶R̭��L:$I	�d"�XW��$I��b
c�bި���M|3F���yF���=:n�:���k����M��]����44���m/�
zq����f�C�v�|�gO����M�M{{{�1<V)���A4S$Q��z���a�1��cca�ٍ!�]�С>]*aq4g�	���Y��[x_Q�XLPLoh6��������H$U!n&��Ʊ�.��A<]#_�q��,��k�D�����u�h
���T��4g�"���V,t���Dv�jˤ�V�xy1��w?^�����tTՙR�J._Q'����K[bn��p��\�4b�3��X
�%��d%&O�/��V��6֦��2���&��&�����d�E��(��8{�;��A2����Z�c�n-��`������]W���e�̸�j��
�LKǡ�G�Y�$^��@G�]�m;E~v�[\�p���x� hVe������eHL��rM�X�N����.�M��,�ϪMBI�1�WoRZ�>�91J�`����U�E�ؗ����j���4;;��Y�@�ԛk-ػg�
:9���������)>�"�D�wO�a��G%��Ȗ��3�o�%�αo�>BA�d���uҹ�b�\�L��&J��EE�Ֆ
��H��ʰ�Vt�����W��`f}Z!y�Y�x�:���0l\?mo���� ��BgHѪn����\nZ+
�{=���_H�-]�a|>3����t���Kr^x5n���w��=�^R��bԫ�Ok_*AdI�Y��t�ׇA�E{�|�KY�w����Ǜϵ�'�(�ND��g��ϩ����Ss��YzI�&I��^���T����Y��u�#$Q)�ٿ�������l��2x��cV7��� ��Ar�*�+�ǍjpR�jD�*�rE�M��J��V�ԕ��dź_���Q�&���wcKXLy�!V]a�]�����F���a��QE��u�"K��ߥ�%���]�@�d�TUW�9��&b��D"�7}�5�>�;���<~�Bk�Cc����:�\Ry&j�wx75�z&�.1,N�W݁(�kY	ָ\�Y.���Ȟ]m,-Gy�z��a���?1@z#���
M���Y،R(I&��>vd?.��kן�VXU��]�j�(�D����o�&���[�Z�19�E�$5`n��	�����B2�+��$�&]��=D�.�-R�bRI���*�[S����Z�"e�>�B�9	�Cx\j�����./m�ķ�,�.���J0��; U;�뛤r�RK(|��Ξ���ܸ~AQ���[x��475����Y^^�퓇9z��k�n1??�>`���n�}�>�����IJ�P�$9�RH+am[��S�a*l������?ė_���r����{�li���k�/-��ǟ�;���[$�4�T����_��s���R�aw���P��0�s�`���a{S)��k����b��.�"W����B<�ѭ�`ܥ���+�"�M�t@dr7��P!���Iz��E��6R�<�;���l�Ͱ�r���kj��2(�A�'�CK���]g���akh��R��Z`s�9�_�A\<�s��j7���k�Y��	6jNdc��������2K�:�Jo��uZ��5�w����k��#��M���1�h�N.avoK���-�5�9�cCfg	���T�ᱚ0���ݽ�����򕧼x���	C��v�p��}|� �`+Ӌ[DSn��ht���|��.nݜ����8}����ʥ�-��t����?=�)H7�d�����9��~L[��:�l��ڎ�-�Het��/�&���®	̓j8�ރ)�z	`�Q(��b-Gk[����&�����9L��ؚM����C�M���/^�E#B!�Z���SM�D���y鎑��@e���<L�4g��2����BJ�K����!.>]gzv�L��6���.v�hѵY�O�~Z�l%ܺ��6��A?+B�u��E}�q-lQ6"|�������O��Wds5LN/�[�L��� ��l�a3c���yy�/�����Ü:3ȃ�K\}��5�������t%���h6��˨:#ú�����$���?���ͤ�E�L�rJ@�ٜzYj�|�զ+�m��|�(`�ډLUUł)6����X��O%�PE�p�1{|X�-�:w�څ�aoX�p�©�;r��b�D!e!�uc�V)Vs���������^���&�h�cG�oOF"���$+K�jՖ��F���Al���.Ģ���.�����ek}�h,��V�\����څ����>�>Kv���+�Z)�4��sh�C���_�i������v󳳇p;�<}$��MN�{[;���͡Jn�fd���	�}q�%�OUdQ%kT*[5��V惷r��"#�GrH�S9���X���N����bs�ȗM�^����:[	 ��`�L��c����j��7r�pr���(�p�43��MT2���g�e�j���0�h܃��gc���/�;y���tu;��ZB�W�XX�$��J$Y�b1�������o=�fw�������
���?Glu#[`m+A�b��،�Qz5�t�x��G;�V6��b9%B����Q���i�bq���R0��,��ƛ��@!қ|pr��C~��+��B���r��A����{����w>�
���'$��>{����_��fr��o�)E:+1��I�Z�L��� �|g��L9�����p�|a�K�������{.(zy}D�z9���Wd� �r(�KN?�<KU�ņ���(	ѰJ2��)ܤ�A�;Le"�u\~p�JzG����AV)W�؛��u[�{�I�AHe��ީ.:Bfd/0��$�5�~W��Q�B�/V�qwR���N-~3��>R��3	2B$,䥊��X�hl�|}KS�#'��F"�n*_�O�U�l�(Xy��⚕aP�K�(}���'��W*�,vb�(A����vښ�y"b���u&_�c��gx� �������K�LN-kv��`�9U-1����}t7CL�F����x����)����N��!���d�h�`-�f3�'UCz$Ŷ�	gMr�V,6�ރ�9�2��jRs�Bg���׮����d�f�V������h�{�1�w�Mԁ3PW��2mA��B�v����O���8ȗ�ZY�gio�K|���f������Bf�"�l�"��ģiҙfk �۫�A0�b�����J)�%���D5˷�&�x�G�,ǚ\�%� vE��ʹR�R��������W����VQWk3���
�Ʒu������f�SkJ�����7q�� 3�?�����'�y���e8�g��� �t�G��f
5���˫�L�`��Ys�FI�5��E�6�$�RXo�.�X��:9꽉��{�օ�,���>~Ã��R�.b6�t����o�^|M�p��ުà�V�c-jN]�ֆ`���J��jQJ��M����\�Z���4�t���l��'�D�J�0TE�Y���b:[�������P��}�R9$�c�����҅�n7�dh��)W	��F�H�*��;2@o����YX�`T�7MgK�&��,�\^���xC��m�J%8y��Mnn�|A.'�s�������X�c��o��&�G��ʺ����|L�A���4�{$��U�LQ�˟�Ac�O?��TK������4R�v����U�,6����+�����͈��UƖ��]6-6�z�k��Ҵ����xܽ.�ك�]"�\ӌ`�d����u������IV����ɡ�;���(�ld3f� k	~��@I�r	����Q6��J��=�o?=���?��oq�]�o�0>�G:!�L�?�����V���,��R����}J57��dK6����pb6K�e����OO��o��(U��������:_���&����N����?��z�}B.�2�I�<�-h����(JX6VV���l���T����������9"���ZzE-����\K�������Ή��{wa	5�
��}DsЊ˖��U7��)V4*ZN-@�o�C̨��N�4��K���R�����Ck�\��n�l�x�ʓ���lJ��df�*���:�l6㬯S���N���z�Lѡ�hQ�J�7%�yPHO�Ɋ�h`$W9��~l�O���JR��|.�d��>�t(r���&O��)�� )�s1�Z=���Gx�z��/ޢf�~3�^%�(8�Bl��V/���Y���cz��d��~����^�{o�L����z���8��������o�n��D,i�Z�\S
��\��mi�*�����'����{יx���?[    IDAT�,&ٞ	�&�c��zZ���C�U�uc��Ք�H'/Ÿ����^�KFgz=�V������l��5���W�^S��]2�&6�Y�Sy�7sZL-��>�����<�
U�D-Kf�DS����KN�s�Z2$O {B�ǘjI~�4]���N� Yy#��@��L�ҹ����r���~�$m+$�����p'���s��k�ָL~�+��e���6�w�s�x?FZ(�U��"�xr�?��kv���W�:L*m�(Z،�]�`qs��QF���b�@EE�f�A��Y7�b-K�'��N /����W�{|sjM2��C蛡ܭ��w��3Ac�nݼ
j�$a_��6��Y��ˌ��wO0?��wP��ġ#�����gĒf6�I%�?2N[��P�(o���X[�b+�f#nhV2mTذ��O[����
�J����Vf�6��w;�'�j���dq+M�brԍ쥴���?����=���GR�*_i����?]Z��O����ퟝ�����.%0WkX*>}���N������W���T3y��k%Ud>z� �N*B�4�=a��4.�P�Ư�1�-������<v^̥���;ڱ��T1��	�h��o�*@�:XF�{��e(hG{s+n;,�~Jt��VKl?�N{_;Gwr��r9}�NP��bk�{p�b�*��ʥ�G!�"��D���P7k�1������x90���E^�Gȕ�����N����}]8�f���<*�]K�pv��a��ȅ3�۔e�����'0��aR�g�F����6�kQ�7�j3˳�j�|C�'Oj�s'�	���z�x�T_�����vٸu�_����~�[v�|���-=��^+���ɴ�//>cm;O��}�����!r�(�A;?k����Y);�,ǒ����d���U7F!����av�x1����'d�5���V���7��t��U�v�D��/�6Y��2��H�/h�l��U*�(�� �c�Z�0#����������v�kj�PL�9���NQ��4��5�ښhjke5�A�P I��;D���ֽ�,o%�����aNh �ȑI昝_��T���Q-��ۈ�e����=��UJ���8��,���(Qs����)V����)�	�^��+���|��n�׳\����3�����l�Y^[��`����/fWU5�^2�q�u���
O^̑�X���10L�C��K�q|� �}MT��f��v)ϜK�oK�9~�0�]�"1�v�(�k̯�x�|C�-f�j	�݁�j�gG�Vw	�M�ۤsY�5�J�N�ӧr<�|���.�ۜ�ZI��^�n�.z���i`��U�%�tH��V�m��sV	�*�)�Y��=���n�ᣧZ?$���G���~�;�j�wX�|^M͍
�xQÒIC���T�x&��n�3�!�`|� 投D"��eam3�J��v�dN�-~�B��!YJ�S���4+�82�KO���.?R��!����=�z�{�3s��l��s�g�����>����!	� �I�")Qޛ������؈�ދ����ec�g��T%�TE�{�$��{��4;Ɥ�P�F�4��;�{�s����=�R��(8\�Ό�����*�o���g��U1�j*)�88ŮA7��_$�dP��O�X\^b��$;z-T���T[<{���V
�ͫ�s�������J8��B�V�c��?���.�l����r��O��e��hZ������G�l%
����b�0>d�ˀS�a���=�ϩ:(ɀ����Q)�XX�*�e!�#�4��
�P�e� �dDE<�&2Z1�m�Y��(p6Q�?��N6[��0����CKgS��8�$�ِ�q� i�X�"G�N(j��;�H��Z���m�pO;.��f]`=9淶(J׵,`�E�L�b�����j8!=ǒєŊ8J�vj76�;�E�ό������]�\M�h~S�s�L���D!U�T+�-�.�]���;.}�;"4|1C��3A�����݆�1X���'�rdh9pڽ*+�qY	MT�,�dB�$J�|adS�۔�>��+ѧ�[T�G&5�>���a���;4�:"���@�w���Yf�'H0`U埪�b!�m��TX	gHe�X�^�'�7�\^:��4�&5�ohY��-~��A��&����!�e�h����׏��"S1q���Q<.?�N��9����n��p�LQ�%���jd���B.JO�Η���i�S�$�����d1�7?������_�)s0R�"K�1�"+�q�2�6���o�T֨TŢ"�;�	J���ji�
ת�hW��K+�?1��-��l9�9z�8�{`7�`��׳4vwr�@�ZOKA��F�D<I(��3)D}Kg'[Ҹ|{�p$�V�c��X�e2�5��5�D:[SV��f���O�����s<H�� YG˖��"%�,�n�q���rwnOud�d6*+���F+�jQuӼ{� ����7وK^ª�k����몐I0�;YX�p�Ɋ��	R�i��=I$�����(7��L���_��6Q��5�]'���ʈ��n>|��.19���?>��!��J��T�Ka֣U���ɴS6b6����45mԛ�ʒڪ�0ɥX'��*,��b�bp���2z3��혡mt/��A�ҥ�o�q[��I:��Xu����0�a��)K���q��+�#�z8���Ĩ�1��g�����cJ�4�tVeT2�*z����Ѯ���������� 'u�<�T���M���baT[s�� @��R�l���	u�O><*�{~���`t�,�⭣��?xL$�g��A�ř{��]�Q�3:��G�Ns�Y�������a�\V��)E��-�:6@�P� �t���̽�������a>������M6������������zJ9������Wv`�T�xhP�V�fP�����xq�2�\�blI��V���߆=ԋ�3�W:#{�0Z�XmbL�,���\L"�O���Oq��~�x	��̩�?d|j���ɺ�8�RV��i೏Ϩl�Xi�z�	I��'d�\�����(�lb&^��081AG��jMǽfg� 6���Mv-�zKYG,�ЊaN��ȡ ��p�D�D>S�c��믎�Xy�t���w9q�-��ߝ�C*+�b#�V�_}zP.���W(7-ʺ��xĒ+{v��6r|��a��Vꕒ�2卥�\�rS�><y��?�jFٝ�^�9�^�O�h���}�������D��RUE�8ۡ���u���Ul�����!ѕ$W�p���^&w�V��|I��#4!̡!z�w
e/��$�/�r6Ɖ��9~����]�>�Z8�����$���x!B2_Q��|&�`��/�s������n�}d�q���8-�Ll}�������1��4m���	R7�v/�`@ɘ�|����v �r
�������r��ﱶ�V������8n+�/_�zq�}G�S7Y���u2�
Z�L(��O�M48wm��dEY�EmH���Q)$��Y���N�./ћ�-¹���K��ן���j���*�g��y�\T�T�L::C�\g~�5�bYe�d�V�dB�CoE�r���&����d7yx�g�E���}�&*Y.)��7��Av���;���{ H���b�B!N��H+����r��~��'���1O��)Љg�s������U��"m�ѥ�3=>�`�lA�Mf�\�h*�F8��7�tt]���\�+�`�eP[��x�Wk	�U�K{��P���2�j��#�lM��C6����9,7&�������"s���L����&7�=Q�!��sA�c�lEu�eӂU��)C�f>���A�GBh�
��V/W����K�9t`��ސ����l6�׸r�!�^��hҽ*"�&��`4�̫��Iƺ�6�b�n�����w���B9��A�`�L�� _}��	MR6Y�{��vw��j;E��uꕔ���<>�8�?��ʥl���y��h��;涫E*Ť����EwO᭨����٠c5����:�R�R>�6wR�&[qq��N�z�z<]W����)�E�/�`D�'V�䔳��GO���7K�Ѫ�p��ɝ�v����llE8��[kv.]{�� l^�����m�x��5Fc�n��'T�B��&�9袜�T�l5��'/^2��5�g�(1(�A���0I2���Rb��g�&&M�_}NE5�sR��ҤP���z�AG0���p��/ܻ���
&cU��kF_/���z��x�~zzXe�;����gj�X�4�}X��JD���bua2:�{o�xJe+,�<�h�D>�R�P���Dl�n�	�
���\rKQ?�P.�/�Zz9k�
)�~�PFI�-��VKa�8:3I���֭��j.EI*�]�-z�[Q����d�:O)V��&�Cm��`�U����V��K�!�V���
)}f��^����8���d�{/V�5uLO�"���$~�'����4�Qe�ّzX*V ��RI*����:�w^'�2�������V=�f��ӇV1�sն�a3���;Fd%�Q*�)��-�(�	�UD]�7�����d�-���.��&�B�J�B^6p�����Ń,����vވS*�'R�#�N�I�$,���Q ��P��8!n2���V���i��/�����i��ޜ�����ik*;���t+��,�2\�K|��{�:�����*+b���T�K����[t8���>��zꅔ�f�>����XN~��;8�D�nPE��|��'�S�V%���i�o��%=J6je��	uK¾b1�Z��PPٱ�V֔��zN~}�Vq]��� �hY�i��$ή>Lp����Nv�9д�t�p8���`���9���tv��U^̭�m��e��c{�iw����|.�:�j3��,�*����;u�}j��ظ�سP&�^����\�����Z)S{�1���-�;%� �\b�9�->x��~��w���W���ϙ���&޽ã������x���{�4�g��5����pF�l���Y̓��.Xs��L�f��'oM��� e5q6:<\����|���q>}�8n�o�g7PBϭGk�{<�]_ ӜJU�g��T(Wh�ʲ%YIC���.W�����MF��߻��ԥt^6��I5;��hE� :�x�x=V��젷C~~�D,���}A��������r���R�۰M��fנ�l���[Q5�
�s�����$�Ѭ��3��b��K_�M>Q��˓-VXLf�����-�5���=B.f�a'�M�chf�u|��>e��ÿ�	��A��g����Ҩq��x�ė��'�N7���y�i������W��}�/�����A�Q�~��84���o��K��/�h��lFҜ;���A>���JSU��|V�fWfW���]�.����)��5%d�k�WHb2E۶<n�y��c�5��{�g7/�H�R�-�*�A���8:��ً�s���i�r�k),f���65����N��{��3���u��ߐ˗��/�wd��}{�׫I�� �z���k:|V>���i,������N6��H ^�G�����5>��4�k�4��LV=�D��b<{������
А�z��F}��N9����ݼ��?�{���5X�|��A�����8}n�\���,� �l^m��<M�h囟�
��U*!d
�� ��z]-�g���͊V�}mS��	b_
���q��� �ZZ�A�/��?_��n0�ŗ�G�<}��|���槦�P�)��ed��h)����{;�T%���C⫯H�>%v�:#}�9�N����7�ף�R�Șh5K�dk�q��c����O����d9q�$�������ҽT�lXIv����3o�\��Kg�=����BN?_]��܂h5�Y�:���Ӹ�z�E�W0b��Y���g�,��Й����I����i�i5+�2�:�S�1��\����h��x��n|VЪR�"��o�����P���e�꫓,,�2�B"�����mxil�U>�7`竷v��X�� h"c�2�����3x�f�ٴ�l�^�����D����ޛAk�T����:�b���\�AM`v��%��h�T?eb�%����ʽk4
q<m^v�&�ɳ���Y����؇�g�P?v_�R=�ݤ�x����T��s�9~l?ã}���[�n�o4��p����x�2�h���~����۷GAnd384�C��#f,��R��'Yfd��wO"����l�w`�]V^����`�p��N�m
DW����mT*�>{����(
�T�EW�$�I5A��\�y���!vO�2�p�X���nG���ݴln%|Dp��rS��-z#�z�F!ơ�a��iT$o�ݻ+}fWn�c+�`��i���U�H0jV��X��U����0:sSU�����
��T�H�W¶�:�JQ����hf
ܿ|Q�DK�e�,�F�.�uг�(mC�T�v\>?}B�4��QRbPO���E����[��ǯy|�	����|c�J�̣��P�|
�^V;e�C�@�HF��|�mZ�˥(˛	2�F}�����}X-B�n(���|�ų�[lDRj �l	�ф�fW��R�DPUr������ǋ�nD���vy��(n����MU���{��|X����2;F�����ɳ/^�a���tR�j3(H}-�љ]u9���*�-%��R]�3{��͠�2��h+6Z�}�D��NML�-��f�T�A�,x#M9���"+�6QU�՝m���e%g�O-���P�!IG ����������D�`wOPu=��U�mz�@)�R���]cjU�?��=���o����W	�
J�t�������Q���T��XBY��M3�tYU		���Ko��B.G��T�l��lΙ\]}F�&���֠ڨ�ڦ���Q���.:ڜܸ�tF�t��K<<BWl���m����!�y�j�Be���������r���U尲�}��@�Ӓ� ���>�{K�`�+�V����K��M�L�TUL�Z��L^��z%�����LF5��� �*���$�eۆ�(X��"!^���)b��jI���<ސ�;�yڰ[�T+9v��fr�C�T�L<���_-��p`wz�z��.���}~N�1�Y_&+��b�|�J<�Q�ɺ�N�8i�
rhf �䯌��BF9�ΰN��I�X�aE0ץ~AG�b�e�PjiT+)}��O����R���:�<���>7�+��t�w���=fŘ�}���L�/����'�|wIQ(-v��
o!p�r!��]wj���y5�k�]̯����e4���p�Lj�+�ź���K�~�����eT�\��k�k��	��P�t�uM_y󪴵��ZLDV�H�bp��F���)�Ġwh���.;�RFy�[�tB��&3o;L��b��Mҩ4��N>��-.����e�B�jV���qt�BD/.n��%�ϲϱ.N�)ɥ%h����M��[���i��$�q���k�N?u������J�r�V��F�����CLM��7�X��U>T�f_|8C�n�ƥ�ܹu�Ͼ�-��n���!������L��x�\��~8O�*ۯNj��v���F:$W%b���YV�v�����Ξ���a�>��P���`pY�|�5��<�����`;�h�j���b�P��0���^�a{�@#Z�J���Om�0��X|x��l�R�n�ر���)�=C�&*�W�֋)��RRQ͎?Ǝ�������#e_��˯)h&.�|@�fP4]���L13���L���v.���l����u�Ջ�JQ�����#D7��E`hl]�ēe��w����+ڥ<��iuک�0� ��4Vc��?<��i�������Jp}ǎ>�zwK�����o�y��3
����tH����W��u?ʅ�/i*waS��M�`.���!��G+o�`D"q�5�\��~��;x���J,�˒+u�����p�.=�#������x�bMr{fe�R�P�(1�� p�|���.������{���+J[�*q0Աw��������>JG�^���Pɤ�p��tmڻ�ѡn�N������yr�#�������FZ��6�wy���=։Ѭ#�o���!K+�`"S _���ws`j��6}җ���j�H���j�x�H!/X�ZjS�|b5��v��WSr�E��\b����8�     IDATo����[\�x��P������@_�� ��[�������Jfz�w�L�����7Y]m��wф�+�:9��NK+Ъd��������\�j`�F���˷�E�|p��=Ajմ:ׅ긲U���3��w�TY�\"��Uk�e�8]��I"���AG{ �IWgm� *@տ)��
�Ň�g�00үJ�/^�M�b``� zW��NE�o�Ǫ����g�x�C~6F�T���KD#if�'��,\���'��-�x�t�\���3����Tu(�śψW!Q����EO7GgF0��ck^-���w+�S�I�C:��$yt�K��9��*��"W�9���'y�"ɕkwUՎ�&#m6vt��jW0���(��x�\]G��0[��L����q��7�)5�꿕��t$?ߨd�ks�w&񊷴TP����N�PUY&ܿ��=�#�\��%[E����|����w��B2Y����";�^JM���љ%ja@�h��$6�΀���K�\?���*���2�k�X<��f�j���`hr�m=X�~�Z������R���n&����p)(ċ�?�=��l��?�`s������O�U�R�đ�nf���l5P��Q�[��u�lQ���l܍v��qx7�|U9$��戤4�#E
e�g�vB$�A=���Z,$1�
x�N�Qg�/�o���0���Α ��X�Ӫ: N���"��n!P)�L(�wU�VM�V|"[���U�8'G�3�Q�c0��K $&��|��fX9vu�,��K-&;�x�7f��ȱ}�=F^�Ze+YB�ey.iқ(w ����kRQb����f����ܻ�3����XӋ`s�s��8B��u��?@Og'6�-%}����@�_���ZI}^d�$��`��vK+9�̭���0Z���%0���êZ��:�EtȳA�q�s:��F�C�{ʕ�*���fJ	�t�����o4��.U��$��)&F�����O^(�hG��@�����ۮ��ssK�Zؠ֒,��b)˾ӌ�
p��+�)u��a�d�k����V��Sc
�U��)�ܦ�ȳ�<{:������3��:F��R�ŵ�w���ؑ#t���2�E��R⠒��KTmASh��F���`�t����1{�;j�%��&� ������}�F���xۂtu�ѷ�8����NT�!���`��q�ؚ��K*c|l�S�x:e3��)��jS���i����])Uj���1�D�ϭR,4)E���bzj�R>��b���b4��^(�y�Ӱђ��\�hP���*��
c�=�y�x���2�@��Ω��*����sjZ�;w/�x�r^�U-V���L���V����8\�&|���j����7`�"5Z�w�H�Ľ�
�3�{�΀�V����>�_N����=Ғ�L�(TD�
�DFE]���#��*f����gK
�[*��ZI��"Q⎹�ݮ'���jgblD��?{6G4e`���3\��D�h-v����\zz;]L�݅�b$�)k��,"�r~�tZ��F,�����G�ԗ�X-�����\.����D}ӌ�)�����F�l�(v�j�A���}��Kp��C�:'�Z����C�^mr��y�]���	���b��\N�b��>y��n�}I�^��!���t����՛���eԯ[��E3���O�:��ˏq���\Q�n�&�>]��K7i�$��A<�"��*|�XJ�R���������74�����j"���?�ɿ�D-� 5c;��N�͠)���LK�)�R欃�� �wJ�1����W�}C;����8s��+�R�j.��
��I�N�^ͳ{�4�6���_���p�ҏ�I��X4>y�M:<[[�����R�����:ϟo`����tJ���Km�jZ!������=:���g�d1��ԝ~_8C�����H��Mΰ׸x�9��M�h�����cē%�=w�l�K������Ţ�QMG9�����VYN?��p���?�>S}�NYo��u����\��=�Ձ]O��z�\�L����mS �R���l��؆�l�A��J޽������h۱w�N�tC
 #YO��FW/��
�C��1�� ������G8���?�'j�ku�يXŶ�r�}��$o�fye�H2�����A74��x��r1/�י���ӧ��?S�gdK�ţU��7���*(PKHiba0����hlR/'�53���'���r^M���c���	��h��M�l�փ^.����R>����}4�՛��x����Q)5F�a��I6��=C�{��z��&��x��f"�(r��UE/}���r�ʌ��;��~����o1�k7�O�#�0��9�\��fDgv��z/H��*/�X(������Cta���W)l��_�U������_]6��.��!B�ӊ�Y(��kI����~z�-�VK��$ ��?;�����ڶ�<_�s��=�5��O���!7:���j�x"�~�Օ0�l	�;�h��r��v�ݏˮce!Bx+��z�B�E./. ��135Y/���Bi[�u�ҷ�j�WH���3�O�H���۟���6&�~���{����D�1<{I8^R�L6C__2ɽ�InܟG���AS ':���i�r���'��Ѭ�Դ�f���jJ��#Q��M������1�.�_��n���f����XZ�s��K6���ʢ�]�,t������1X���\{�ڭ���ntx�ܢ���fP�M��{��\�;:�;�=����*�z��!��̔�-Z=��M.\�%�)`�X�51ʁ?��(��l.����ٌ��LhZ]��+d�9<��������Klm������-F���D�!� �F&����ckP�Fy�K�-��"���������0JHړ�!��߃���`1�چO���%_(�n���Ӽ}f��e��/R�M^�P5-�;���B�ޠ�_�;I�l�RI��;�R�����6����^%�M+B�be3V��~����w����X]Os��+�&{�B�m���B9�Tt���$�����ϳ&��|�P_c�G�؊�NP-�0x:�:��g[��_rVy���#�!?3�~L:+����.\>s/W��}���;�%�DK	��;�j���N"UV���E�IE�q�p8���g҇]
ΚF*5�ͭ���)����l��TQT���һ��T+YZ�F��q`�����W�J���ux]f:f:���#I��zH4���oWuC;~�b=ȟMd�c���;� ��U���F��Ѩ�I(3���k������26֩��b���\d�7o�'��s��Q���c%��bDRe�y�L���F6��~*��l~��h
ܽ�w/�H-���K���6��v�7��ѽJ:|~:d������b��I�j`i9�f$J�=��@N���T�كG��ne��t�:��������Y�H��P;�X؜����`?�#��F�ɂ�8'�I�媲*��,v�V�6�O��E<i-�oCCG)e�����}�u�]��Q:��U��:���I��ٌ1����BS��<'O�Io����؊
�E6��.�8���P`��(�]�=��+ǉ8z������=�E�.C�2v�� �]W��7Oc���t���f��h�|YSU]M���)J��l����`��?�����bP�/o3�����A����q�����^Pb�"��ؠ��G__Pu�Efg'��9���C<|eq=�쫊���3ef��Б3�ew�J�D���¦�Q�sC*���ٽ�K��f�I�+*Z�Ս�"�"c��hHlD��V	�͠��;C^�Lv���fn.J�Pg�;ľ�6�&��U�x�6b����덎P���=�,�'x�!����R�a�՘�/hŬ�@�B��}�@�Tbb\X~Z��z��t&V6,.�����p_�l�����d^�4��/!��ŬWbP�=�f�_�`è|���VÊ���߾-H�)���J���c�qh?�B���.������>��Wo/��Ų�3��uc���!>��-�4[���v1>�M2��P��R
�Y[��'�g��Q�h"��� �;��\nq��sW��V��@��+dA�}0��/N�������)/�٩i�:�Ir���zW�������U����J�/�<C��P$�DZ
6=�J�S��R�����BĠK���MN����ϘMz~���8Mz��uz���ѫu����L<���;و�}�\y��%��&(_�X��Sm��B^e�Z^����z��)�Z>��.z����@�	bq�i����"�4�6�� N���=c�j:~��wlm�9|�${����9ֶ��FB��__����Yդ���To�-׸�p��pB��;�-��>�m.7��)�t��B��Y�9�K��(�O�Lz�e0��%1�R��=��o�p��B�K�u���[����ъLV�Wﯰ�����Ϥ�
�����c~!����)�:(�\*�+��bG��Ìu8���I�:�K�U���
�h1��g/����[�	�%L^�b0c���r�9��<`��)N���^Գ4�ƋW�ɔ�][fr�B��u�a���M�[��^gEl��41�w1�=��{W{�j�FS+Ь��;�t���թ.�eMcm}�͵%�@���|N��t���L���&��o�ˁ�^e���jڕ*�U^oy}M��q�s��'�h_�����֢^F#�%sD�u��l�
.SA9�ł�l�$�J�O>8��.g�����&�f�������m��!���r���vmà��U�����9�O����0&g`[��F��W6�Z&���{'�^2�5���n���w�����>|CM֌M���>7�����s��G'A���׬F3lekT���2t:�gU�M��F=��.�Z����xt�J��P��ȇ�����݁f���꣭g���l>FW��7��u���&s/^'q�\LOL�j'䷪�3�6�V1�;�fs;���TH���N>_Vw�ɉ�T�+���Ee_�9Ersm^� �Lf�EUǈ}I���cU�^�z��A�%��2�V�Z!��U����32�O��D<���cfr��K�PR6�]{F�%A膯V�d��L�������-%��ʆ�|E�4iVs4+q�|�$�v��*�Ĳ;�f�JnE"�>u���v4�]6�x�A��2ߟ�N��cz�(3�tmrun=X`vn��=���٦��$Y�Zv��������>��ה�K,�<�Ȏ>��p������CX�8zv`tx�K��ݭ �=F�6�<x��k�c׮1v�Ǥ3�����2�X�Ӈ�lVN�� �X�|&K%_����29i��(�k����8MMFz���,�g�ԍ�l]��js�7ˠ@#�Mau��nb�,��#�:,�vZ-A!�REFƂ���>O�<�#೷���g٤�j5e�
�:���)<��o��ǟ0:�ÿ~���M��QP��2p���rq:��>3I�"7ĊjխV2�?��2�b����na�1�4�V�i�o�����g�R��\�r�&w�.�|)�f�Sh��(6'q����b0��s��\���_X��`.J�� �&��E�ej=���<��w{{���i�<S�O�2�cGW3���k�<~����艣t��:������+���Y�س{��u�_XgY�D]�����>(e�v����nvO����)`�` KOg�9��,R��2P�֕��˛��.6�zMKҬe�ٽ���=<x����:f��J1��@��;��y}�J��fX]�"�+P�4\n7o���J�¥+��+X�/�;yF�R���C{ƙ(;���.[�뷟3�z��gԥZ��Z��"��s��"��<q�ɝA�u����ٌh�lj�&N�QS6K�
��i�ܹx�;~�]����
�l��ϛt��fq*�L{���ClL��
l�EX_��������O�6d��T	��h8T��f�h�Q.���jD�EE͵	aմg1���CV���g^�V%J%��3�Z6�q�d�)IR �l����lU��I�a����ڋ;4��7o�!N���FO����h4��r����� \Y%�N�a�����q��"�*��:��pR�'�j�ji�M��{��d{R�aq8�����������h͚^e�\^�rq]�z���5�9���~4MO8��ɩ���8 4�v��U:ņj�3�A5]Ubp���MTEptu��_��4m���=x��hk�Ш�1i�{w[�l󩳠)"�d"ߢ�������uq�цb7��B~'��V��@PU�������jr�"�f���v�:��}X-z�ጂ��r��vm�&z7&�����Th��٨���b��N��"O�Ш��9mt	 Ќ�c��	+$���庑aQ���>�Fܛ]%˨^⊸-m�;��+͌���b����,��1���lHb�ˤ�]� �d��st��1�s�f�@4�gq#F�.|�j
����A�"�װ5�����C�A�'� 0.G���΄�.�i�0V���ig�?��F����0���I������O�1Z\h��FA�z�� ����v��U5^����b�|���f��df�W��^���b,��Y\͐-m�s�R�-�c�	͠���Rep�*���X��7��XlF�w96݃��VŘu\�u�ŵ-�SUH	�W_��0��������Á��V�L]-I�W�g���7��X�5�]U����j���O�(�J�&�s-��WkQ��?����4�}�_Foܖ��(����CJ��^(�4ܶ�J�[{ȏ�ffsi���2�W�ȯMTl�����{/]��Nbm�Fo3C5GG�I��ׅ��cc=��Rr�dSk
�?�{�����WO�gK*S8=�%���wP�I'K�
���R9)���$�G16��ԀL�@t�Hx3��V��VD f�Gɫz	+7���#.�	-�TL2����fx>���+"�P�2$S��e��8����*B�����#�0����?���9�<|��9L��P���ܬ�SMG����n]c����c��y����/������qBV!�f�Lf������f���ϙS�T�H2Z�ѓW�\ݢb�P3����fh�Q�ⴛ)W3��]l��kJ6��fS�� 8<��o�V��U���/dbj<�P_��P/��He�x�>�ֆ����u�|!˹˳$KF�����yp�\�((�Z:����&Ѵ§�8hQabw?�@Wk�4�"ɑKWx��FYנ$�6C� d�N$�A#TUAH�;]�dt���x��n�s��}��Y���7�S�|��`�5�ד��R?SR��S'�`zo�?~{���6w�`�%�b����'y��A�V�Hɵц��dq1����������D߬�+V	�p*��w����n>��}�8���8/֓$KMՓ%Iă�S�t��v��}���<�r���|��^+b��?D``��������	\��j�Y��Շ�����f��>tM=�xc���hTd6	~;!�� �l�ZU��u1�����E'Z��պ*CM�wU	�ZQ�Nho)R��˄T���q����P"�P�@$4t�-����R1ab����j���˜��.��_}�>�._���V�CG�q����_���g*����ǨV�r�6���`L~F���l"Z�F9��g��A�RUxmAs��.�a#�����1�^��GM9G�����l�ӧ0>"6yz�X�����s6J-<�=2sTv)�:�v�z�T��맳�6^SI,�p�F���e��Z�} ��k[پ�͸z۽��nmc���e�]�d�E*�<V�N]�N�j�ؽ��P�M���!#��E�mR����<d
e~��n����:;iJ�V�N���Lr���:2��T�lL��ʥ��IJ�ɒ��`��Q�yw���4��p����?��=��W���%��N�୷s��,wn�U���=E,���_�(�iY��V.���V�.�j�����'X��P�A�2�|�
�t����m;o6��*��\���Z%ǯ�x�Π�J����/�r�x�H�b�f�+ܼ<��F�f��DG���ֲȬܾL#�o�������k6"qu:G}�����эK6����    IDAT~Zݻ3E�HJ_Y��,�m����̦*�UE6�zȥsxl�:�l�|�BU�f��J��X���?R*(����"��*¢dބD-=g�E,�O�
��M=�eKg��pȖCġ�Y�:����ccD�M%�����`��^���[X,�vN(����
�d���>N������Dor*8�|?��bk�V�Z����=�
����p���ܸ����_sp�S�=h5�u岊�jܽ��X$Ɖ736��?�&<[����R7+jcY*�r�z����6Z��.��ɜE�,4�$b�������G�h�����.������[d�1�1[�FG��8�D�.B́��W`)�6�N�6���x�1�M���#_)oW}I�b���%e�(!�ק`Xb{^^�`�="�v������F :z����ΰza��]]LM�����ͫw���dfϐ�˻7{�J���7�PC�K7�����ɓ�F�_�5�L��M�_��r�A���b���Ot���hTkT�\��y�z�{w�+x�t��c�R)cu�h��\�}��U�������2.Ta#Veay�LAz��^ �u��m`�[�tPK�Mt���̠���&j��r���}p'z�_��@�I����o����ڌ��E^�-R,�����G�&N[�<O^n�a���bd���Q��h$S2�H(�}]�N+Ւ��D4�����&{G"9�rS��Yt���Ɇ�� �������e0��Z���>�^3��*��GK��-*�,����wz�	��B"W��JBY���2뙚S��+��*����Z�ݭ��u)6ٽ��u:0�JX'a��Z�{/T�nr�Z��9�V.���|�Ǐ�+�����Pn���z+�8@��� 4��v�̠���o�T���S��p����U����`|g7=�6�;줣)E����!�̰��S�r1�tm�WK�d�FF��?#�Ҫ.}�r�p$F&�!,�W���H�eKL��s�t?:��F��V4�����6�\��%M���U8[���6U�UH�2E��K#�3'�;��on2��d1�m՞���U�$Y;_�~[�k�l�ɗ��o~�&�X��~�BU3�2y�j�"۽V�V9F����o&d7a�K!w���F����?}��E���C�B;���)�����t��o*��f$���U�����5m�u(�4Ir3���q�̬/�&��H��3�ks�
�LchTq{K�,���7�L��bv��7+
9������1�<����p��A�L��h#V����o(aZ�י�Ќ����jJm,ҙ��(M�dqbuJ^���oa�L7c����X�LR���)/�ɥ�h3�lJa��w}�kP�I�27�x9�_����P�o��&��"�{��Ơא��ؿ�cyf�c���4������ɷ����B��JC
�Mʶ$��J.�¹_�7�G'B���1��Ov�g���\fJfN)A�TRI*v�ܶ��abv7��D웍�?�����t��q�.�X%�fJJf��|��y�����+JY7�9�w�~?_�r	�����]��/��?9C��B.�E���txx28ν�Ϩol⽳G��Fʢ�݇/�2�UPx�am��r%�N�b�RYRqbe���o��38�D3}��Tu��}/��V��
�:8�Y��d;;�$c)޾���Fg��=��UA�maf>õ;C�̬b�W������B����$#c�,�Deh�Җ`�Z=\�l�\.F�fv���gjl��u	����)�vS����C*W�0m3�U:�y\�m˳�t4����XY�s��K�������N*Ba޼%R�@Kw3��{����eBA/�~z��z��o��_M��G�$�yM%+.�L>�đ�f>9Ӎ%��(�(N/.����	~�������/??�-�.��Ǌ=������]�����>~�K�Kar.ʳ�y&Wb�%�����5�����N����Q�����+�S����[	��`Zq�ۈ���Tb�K����Z��\.��	�p�N��V�n������c�M���� �Љ��a�R��7�E�|�C)I�pj(�s)��Jx�@�>	[�̲�0m6v�_�~��&5i��%٠������)�+��㷇������������������~�#G�ŗ��pi�;w�kO?_|����q.^{�:L��߳�tkb5P�l��Gv��4�b��~�����KGg���e�
�Y]��å[�om��/���YKjkC��~.�������By�������P����7�5#.�8�Ľ+�����k7�3�4w�n�[�E����N6�����\\	���J�A�̀�(hv�4 "M�x��s�F݄o�7q��|K�h��Cd�zY�x%1���XÙOh�Z� g("���IV�,@d����������X$,^�[K�.G�Lt3����9��.�����������hŏ��1���;�Oq��n����x�>���g�q��7�SrTk�A�T�l�\&��R�e)P����]Dv�b�b��"�)q��]b[[��W��4����dsM��|�����'꿉nnRYS���������)��
��I���K�������i�ݼ���k��h۽��=}�|���*%���V��{�Pc�6ׁ�Jr�.�=�W��!�`��7@2�Q��lۅ��h�/�Yv��֒N�A|s�ӎ7��v�)�)�v]ֲ��h������Xo�S���T2���s��eI��l�[0M�Ld�]��D�BzG)Χ�"�uq���F�9y�0�;��36=�����O~����������;����K��-ũ�i ���k�fPJb
ir�U��foo��٬��*Ml� �����7<������gӔ̂��67�<|��EN;DkS%eK	�����5��2�a��^���JsM5f*���xt��(����G�h:p��νd�܁Mu5x�I�N�+}c����NC�mT�lZ^�6�.Qy�Ԑ��I'�lig&W�Y�RP�d�	Rb!�N�g#g�-&l7�	��� Gj���ZVR���LA2;-��A�"+3�i�u�޹}�
&�/��i����ǈF�\���X�������*���$�i����Z�ޛfrj�Lу�[�rd��E���([��@_'�bfMU[���3:���O8�w/{{Z(Hޝ�Xm�`y���������܌�.���*�������%'����	-���!�)����=��)��(�JX���]�Դ�`�W��!�K������M1euq�͍M��567�	y]*q���TB�^נ�IEH�ry��6I
�Xȣ�^���,�<Jt�M��7�ה�/��O�����u��d�94"�l��®*���(����t�p���,Ks+8{�;	���ϓ�%ijߡD��D�T�ʑ#�ع��U�tS�b�d%SPȻ)��l��!���UF�(�"o�X�ؤ�������ʖOr��"/^�&����ݥ�a��F3&of��L�ZJ�#�zY��f��ߦ�i����\��C��r>Od���RK��*CN�kL�eks�#G���B*]R���\�;�HdsdKYv��a��2��KQ��,oD�dd����b���Z���������Xfai�h,C� SN�J�c�]�D�)1"�fP��M��\���*��q�X��y������Zٳ��677ihl&�N������㚛���Gx:���{�)[�p���D򑧜Z��k�ۏNQ�w�VW����J<͏���D�o���l�2)�`�Cp�.]S�g���a �i �XKH�T@	b2ٗA����\Q�����3c,���yC9��Q�#�Ka�bk�^���]{q�kpd������S�+L�͑��qjjjin���m19�J��a�MZ�W�d�[l�G^V?�M�4�D�R�(TTx�o������ba��u��g�U�hrES_���R.�gRų��딲��{�Vs���>����O?8����w�r>qo(��7�e���/?�C�/�K*e��W�͙Ե4O��D���(��|z�
�IA�bN��E����ş��l|��T9dy!8{voPɰ��ߦ�����V��ic+�d`h��K��Jmsy)��KB�*(@�2"�<�Ѓ+�ޡ�1	���a�
S�{������������|�n�f��ΰ�g#��nI��ƺ*��u����L�}�c�9��%��E��H�����&�K��%�f�b�ɥ�����ˆ_����$iKB,�8+mZ�:��̜A��-�8#͵�-���0mM~n�~���9z��~r��w�2�+���oCkk����U^�fߞ>�����2���+X}A--��	����OSJ������O��]NSH��n�v|��WoP�P�g�����vؕ�hx켙��╫TUF��p�)�L9�����+��/��8���L�7TWI�"+��<�u��ї��`����A��S�~���q��0�Bc��]�5TDm��!HfŃa�J
�t���BDozy�l��"Yӭ���?�D�ir*�h�<�I�D��n�>�2Q�֓KnjQ���F�`�cG=}=�};���,���P(Ic�a`6+玁�%��%r��������;-�Nm�O��G��;���\�4���������?�Ῡ��W������ՇL/&)�Z4T[P�")�I����BX�|vn;�<���\ٻ_�UW~������9F��V�ɨ�4�^Z�r��#%޾�$�]���z��vw_����	pW(�\�+�K%�Zu����C����a�޽LoO�=;�t�&єA������q�B:\tX��U��h���ߎ�{Em�l�D�K˛Z�W��Ř�p����-��@���Or�!�R"�I�t�5Ƿ��൘�ӡC��/������~׮�Z��Z����@��\�fBoN��֬�⓵۱�2��UzZ*��{IE\��;j"U;v�[���Mq��q6�ֹz�;vt����~�D���{�j�I���S�Y���AVt�(!��o??�G⥒)U|��Y�U?\����2��/�=����d����槻���7�~@Su�\J<�NR����<_&VtP�����T$�aj�^������_�{z[�'Mݭ:|�'�Y�[���Uш�����.�j���}�"�r���#��m+�"2��T�YV��5m:�5-�%;6���
��".�@����-��
6�����$�^�J%�Z�TU� Gj�T:�!ԡP_�L^��G�ek!2��f�f2���ּ��z����/�ݻ�#�w�|P gOhli��;G��oq�_����N��9�V���헤�|�0Y��W�x�v#�������==�*ǔ�Y-O��fdx�޾�{۵����%����_155Ñ����Ur������1���"#�E�n�z����`ͦy|���@vqJ��'�X�p=M-ѽ��ݏ'��&��yr��ӌ�#����oGפ�@f�餝����\��c*��޺na�~-dN E�.�'��)��d*�?���Qs7W���A�nm���DM}����c�nh��e�+u�4�E!o�<J/����w���Ȯ�V�FWx�j�wO$	�Å
(��l�op��ڻ;9~�0�L���^��(cqUcZ<M ^hy�;H�ޜaOW��㢾7E�"j�ə%=|Lߎn��(�]9�}�^��P�;����$9 8]V�I��#sL�JT���l�L�OJbP�C���Ky|���7���
b��`�;�k3X��UWSQ����wd5x>����0�z}J��d����%vNH�ܾj���c�%�Rr*C�S�6���5�N�C}���/ɶ��z�?[(Hf�
�ҿ'rN�җ4�^6�gg-������&�ۤ�����Z6�<zFe0����ꕽ}�6�B����a�'/XY\�����{�Y^�����@�FZI�tyHg3 ��BRe����^r�/c��Λ��"��ޝ�6�P�&�~��`<�chhDL;:;��"�a8�̬�Y�H�͗�ֳ�)z�"��è��?�-�._�rٍ�]���e���VOk{D'����/-i!]_WMMu�$� ��(%_EyY��������ƕ�(�_Yuڌ�L=�;@<�-�q�?��Q��nOXQ�fɊ��A��fA	��A�l���o( ���!̇g�ȧ�����E�p����4�4p��5F��r��Q��ϫ�q<z�����eW#�����9�΀zE*��Xڳ+4z�����卵�S2K�.��^�N1���o>�+lF�:1���������v����u�d|y=��IF�H�<��JPd�T.pXL�*+�m,O��:;��`j����RB�=J�����@u�)"-�8õ���Z��6@*�D:����:�x��~[.�tG�&	��تp9k��,��ڒ�od��)�d�&͠<\b����A���[��t��(j���/Ⱋ��J(D�'��H�N����+f1���g����_�33��������ǿ�����xQc.N�9��c�\��/_q��q����<O��u��PMmC=ф����\"�(����P�40�q=��Ë1��x]��o���*{��&6'vo���S\��6m���{��J��ޣ�c�<x9M"/2��nX�eCW�2y���P��2��W�yu���8�cڔ�P�s�t��0����+����<e�W,oz��̂�+�hp�sVR�V���d`(O9��i�(�{6�1*�a!����V"[�Z�a��ɗ��%w����2��]�K���Gl:��*c�YXJ"�3�Xf��F����������#�mm|��y�/����J/���-�����3���A���3t��q�������(Y��V�nJ��PJ.�����N��6S�532�]���46���'��粸�-������\�rM�ŗ�}H�-a��ӵ36���!� ��5F�(:�����̦X��٭k�ƞS��`X��+0��'�r��GpU�+$�l�O��`_29�a�)�Д�D��g������r������J�%�8I��֢3��`��*=����3�M�A~��.\;S3<}>�����V�?�1��Ӝ*�l�m~
�I��A�[���"��*`��g�i�ws�Ơz%�y~aE��u���/�Ol��������?&�sbz��b�ɪ�Kv�C�G�K#��g��m�BjK��s3h���;�.�+�b�6���r$Ori=�O7���y��ivu5�KD��4�������1LGe��_�MMgkB�z��||���(�o_�������f�����i�߼O�J�[9ƻ�����*
y�	z�v�X��1���\�6��y���+���V!�IiN�_me9?�qNɸ4I�Sdc�k+���^�.�͔�{�.�o���ɱG	V:��p���\�jRy��
 Ȣ�Uؘ"�-4��L�_���>>����&/�� �*��#�)��8����Z�G&�s��C��
dJAr�ScH4@���g -��ɷ�<�[P��U�9��k���[���|EM؋�Mⴊ����F�+w����ן}���R:�2؜���B�{����Y(�W6�3��6RA�����k^޾�̳�����ʑ#�x�x���%���J3��k�h��_U�#G9�����N����x�ꯒw��%����:,�Sp��s�ΐ�IE�ɶ�� �d��U6�B�g5�4T�ػ7����gψE7���޳����r���%lN/EîP���@�,J��#R,�֦���9ud�-n\���{��c8<�z������yt�&��UΟ>O�����y5���'j"�*�G^�}\�]2�m�����};k��9��6!�[\<}9���8;w�C�'��R<��������Oq��>v�l"���Ĝ�y;��۩LW��|�eQ�u���P�-�b��e^����P�h3(���}'�ܱ��#��j}U g9I�����2�Z[_��S���զ��B&F*�������"��RD��l�-�!A��5L�%q�Kj	��I"� �Os�݃�����$�`bd�L&��}�Ֆ0<�����f��tS|��lxe�%��ժ��Q�FN��������*�l�Co'4�pGg���
z��#TTU���4Cog�Ѱe�    IDAT��"���S�N���_������;4��"�N���B}��	����߫�����.�Q�^�jfkWW;�{[)J��C 8��k��#]8��D.��13_&���2��ſ��򿒏��@��n��:�`W���wx�WVQS[!�<�4�~C��v��d򢀐Z�@��W�l0XC*U�8,��*$K�� 7@ȿ|q;O]��U=��21�!6��r���QN�=�Wd�%͓��X28�F^�b-���@̌�)�C��n�2����+�k��8z�L>��;dJE�8L�"���$7�9q��`����߽�0�=��y|>�F�31,����R�(����;ɶ����:{�졡>B>�T���*���ʷex-�u�
c��,��ٌ���/φȧV�x-xIa�~��i3(r1�+��]�͠�}~;��A2�It-A!��e#�4 "k0����:��Ti�+t��%G:�Љ�4^��,��<n��t2��L2��L1�*aдۈ����"�e�b��$j��a-h��r�6�R����ρ������|�o��5;z[����O��������LLo�?��?�?��/ɤ����7I&
X��`�pl{��y��%<&���5>fZ�PK�\� ��^�Iq��~�9>��e�LD�1vF����?����}�ɍ*��|�WcK<�b#e��
���5V.TUE�����8k�c��͠��Z����dx!�H]�)��;qG�Ԡ��Q]�P��r�l���|�͡�!Ѳ�����p�XZ)�H[t����>[���Y��G<R�[��Xʊ�/�28m^��$j�T�)���W��N��t\����L����M�4�?�����z��SW����<���w���p����69���4�U�/��k�����~�?�ǋw��rWP*�p����O$�s)������Ժ,�JX�3dx1�_.^�f�_}H�4���fP /�ft3(��s��F�Ԇ����:7����魦 �9٤ɤ����"BU8���C��2#��͉�7�6o5�G��8�+Ҍ/"_
�߂ו�b�ʣҳ� -PL���D^��-�mL�H�^v޲4�"�Dib�ЋwAO�$�E�,e���N}�G�>�g�t`S[S�������678�~��LҜ$�i\>�nG4h\$��"��ȍ�8���v���[���W�$\]�����@0���,S�k����9�� t���2�_y�R4�>)�j��q*uN�4C�:�u���D3��;�*�g/����65���g�ɧs����q22����W	��w>��&B�o2����
��:�*�A���j��J�4>ɋ�?{���f�Q�$=o����Q�}_]3��0�|T�:_�=B[%n>`q~o���DF7��EH%���d߁�\�3����p��q�.x]�6�qdqXd�(�[��4������t/�r�K��v��|[���*������1<y�t���ˆ@�xs����?�U���ٓ�DN���z���	
�"�t���V�?B[wHNو�>2��ٴ˔_�Jnx��Y�����gW��2��f���[����������i"�Jiq%��\��@��Ͽˮ�:r��v&��ϫ�e~#k	�@�"Y[Ţ�?;:;�:,�zr�����1�޾@{�@�:�"�`�J��s8���MԵta��a�>8D{����\KR�8����EƞH.ӷk'��tr��<c��N��KA�LfT!���i5R�l2�	O��F���j>�����%��먪���x�"�]|��_�f�����N�e#Q�ԛ"[����v�e�CIݟ$�8�ߞ�3�9����z���n&��Jd��Tp��*���<�����^E��W���ć#[Vٿ��YJ�u��2�����\"��z�M����z�����7��X�ǒ \A=�|���{�/�������Nn{[�ײ\}�U���W�FF<�;5B�x؜|�����{�Y:�[9r��<V�re���JJ�
*��	W��f�Q�`�'9w|?5.�tp& #���6�j%�Z����HU����x;���_��Q����B�c�x�w�x5,}.�k��6T��G���V&��x��k++�������ڍ*ۖ��L��%6�W򡆿Kq�Z�VJ������Zɤ�i��w���Қ顠����?r��-�M��=0��1�[N�A:y%�+�I>��������=-9�˹3�|��Qz{{��߅Y̪/MW��̓�ϵ<px?=;�)drJAv�=�,�[ V�͉��MYʹ���^����.H3�y+����q�)�v�#���V��v3MО�������x2���;H� .�"�r+9��8MQ���ޒH���IN���t�ӭ~�j��R2�Lg��I�?w������5U!�<x���dΟ?�Z����J�
�Eid�Z)��v�7�Ģ�
;~���`iv����bqRɸ6 �H��==T��2�����T	���N��H�.Ϥ<s�R�rr���0�v��>��1 ���<zB�6�}*���l��y��7#��������V��%;�h0��ŋ�Y�;Eid�%��Hz��m�Kp��ܿ���c��F��^��Z:��P�ң͠,�jj#�2hk𲯯��8A
&���߰8��$.�T��O��26��6"�Ĵ�9'B	�0��^Qՠt2q�W����b���Z���njw�v���>K����<Ks)�o[I�[��w��(��l����3�b��K�Zw���ph�T���6�B�����h��og˫)��x���� -�d�,��`{�Q�k3��\���VJ�����/�(�xϞ���ȤR
�t��
�y58��`Ϟn�>b��X����Y�H��Hi޻ܟRKI�r�,����fPBk��*��j��
���q|	]/�4�1���Ig�P'ݬ�#��X^���	�HԬN=�����'�Pw�E�w��	��N*�2�Q����*�dJ_1�VE"���)��2vkP���m�P�,�dbXLܶ��i�������D7����L�"���Ϲ�h���np��iμ����s��3=����ރ��{��"o�u�!!�y����->G����`�ǆ��)^7��4�� �-���_��4�2��rñ�9~�����h��O����Rq�_Hq����Y�����E-����fP|���ύ3?<��Ai~"Y�E�������w�4���h�-�}�v��G���x��lH���Q��������A�̫��������Ŵ�|Wd"��2�30U9R,&�LN��m�3><���<�h��]}�>%Ђu&g�X���8|�,�$:�3�	L�)D>M.�A��&N�Ӆ�]��������6Z[Zy�b�T"ϑ���%�ܸ}�gӿ����un�~B"c�� _�{Ǝ��Ռ%9
�-*\E���4�N�TT���� #�)mE*'�`��DQ2%m.�� �o�x�&u����>���+�j5��o����	�ih����]M�"K���L��5����w���_EM�A�;��l��"�Sqp�T��>�v��D�\~/db��(����Ĺ�h��-	��	O䡥����$.E��rb"��L���-�<�L4������ާ�����cm-Ͻ{���R��0M�n�D�d���u)RB&K+#C��'Ghy��O�cڜT�5���sm�wt4���C*>��cB>�ܜ���
e{��6+en��	^��%��&�;���d.3�]�(��y=�+�ih��/O���$WO�ϭm�t���������\"���h����7M��s��k���l"K8ॱ��R.���4�n�9��bl���iD�P�`��^����o�[�H�Bv���;FWC�?��?���8Ս�RN�����`m�-�9�{��ʭy�\�b�PT��y�)����7���F�n���r9u*�V�gv���+2�$�N����)]7o�9��^���~�ɼ2E.��-g���Sd�	��299�3q�Z�8�����������N��wJqR�����>���icc+�>���F��UH���T|r�->9�Ǿ��xC��� ���+��069���'��ߠ�J�߬n[��n�gey�Ͻˮ��	���!�淸.E_�I��Ӊ��"�������G�H�ΐ\c��E�w6����ŋ7Ie�w��l�[�Cus�naK�(�����Y�ӟ���R����3H�c��	�8�Ϝ���>�ݙg`d��ţ�LpD��B4t��w�B1�0�����;�[���<�3�۷�|�����	�餢���=c~-G��I�W�M�^$7N�����"��Y|�{��`_�wth�+�Wɸ��C�Ӣ������1N2o��U`�^��U������!�7�5�v��|y���I.��V���-v��z�Wo��կ��͟fri��D�z��E�����h�PL�U�`8},�K\�3�r�@N
4)n2�zy��j�^6&^�B6��f6��٦����259OU�ʡZLO�P}��jjp���
)N�M���ڵ+ĒIB�$'��+�����͎�v�=����v�PjR$��zY#td�-0�|A��h}]�������:X]ޤ�*L�L3��5c�|�,}��~s���$Vw�D:�͠8ݷk�����t�%[����VK_��)L��Ӽ|=�F"�f��MoW3;[kY^Hp���7\�����e#mQ���Q�
R���m�@��%kP�t%�ɳ��yî�^���"��`H���F�n<z������R�R����g5Z���iVby����)�RkC�v3(2ѫ"�B�9m-�:����z�~�Q������iB.S�>���C�>_D���Y���	��y�9�����$���$��Ŏ!�X��|>����-���D!��A�G��T�3��m��45Ա��������ei����a�V!R��F�ͩ�G��%��"Ϥ��01���8���5D���JW�+ʏ���@X��f�'s�=!�_��W���[�5�r#�B�4��mJl5��-6��<~�ֶV��J�%%���azZ6������i8��*�iW�%
V����n�X	y�xL�[�~��?j3(6 ��NFE���j�I���!iu]�����ٓ-8��K��W]������� ��45�y;�����
��|r�z8e����-�t8j�/�Z����\_C�.����ɷ��A[G#-mM�e��V��J`�Da�e�X��M�>�(�ķ�NE�ž�Z��N����"ϲ��h*�ӥ֤�Jv������s��{l�MQ�ںnSΠ�`__+]�!l�Eٽ��ūa��״���ހS(���R����܁�f'�����6�6��'Ҙ?�Kλ�JnX���e�'�!'P��*��J��p�hi����9�K����e���"�]�2��O_�+9�Tas�7"�LX�+-c5Š,~���D�'b��u�pho��;_�0�z����#ij�brf��g�X9<%Rjyx˔�b`_�e{�ݠ�����^Ο����q=�ñSXX�d��3�>�E�しTIA��	�E;?^PR��WM*k���,VҒ$:����"��;T{-�y�ù�������şT.��o�"��P�eu-ҽ�y������/�i�!S���J����C��ZW�U��,��i�2�i���$ksc,��LtmʹnGe_v�Ҹ�4�{43�������8TI<�L!���RV�b�6X]KSYWA���?��ޣ7`�k��i˫9\������=:ݒI�L^�BN-&�M���#�K�4efFLʏ��u��a�v�tp���9r%S�0B�xO���H |Q�<�l�����;8v����Q�Fg��L�����p���T�W��Ǚ��k���X��!�Ω���K�l��D���f�e����W8��r�?���n=��GT�K��������"�ޤ�������W����۴r��C�+�=UPv(UV6�B���U���Y��KI�#���$!XMe�>j:�����^�����_��J���u�nJƟ�c���P̦u�����r�ōGc�mq�C�������rMJ�gR���
�%ʞ]�>�B6��h�y�f����>��yv�4q��+ݪ�JV�&��V�A�T���B�=��la�%M}��o���V��b�����"+6pTY�ܹ�	V�y�|�{c$�n�V��t.��-Bȼ���5�Qv�U�����"�йF�V���e*�"����T�%s��������e��������Odp��*���r�C���`��k������|��`&���o�cs�%��)��%0���ZqVv@��`S�6��p�\a�Bz�O����z�������c/��:���;��M\���דq��q�"Z�@FCc-6�	��f)�[�bk�kt6��?}����Yn^�ACm5��Ż�*=i��\�ۏ^���t�H������+Od�\\�niC(A��T���IJ��{vj3U[���J@�#�2sKe<ֈ����C
���L�!e����Q�A��1�1>8�Ñ��Dr��09�Ƶ������ؽ�N�e����QY���w���烳g��[O>�R�?�73\�?�Z���6}��������E�����D��4Zb��:w6ӷ���^�A&cе��P3��]x"5�55���省��O73�f
a��M�\j�ba��>��cG:���/&S����{(�E�Jp��esN9�0���>+��-�����nV3����;�� �Ο���J)~����4�r��S�<21(�۹�Ҹ��)l�$.k��$���V,A$bGG';Zە���a`}����1���E.���R���o��om{^���AT.���V�ן��&�T����S��l'�z�gCo����hk�`�0�#��i�����123˗��ήJ̔�
N?Y��ϑ��H��Y��,T�g0�eut��7/0���&]=m9z�w2=1K��c����m&R]�y\2H2r1��ME���?����5�j�5L7;��@��~�=��R�dwer�9ߎ�C3��$]C�
d��w;�m�rho{��\�p��͑#{�yFǖ�kl vq��3K[
����%�?��bų�[�jCv�|:�E��^�6��a���I�����K��6�v�s[��3���lH�����DB~�l�d+-n�\j�}=M��H������8�V����d����ThY���<x����1�Goo;�\�RF�e~6�e�9Kh�l�����_r�C3�-�.�m{ͼ�#F���}�3(�` �?LME{9�ۚUg$�abj���ir�(KĊ���iml����,oX�v�f�IԆxB3y?�(Z��]��E
ٔ6 N�����<ާ�74c������z�.�o6:�����E��z��HE���FD��f6NEȫ��Tb��%Z�*��i���9�Yb�$�s"?�`mS��^�#�d����ސa���� �bɮ��R��=m����J|�-��H���fإ�]Q�n/���WoF�������]}�ۖ��U��6��rivM,N���� ������sG���2iEI��a�����0����.|�ajj�f��ZgO����ٓ'x�n�n?�tN�P6�^��=��������v�9ԶR�{W0�v����Фh�(�Ҙ�(�����)�H�=�Q�|�Fs��=w�L���̒*NdX)ʵ�l�>]���P�W�Lz��������JU|��)�f֙�_�X*
#z�[U86���܊Ү�Z*ûR٪�r*�0F��r>����Z���i΀*���Qk��={hj�Iep8$�����W��p�<��׃�%�4�E����œ�$�\�l�m]��\�2"����A�����o7 �����<+��A������6׷��j����P��Kמ�zt��
���K>��$/S���lX,2�"��,��E�Ϝ��ocf2���(�#�q�m���iy��f�bɩ<2��L\����+��Sr�ٜ%�(���������c��,��+tD�P�hm�d�]x�A~�3���i�I��_�2�ݔmY����2�gV����P���4LO��d�?�pI3g���B^�b��~�;��[�/.Q����    IDATW]�/?}�æ���&Jn=Q��S�a�2���ˡ͠�Rfua��Yȼ��ķ�A	���eI�3�U4�>K}����v-����Ǐ0�vL�얐���W�+f��i�܇�x�j�{�0,A��H��/�C�S�"�4���A��0KIn��?<�z�\2���o��p��-�� ��~Ã�Q�L��;0lm|�!�i�Y��?A��G���\����=�;��_f��Q�h-og"�<T�V�ֹ�d*�݇#LέcsE��WO@�p����X^�&�疒T8�|��Yj��\�|��fpl9˟.\��%��JO�R.�����[�╛�����3��BK��\$���O���EÇ!:~��H�^.Q]%�Ai綛�W�(m�@.�-�	VSѺWii��.� �4�������MO����tfL1�;��dQ}�?y������d3X��	㖇�,�R�l"ؖ\�oA�|,"!-g�$�9w�0�z*�y�.U5�������o�����9��_������@=e� х�)�^&g6����
�I����U��n��R���]�B!=l���6n�������_�r��Y	Z��������s��H:bQ6��fz�������g-R��&^P�����ˏ�x]��o>�&����~f�|�6���W)����2���p��k�+V_X��l,Me$�Y��t���I�>����+���!�iہ�n'yW����q����ܜ�H3��t���۷�3>�P:�lq�>']�!��n&�0���]RE?N_5�t�x<����I���S1��8�E���i�z�����`~f��8z� ��$s9�<ey+E�����孬�|��M��"�i*���e�W73�O�$������hOdRD6S9�!��)�d��]}��d�����R0��s3��ѝ�]A!���f�5\������������]O*�����i���kw������S���D)�!�N��T��.�כϙ]Kc�"
u��q���\�n-MR��3t�G��k��h��ş��mt|g�wm��F��ȵܿ��'*I&&����R�����w�)��O�2�e(N]�Q�k*YuX��^�?e�`B�ܤ2�aZY����Fvv53>1����=�5�R4JL/o�xh�]�g޶�^��-�,��]��\z[yS�b�#���rh\7_>o@�;�\a;72�"�JS,�ֈ�O^|�?+ �S-����24@�Bj'9���q�*�*�o�O�A������W_I[S6i�3)<?y�ƥ[�x=:Χ���oG5f&�A�WP%���av3MF��?{�%I�Ӻ�O���?����;���t�tr���߽���,5{�b�+)8B���o���I����*��ag{��W��/,(�%��+TJ",�|�8v����/���a�"�0Kd2)%IZ<cڶ�$�q
����b�	Ӡ��;�x��	sӴ�4��.�/[�3�J/ۼ�
V�W��"ߕc�*�&�J�(g7U~*`���M�ҹ�v��h�h#�ƷH��d��6��$`ދ�[�2[�+$�.�T�4A2h�I�Bl����8ئY�fa����T7��9}��>�C�m䙵�
y��%#�#8����N��LJ��K<�_M0��!ow�C<S9=����2?�D �0�1JY�a����9IM�^
�F����f�pi��Bt�ưd���eccK���f'�P_�HCS��4_��|^bzrB�.	WVkTV&'5�S?�4�"u�����hm������Y�V�����u`��X\�bzaC7��KY�Qv��F��DRi��`����k��4��Zb+�E"�f3T�+�`$H�Tdc#���N%�J��\+�uE�) 9y
�'���sr�Vrj_�H.#��vW@���������1�<yQ0y|�
x�z���i���oG����h"/G�Y���z�'��+K�I�mefUV��U���O8�-gvvg�P��e��î"�?C���J����$�6 �}��.�K���g�FL��tg������s��� VC�0"pMV�"�*��O�⛘*Y��V,.�]�ϩ,�xB~�$r��+���Z�_�q��u*���d+.�j.N{K��N0�Zfln��Я�%V����^��Gm"|���iY�:h����[Э}Ow�\����z�O��]Xc?�W�,�m!�O��<'�,��N,��l�����d�P7]m^*ee�����M�)f�2��f)��M'�6qiՔ ��!�}ːM8$�G[���)CC�-N[@-��L��������(fX�2n�L������&�pˢ�X�>�x��Ub��<$6Q���z����\1���F�O�y����7���3Bwo���)榖��xnjՊ���w����s�/.=cznL����Jz��+D����C������+���^�ǧq����z_�������q���~�L{K5A��R�29"3 �i.�JK%��P�׏������{����e�
����Ԝ��G3<�VK�L̄�g4��!���t1�pK9Aԉn�N���ߤ�U�`����E��կ~E���/A~|2Q��Q�������ɦ��ЮӍۏ��pZŠ�1�⿯��YJ���A��O��_zN=��I� b�hP��h=�2���X<a���Iw��χ���|�՚�`����T�r�D��y�Ǐ���`�5L�j��
�{]at`������?�����o~~���<ypW��]�.�h=B��0?�[���*���K�T����jb�0װ
ᩔ�d�P���t
��NO���[��(���R ���.OFfX�L)Q�n��Lj�����Zhn�b��.��dF�i�U��3�Y��//�V���C��L]�N�6/Ss�|}�^��w�y��L��j������[ U8�CZd`Q-��6j ���b�[�nS�_<���T��D��n��ݚ�MOKk������|�ɧb2V���h���-�|n^y����ci;����)�U�P�jJ��br��:#���V6�K�R�q��χ����V�7y�7�mb{#�}N�L��7g�[KS�1;�j3��%�+�5U��P!�G�A
���ۘ��1̑#C��\z��9����~���M̱'�c��{{Յ f���_֌d%�E����<��V��v�Y\ll'�ӧ_�(��o>R��tD	�F���v�Ͽ�Js��&�M�|�����l1å[�le��d[f��Me}�,eSl�f��m��c�f�D���"kn������J�Q�mry��!�	S+Y�ǋd�2�T��h��\���[�ܸ7���B]�Y|+�Cm���N���f��W�i��R̥�o�qz�_���n�����X\�����~��T�� �&�"�l^���f*��_&��'91�fg;����<g;!P"�A�L�rl�A.S2	.g�z�H1/����p"Ho�ѡ C�������}�t<L1��\,`�y��]\��ǣc�����1��N�*n��R��7Wn2==ǫ/�ȩ��KER��P#銉?_��ϫ�)��.���&}������ȃ[$6�!����/t�"b���R(��:���l�v"m]ح��n'?��ᡠn槷�3����5W$¥��o����(���
YJ���h�.��NJ\MM><^�;�
l�,�/1����u���18ԇ/�eys�D�� Q0�p�M�@�}(�lr-�h!�E{��O_?��.+�L�����g�NfHH�dx�R��@���b!U��P� 6[������j~0�.T�Z���u������T�)-���˗��121�G���Ζ�2,-�q��1q���<��?}���r�B6�b0[3�Ս	���d�g���X���k������o?g��5��]z�r��ynݺ���
��c�,[<���c�4��R.$��783����]����K39;O*���v�r8��򰰜�a��[�Rn��H2��8@� �{���(�RIi���b*� �����R�;;�t� n���=��y<Md��[��&��[�2(�F���)`��P+Ţ�ёq2��n�����X<nrr��d!��Q�K�ǋ��� u�6w���a�i~�l,���r�'��g�1KMHE��2��31��`��<携�	%dX����cLNNr��1��HI� �c����OfY�NSx��E*+ 4�l�a*��&z�����f1TR
��͠����/�9B��kjTw�X�*��QZ[}��E,��z���YDg��n��K�����4K&z���,�n���I8��9�ΣݭM�&��u:�b�$�N����9�Xk3�x�x���^��t�L�D�d�`s�FN]OB�-���5���'i
[���15����{�$�B�;�A����.R(�	x}
'���QpQ1��x�ڥ�,6�
���-A^<с]2����V���w�����v�G��ǧ�YX����#��*��ɪby|f���$%���e{j��������_}ƍ/~���0Y-T$l�k���D�Khl��|��^>׍�fb�ٔ�{�2�W}T�c3���Mkg+c�[�mŕ2.�9�,)�H���eY(^���Z���)��hj��������P�h,��#��<k�Y�7���!θ�E����P�_v�lv���,L&�)�j�n��4F��.э�]F'7Y����l�+U��'�ƃlKz��J�l��;���j)����ʤ�O�XXZcxx���E��w.�%�2cOg�^��ۇ��<�%�I�����}Vwz��A����X�&���������vޠ�\�Fܮ �r�����<���)�2��zT�H�O��Gy��^���(��%�Yt@H���lF���DT5,���.��x��.D���p�B������67����U�V;_\e+e�P�`�e
^SpJE��Vy��p�*��>U�PΦ����ؑv</�m�?����c��y6%�c�;1Yܔ��3#��ř\�p�~;�~�!��ڄvf�h4k�?��R�4���#����\�����.��+�;���=B~��0%�V�9���ʭ�Zr/>.���NǍ��^�-��4���(y)�1X�ct�蒯�5�~�U�zO`�7bq�T$G�=��u�ɩu~�~���6{�U��YV��������<�X�f�P��)�DK�+�uJ2��ɔ�F�/���OB��=Hf�̕���n���O^V�+���b������� U�����j��S�˺��/�4������J*�ew�m�o������H���LL-��%VK'nwX-�2��qU�G��v��{%�E�Q�Wo_ "����y�X�>�v�|v��'?|�M�>�S7ڰ�}L�������F��w_�ڕ�b��N�Lms��$ɼIIe��JN�P#*%�^/���7���w�`�/b��@�Q�z�h�����L%E����al37�}���%��U����Cgs�Β,�Ɛ(�ץBW�6j��ݥ))&�M&�6s�j!E�c�͗�y>��w�o�����A1W�ggn=���H�����Qx��-C�B:���!��i��Λ'H�n1�|�r�J*���v����;&�+��'_3����B%�/�,9ɧ
�9W���A��v��w�i��ׇ���:�ԗ�|�;{>��K=t��y�T�y��[\VvD~�g�G�IK4�4R�\8|v��K|ss��x��$�4��ǚtS�9;����$��ߛ��]�^���7���0ic��E�-8�Au	(�ޝ'�q��a�����Bl��6��W%���+�N̐)��I�2:�y��c��Y��1)��%��S��n���!��{���T2�������o~���gau���1<K��ջ`Q5{�K��J�P�i��W�&�hnp���E�PPʚ�<x����Yv�B��bu1���gRj����n�����\P�J�&=M5�J݌I�U�2�|�WO���0�T�� �mN
��zw�����<}��lFlCe<������-&'gx��8y�K�S��pD���|��K�X\MX�<�@��������;�M�����}�]|��U�9�9�*&_�p��.��	,����T��pmͲi���9ilv���ۃ��m����̔0�,d*B��k���(Sϒܽ�@�2�;�����r��M�����l㵗t�����{V���ͯ~Egw���O:���F�O/ߢ�KsC&����jT�\�Ŷ��P�D_^S�X��P���N�g��<x:��n�P���TFX,��[�l�,��tP�1�Lڕg@��r�͠L�%֕�TN󳟜�+j�R�hg��f����?b��4��#ڢA,��)��}jM1�`l����*ǆ�0U�\�&>�u#_^{��N��l#�.�Y��S�`��!�2Ã�_0��{�������}�.s�D����E*w<�Vܡ�X��s�m��2g�0<І�a`y5���HԌGh�%��y�h�͝4n_�\����H�����3��z���j�A`a�{;;z��m���!��n�ܺ��b�ܙc��e�t�d���2Jb㔔�Qz�,���&:�H.�Ig�Û���0;�`wk��ϧ���UǌA�~�{d�Q��~�%v�줃�,v7��7��!�	�l���d((�{�+̫���Q����<=�ν{���j煳�j_���<ov��;wǵ������R�e)'7e��[����O��Qpa*�ׁegK�b�2w�|FnmC5���H��7B��9���FZ�c�����XJ��[��Lx�FB>����I�lnY�ʰ�.�����m��@;�iV6I礟�L�%J�����u�g終�s�|ܾy���e��7������ٺ�6�2U��x��C�n�k@8Ҵ͜�&쵉WM�2��Y��wX�I�_�������taQU�����ժ���]��)n鏵Jt ����>�mS�Ě��lW1���;w���ͷT
9~�cO���[����cG�U��d;-�쪁gs[�-'(ː��b�ɦ[z��| ?�GJ����A*�R���J�X<xh�� c�g85�Ig�,Rrlo�O�i��\*�m�5�\�s��$�r�ڜ�w*��@l�.wT|T\Bۖ���T�45�4w���B���)ڈ��c{w���$2{�3���`�sЦ�O�r?����V#�!�hgw7��Q9/e�(e�ۭݠ�y�Lf5�+8"q���G���8�+�5���W����1��n�R+�1�:2�L���lo̄~���hd|Z������R�y@�w�l����)Ԥ�ީTk9S<6��1�>��깚_C��-���S188�ə�-lo�������0��@(�SSS�c'���u�O������&��J�B1�/~�cI���Y����.+���]1�k���	��h��8q�E��7>����.FO�\EԿ� |!�^��+�A"����F�+��56VW)�
�cnj�����j?X�&�������Iz�ju3&����V�!�	�������/�8w���a����8����W$I~��DC!����Z��O��/�Ҭ�o>�R]/�dR/�����4��0B�d<��H�����fZZ�u2������$��cJْ�ysiO3�"�*&{#�G^%�6�=Є��T�~�<?��Y�v6���afvM_-R��;�HOo�d��_�%7�f�X�S(epH�Tz3ݎ���v�N�S.�q�,:�i�3����O�r��a��	�wc7����vT�m~�܋���S�[��m��.P�*o�y������3�m�~"�@�K�"��[�z���P]C�;�?0:��!(M�t��j�v׈yM|��"���%�o�z�L�������	�Z�[�[��iva��?�����	a��t:��n��r�l1�՛#�*�k&/ۺҠ�hmm�<�����]c}������~�����X'&�[;z�=�Q���k��lt���N�l���.��~"���r|��M��
�*��kDx�!�i���9�>%͉��d<X�x�P�mQ�ON�M�ȡ~,&����ծǥ3H2oS1({��H�Er�B��]��@��y/T�,.�03����,f2Yl�'��fv�)W�:�:�����⫗)hY��bK��Fx�A��47����c�x��    IDAT��i�����n�˗�)��g?{�H�MIz?�V�F+�;)��t�B��o~�3�!Ղ�U&�++�E.�e5Q�f�*H��N����6x���O�)� �;C!������A�}�I�#�C�8�b�"*�b�(RͦpRǉS�H�݀�dkw���N�R _+���5Nbk�'�x�l���|��'�>��A���3����U�����[���۟29�Ɨ�� 7@ȿ������@������+�?����	4�R5y�O
qҫ�鍳���+v4�/u��z�\2NKw+.��V<�L(l���N_H/�e�f� �v�/�R��M-h����!����In{EkB>�I�\Zm�6��TѨ��k7p��Y�u��AȲN��W���<㕗_��P&���{X>s�����$O�dZ.��W��m�9`i�KS#����	��QZ[�ܻ7�����8�z���Swx	����|ϲ�����R���Xhjkcc/��z�lɫV"�M��YV7giim�����sY~�����q��i�~Y{����+ַ�����'���;$��|�O&���w�4_������-y��������ճYJ����,�-�Q��p�/��^�fkf���5Z[ct��c�X�.����f� ���av����d�'qi�P7*Fj�r^�~1X�R�\+��_���6^># ���>�Z�,\0��G�����9�Bv[\u�B�.��ۏy�l��_=��Sݔ�b#�����¥�3,l')���`�P�R*Vh�Ho����	|�9�cw�dvh�q��q�OL1;�H��(��^
U��.��c�(���j�bx�u��:��ēy�bQ�v��,k+[�2e���.����wt{4��#aJy�S�$�.!��tuh��ȓq��V>|��绘�Z���=�� ������=�Y�p����0��T��w��{Or�r�U[�d�z[8q����ٱ`����.K�kl��L��]8|^�ϛn
q	Q��o2QU��|�B/S������Xt�+�;CMH�u�]K��Ν�4���v���\2��c�����:�=��=ƙӇU��6y_?z��Ӆ-�Q��S�;Z-�܄�(���ܻ�9Y��e3(��Ί�>|�h�1u�H7v�)��"�h��˝�F.�O���e�㵘p�<d�Fr���+�XN�<2X*I�x�0-a������3g���˳����#X�&�^�����՗Oi�s��}�/^����k��r��9uc}{k��T��MM�-�+놪RLc�g��h�@�@�P���Y7��b�ɥ����U2y���%�V�t��DT��Z�⧨bR/�&q�)
U����cu(d�bj�z�ڍ�Ƽ�����@^`�24g�����O�����B�\����]&��(J��H�B��F�T�T�ܼ�%7����euɗ[5�0DZ�~�H� e�o8L$�^�g:NG���fm��fc�5٦��H�t�X]I3>�J�fT���H�Mtu�I&���I����HH �5V���"���-���deeQ��=�8�[,��X��R���M*&,�����MM�
�R���ѡnZ��B+��7�I���{Za��1[]d�U<Q*6�bM;7�GV|�5��2K���U��(�)���0�Ҭ��D�&���9��:Dg{�b.��7�R�ޓ�)R�҉}������Ww2̮l���Et��u\�^KQ���^��,x����A��zM�ÉS����RH]�R�h���b%��r�����O�K�;|��d�J��i�L���ĸ��f}s�G6LyL�,�z�h
���.����n\Kk�L-n�����R��eQ�@�/�C-�/R�'��K�9s,�S�'�&�x>�E�6)}�p�é�t:�L6��d"$�[�oE�dp)�**�ҥ�\�����oSږ\J*V��d>���?��f�9Q��ѳ�����o.kͯ?|����\:��O.����)a�X��'�����������\�dcz����5%d)9�h�dtQw�h~otW0F �t �$h����k�����-�X��*�-���Mp��,㏗q���T�UgW�1+�R�c���n�(�Z�3���2�#�Op�5�653��cǉ6zyj
�tf��Ӛ�,խZx-�\Yl�����ew���꣋4m�5v6�xt����d�.�������e�5�J)X��r��F9���`��5�V���Ƿh�U���G��q��m.��E��z �}�U�Ay�~1�U�/���˫��n>x�6��S(�T.'Ki��aoї���ʲ��@kk�Z�W禘��kS����`�Mb���hF�X�$[��0|����A<v���%*��
&�"OY^�a���B��GN,ΆG�klf��+�k�=B{G�c�YZ�Wđ�n^:7D&��o���)ě����l�]X�~�;��N�R�O�"��� 6�Q��Iŷ8���2�v�q�Ld�U��A65���>ժE��|թ�M��C��� P��ԚS����A�<���x����:cN��I~I���d�˗�)��w��,M��ԩ�.w�.]��B.ϯ>|_Št��@�'�g�|{��x��U��ɩ�ԯ�������'̏<$�6Ezk�Rv�Z)IC{�����#d�)`:�~��U��{�-f".7��: �3�
k���:�6����-N�w����=�ɓ������a���^�_�����)�\������ln�P�g�Zܼ��+�o�?��C�����t�lՅ�!�(a��4�k�	�4C!�J_[�����r�߾�4̞�~:��j�Y�D'����C������zYELN0Z��JZ� ���P�%�/��%���6mA+�5Lk����N��D���S<|4���/���N6�����/ݍ�:�߸ϓ�q^�p��(	�ZȪn�f#�q1��b��.T���X��9�����(�S�r�<��'::io�r����*�/�����g�O�}��Uҭ�"J�,��: P�$�%� �:b/�B�R9�`����frl���o�9����e6��9z�cS{|��x�^Ν?D_g3Aq��K:�}�x�O����o��&7���_�P�nW�
6`;�T���~�N�$����Ma��������:[imo���G�Z�K���k�d%��R�l�I.""x���x!�V�\[�v+.3Z� y�W����.�x9�]N������q�勼p���N�����T5r��c�=�W�r�L�tV�N��
���9f7�*e�T,��kl$"4��ܻ����u3���䩓�N�19�@�g�`K�9�5�1tB� �\��jf_k&��jDDV�UCM�d�`��n�l�֔�m	��������{�:w���'��bnctt���30����ln���=�;[x��Iu\�9���%n?����6O�˯ ��vG�g��d7�9����TY���~��:�b���,#�K̭m����;p��j?���!�a��5g�/I!��R�``����ۜ�g���.�0�I����F�6�{�.���gO+X��-�����(���44��p�����~0�0ڝ<y�����Ȋu�vaJ�j{s��TK\ᾊ�Y�E����w�����R�xqz4Ed�a�R �I�Tb����؍5�{��n�Ie�D���{d�(��m�8�#��ݞ�J���6���lnl���A�f�k�f��uw��׬T�L:I{k3���\�|�W~�B�n�_dy+���Q
�Լ��9;��1Ws�i�Hw��^���e���D�HOi���f���5
Ea�Ju�XOmzoT,���Dh�k�F�buqeȖ0���0rb��Ψ�,pJ%�f{�,?�p�p���/��1�%�.Y~�X^�����tv�p�̑����0%��	��l!��b0�f�a��i+r�K�����+g�O6��{�EZx荄�4���X�\�*���X�PȎ�Z�..<����<�"�݌L+�c�����������E
B��d�5�7����gc5AWGC~�W�<~t����Ϫ�S,�ހ�G#Kl�guh$ݍ�̊U�Gp��48-�;މ�l��csIerlm��F2��Aw�֫I�pF�l���� �X�i�k�T�حv*�"�B��&��	z�d3��b1���]erj�޾>�����ܬw�'c�ln��"F`De���L:TJ檌O-���bqՅ"���AWM���Q�U-x\�0f�d�b�T�u��A `eh��I�'U<�pɴ
66K<y"ЗE.�A���CĚ��y66��Zg��a�{����3����m��)���v\&�����h�s�ΐL�I�ʔL&n<�g;!�
��!��^7��ϝj�@���Z����aΝ��0[R������9ֶH�����{��/VV�YJw��J��h�`���5��
5�ڐ��b�_�q^ˑ%�"��f���D�/��B"��W|��A�MȦA��{q>��5����w�6�(�\��V+SKi.]B"_?�J:�<������R+!b���J{?�A��|�t}wc?v3�p�R9O���Zݧ�������N:[��r�p9)�,/�1=����눐Ip9,������߸���:-m=���!�ʅ�݌��r��]:[Z���3�o�����I��|���4�l�y0��׏3�\櫫70X�kv�5�O˄K.0l�<�w����˧0	��n$��L�y:��ӉE�w��,BX��HK�����<{�ٕ��T�'�NjV�^J����������v���Sz J�z;^��.Q(x�7hi���&�פ�����_~y��ˇ?}�h� �sj����*��zB�$}~bPhe��W��au~��;߲>���TK䅘VS�]���>�����JZ�f��b� �C�R٬ܽ�$+���$�.%�ք$;���#�$ַ�y�1�PH�@�{{�={
_�åo��M&x��yΝhfb|���������o���8��q�x�%���3���))M�|2Ա�Q��Uʅ'��h"���6�nЉ���.ӓs�ή��.�PѶA����
���Y�JM�Q&�Pjy���eTKCi��^8��cMZ�]�qX^��O�!�H�>RHM� ��V�� �l�KW����/��X�忈A�<�o��/P5INê/C)/�hm�������ȮN����jaU�!K���$�����Z:�E��ե)q����2<��;�u0�p��w)���o�P؍�[0J�������������R1�x<:��㡯/��\���l'�������7_9GwwPz݉��p���r;v���
K�i2U;�Xj����Z�i�SNo��������~���.=�]9t���^�E���	��0��%�jV��e�]�u�&p�-�砅ܵ�
�z!��\<��k���R%)����)n�x�/�Dog;��>����E�P��퇌>}��#Gy���T
R��ɿ�j�{ӌ�l��E�n�i�L��QB~7�c�X����`D�`w���.��co;C��,��sTܭDz���̤��T%
�M&|.o�����M+�L�Qʅ*�B�<�F��6K�����`��N5cd|tL��H�Us8���'S�S'�Po3��hx)d�<�����{>u��DI��5���uU@�&�d�u��/�Ӄ�f��W7x42BP2;�ǎ���IE�n����:ϧ��L�V��P1�I�� 9_�fs��@�z��@)����b�?Ƌ�:d��@Ω�?<�΃'�x�E^��K~Oz�k�l��]�5��'����I^<�O9�U�Y6:�������)J��E��R��p������p�ҟY|t�ja���vN�<�����:�o�![u`�5�>p��G�(��e
2d��qjD�>��M<��$��h��X��M�$hȶ"�����ʅ^���d������Zߦ�ك�o���gL�/�84�Kg�W'�~��J|��f?���N��dr���M�d��|N��	�U@="Oq����b���i��!b-M�����F"���s�$R�FNw��N�V; V�uO>�JM;*k�ݚ����&�Z��'��Pҕ����,�����ct�;q�P��Un"e࿱����x�NΟ;��B��+�����������U��3֬b�ѵ+?n��KX����r�,�G5o(�hc��E�5�b��Kw�ՠ�������$�q59��ݚ�X�\ޤ3��\��5@o��ѮC���]r�f�f�V�%�$3Bb7�����QE��aeyu����ۻ5R ]�;ɒ�fh��[b���`c�đ�V�y�$�LOβ����k'��ք'�%[�����։�+��T�S��(H}Y��ݒO�iգD%�TK9,��� Cݍ4���PV`I"Q�ڵ�\�pZFr�,����k;j�no�q�������Ģ�����'K8�v��0����2�En�c�Z)���U��#�>@���	iP-�p[���5�
�d��8(�
�9�7�����X�6��ku��"��FNm$��q��#��[ik����p��C�,��0�`�X���Gbz�ON������nFƞk-JO�&7X\��e�tęJ�L��)fh89w���O�&k���W��\�l�z���8���H�zW���L'd�%�UY8�RIl)s���l�F��SG;i
�I�ob38�ٜ�����4}��tw6�Kg�Dd�n03:>���.CCC����K��j�L2W���[��B>E��@�`�Y1��깚_H~T,�F��&Lu���RB�eZZ��/��"^�U��ҩ";���"l�d�H�ǋz�`4�����67�D�c������'�	^}�g��xt�>׮|C_|�!����&z�����)�M�`s��+,ɍ�R�e�B�f���}M�6Jp��7���q��grn���d��U�h�V֤������f�2���d�D����~a��Rj��^=Å#>*�Yg����er|��%�{�������j�ho�E���W��)�l��>�l�b�2-6�#ĳ��tR׋�A@_���z������6=��6QSi3v�b�A��F��7�VJ��ߠE��	�S*��fC�c�ʊ�&D�t�p0F�d��/����k�t���ͧ���#ǆy��<|����.o��;[5��������^�i�s��m�	˔wmy�Ͽ������-�q��[��W=���q��!���K=����=�yq���=r��n�a��6�y:���¦�ˏ���b�:5k& �I��I���Dݠ��SH������9�T�Pʗ�x�Ⱥ��D*�{?{���0���CE���.�~zY{�>��[Z�P���+X��/�uʝ)
�ٮ���l#�5�::i�zX�γ�W٘�OM�%�?����=���O_&Z/VW��bv�zvK˲�.�}�+	�jUj���P�)ͷ�O��/qz�ç��;{��cu9������~���w��*�����~�f+cOǉF#�5�ɗ߰���7�1W~X��k�C=
����L��M�M}V.y�|����?ey}�@���N���ܘ�Z���͒�r��h��dr�EV-if���]���*�>��+ഀ�\"_���v^~�[���l�͡/�?��S67v�����D".2�-�3[�x��W__%���G�Mk4��,�<!H;�H��`I��M^�r!��TJW��Tg~l��g�dV���4B���T]����Y҆3���!�bX�b?L����EN�_|�����r��#l��6?��A����8*LuJ�K�-e���p��a6�q���������������Nb��
�N��Ԡ���H>3�/�����Gϔ�i��/��yy�m.)� r��{G	7X�����\]WZ�lغ;=~�ƨ�����~��M��-l�(�@��0���$���"[R��%N0��\��F�~H�5�|Bml����>筷����~��:&�'��Un�}���Ǐ����u�2}w���\�3Ãg�!����a�E����vzM�>ds�9��
c��@�=Lww;#c3���	w'�qg�0M=�Ly��=�&T0b6rt���^r���Va��!���L�d؅�k�ᰛ��-R��9>����\&�;;d�Y���^azq���#
�(T�8j��m̈́�6R��E%3UVv�|&)�V    IDAT��-J81:�����O�*6kɚ��L5�C{��/�=�֦?��#Ϟ��O����li�衣Ě-dRU֖�Lά3��C\.�^�C��b�������b�ON�C�Z^��.gOrx0��$[�:�n>���^x���8@I-�v�$�;��7<�¹c\�0@5+��:e�������ˌͮS�� �*20��H=���������岣���Ǐ2;;���*��^�?��VZz���|T͂Ȗ���z	��JOk3����p��ro0L�(���E��E{۲�]<���a�z�	aqi_i��W����-��񃍝B�O����P��b*��ܲ�ܚZ����Ԫ���MR��$W'��\����K��?�Ǉ��L%�u�
��Zca�/���\����.+�;l�Jq�lĤ�Xj+L�K�ۡ������#J���r�Z6AG�ϙ�,1O��%Od5s&���gO�5Jq{���-��2w���n5s��q�V#��t���͓�k��n�<�Z0Tk*E<��f稗?�DE6�|���cj�sx�����M��w,p'��t�4M~�o=���P2�($R"�׃|���rb�F��F����m����M$�ՖLg��Y��jОZ�´�Dhm���q��'�*Vr%�
�������թ�^�I��pO�4�B�=���3ǃ�i�x����:�z�j9C�5Jg'.�K��q�RG�,5Lc���%/��||�  q$�%�Rvt61��.���x��7n(������t9�zj�����6`��9qDŢؔĠ�We3��膃�`	�ٮ[zS�ĝo/�×��1X����j�����-6LG$�_��4U�|.�<,�0F�1�Kک*y����Ž'CE�OVr4��FT'����h�X�������fw�O29���桿������.D#>S�gO7��{l�)�mjfKw�T��lX���q�x;�,-͑��ink����l��⬬�H�(U-��R����[��r��|��b _�>R��#Z��7������.�N)����9_���}}}��(�جb���{������������V�'�	)��1��d;�{��D2�>GC�����D���5��ђE	&Z�b�H�*���'t�"����G���F��{�9-9�&n|��'�y�������_>���+C|{c�{w�q����p���yf'�Z18t�?~	����??ǥ��<z��Y3��NI�B	�z�rz����3�;{kll,j�Gsg'�X�>Ts��Ϯ17�F:_��i7SQ@�r���L�e#'�P���NÃR�|b��O�����d2���!W���Ͼ`g�_����A	��Y���{|v�;�d��������Ϩ[V�sk��>�^�B�����L\b-l�ޟ��)6��>=B~mZ3������d�P�6=�'�����;��dH�	�g:�����K8=a��I�J >�W_P�L��F//���f,�ܞ�������FQ�[��Q�Oms���guu�r��!�`�v��q��\�s�������\�9B�$Spb�u�#�3)*�uJ�e^81�Gocg5����������ΞVn29�[��/���C��T�|���=x�I	��Y�`F��[�9�o-pt����u��� �]���_�?E"���&�����~WP�_�V��铯qXl|����B6r����e��|5���I)gS��|��|���n�Y_x���+lNޥ�7�Š�	�I��N��j�X@B��6[���&��lR������Bt���;4[4�j����tsz�CZ,[�R�T�F����n����ܲI�U�j����SJD������7��f�����k,/'�XC�Y��\�B>��f&��>�8��"o����%�ݸIJ��>?���9v��`�I*Yc��"7�M���Ijfk� �=ib铁��l5�[_�9L�6�I���r�� }>2����٧_����_�Ϳ�9*������l�Ͼ��`���]m�f�ج[\lg*\�����e���
W�c��hknR����S�&�H/?gk�	�6�I�q����/�5E1: c���JC�y��H�I����z=�ݻKܹ��+@��ĞNh�w-�����79?Ԯ�l0�"_)����X�]2>���R��d���Y�X�p�A��Á�����e=[�Q$y��Y@5�▲�2��֠��O�:I[���>���BT���#�L���Ek{;m���f$�4��`|bI�~*-]bB�vj�0B��d���b�*+M8��I�e��@#�O�㳛�`n&��O�ĩ��8wz��\x�%������=��p~@��b��A\���?���8��-6�)	��K�^'�#�[���^�ѕO78�L<��\4��w�H�I��A����H��2��G(3g���{}���d���wv���9��97��h�D0��ΐ�G�e�\v��z�?���Z�lY��q� A�$r�F�s�}s�9M����#��{�{��<�g"���Rm:q9%G��i�h7���R�Q.��uq�� �Q�U�TF~�r���4�O���iQ@����x�<���n�����c|j����)4t�P[R�.�[�*r5�ؕw���������v���7�@p����L��`��nZ"QZ�vb>��:�.0>�@R"�t���k5YH�[E�*�F�Qxe�5�0�s�H�}A]F޾=��[w9�ۯ�$�ż.�����Wo���޸p���ۨ�0��������M�b׬���f��#�w��a��Ϙ��=�j���v��0����"��A|�A���Ļ�wc�y��kT�����n�z���8���7�����V?��O�j� ���n���$�2{9u��L��������mW�H��-�뻴���v'h�������dy5O� �Ƨ$W5{�Ռ2ɜ��q�L�j�!�r�� /���R���[4��[�ZK����1��E��S9�vX��֥��'�^�Rױ��/U�15p��?��%�Guq�XD�����n�~�I.������uw(qRT`Q�r�wnߕ�!��SȜ��e���G/Vu��ȿ� �U	���-J�}p�;�|���(MTB�>�DH=K��qj6��o��<�nM�Te)W��MUΝ<F�ib��m���L�'
���Vˣ��$�	/#�Y2�
f�V*j��ƕ6r�MHT­�޶V���|��N� ]�Fڻ�H�K<��$]��J,��A\5VQ�*RW�O<����n�^Ϟ�P(�)���@�V&�ى��!��w��/��V�.������>56(���f�L��Kb�B�����Cq�N+N��JW�|��fcϟ9J�(p���D���Ns��mZ[b�:>��4Y��B�i�1����Q�u<���2X�q��7\��(o�c1J�C��݋Q�%��!��O�j��a0�yO9�:��)+c��Ǐ��۹���B�'N�j�V��Hb�Y�Q��(�u��m!�B���u��
���:%�?�Ԫ1���>�]��f�d�)��;�}�� sK[�ƋrV�)7��ªׯ�V�T-��y�D/^���g,,.����t�u��uA/���4�R"�g����W,�v+��`�/g6i:���XEf/�i�{4np	�V���<{����]]
g�3���UQ �6�O̳���6�Ύ��d�`�X���������^�~����Z������à/؂� ��v�2(�e"�^��f��>�Rf������.���D�<+岨nu}��o���ݔr�l����ڎ�\!��bs�0�m�y����>���#݌�@����X������P+��<ϵg��,cRD�є��2��o*�Z�F>��)z[�<����'��#t�ќ\W���f����x6��f�B���H�!<�D$_�����coԬ�Bz���S�[uԟ,[�r����%�;����u��-�Q� ���˟��������C�cAJ��f�dS���W��N�JC�J%�+W:::�~�9?���鱃a0���D�L��U���%Jd�m"�'q�;q���$/�R�{$Z���gX\������٣�^%�J��|�r�d���w�82��h_TU� HafWw�<�<x��+P+�y��I�{[��[�fne��/�v���v	�=N�d�Ґ�<��XR��G%�Ʊ�v>��,�\��~��˴uv�=�OOw;��]/�L����6SKl��Z�4{i�T5�ͅ���,+I�,�C���
w��G;x��J�:.����2_|y�l��G���@�ý��432r�(Ų��?�C��/��ְ�B~O-���W�|��#�6.N��R�
ݽ�D�A�'xz�[��i$�*]J�L��>I���OàOz-{6�1I�^�����[���]��v1Y=��u5_����@-���H�r����t$|��_az~�p,�y֩�e����A���w��IZ���	�x3�����B�ɉ��1�B��V��Y2Je<�v���y~�O>�`}���>��d�A���m�1�����:;e�ie~9ˍ��X�-��5Q7���S��r+
կ����c���b����e����ß�P�:�|��̥o/�m�/��jc2V����a�)5��K�lm��`o�r.�*'V7����z��f���C��� 6Q����8�f��'OY�z�����C�n�h����}�����Cm��y��(Y6d��1ի����38����SS�Ym�%�b�%RS�I4ղu����_�'�����P�J(�~2IKK?��Y.^^���qZq~��sJ=������S%_��m]�|��I���5�3,���gn�Iɖ^#sU����:?{�4mq+7���ܟ����i�\��P�h,�К@�K h��6P(���U�=_#]hRs
�ޠ�D�K�|���PlTv�4
k������f��]����w�����pj��(F�;]؜v��|��k�8�^~yHA��Z�P���%�'I�܏�e��`o�*�c��_���\d��7�F\�n�=��Z2�08M�#�?H�Z��(ig�@*
��D�N^~���[�O,Q��y�_��E�})R.=����A
�=��Q/U=+�Jt���қ�x�4�����}|��r�����4+-�/H!{�ο��'�q��⡪�M��T����Wʌ�X��Lln�ћ���q��]6�2������7r��}��{��>���L)��x+���Y�j��	�;�C�2W�_N����Sԍ\f�D,��s��X�x����)������>�ZI���hz��W�s��o�2J�\Q+q�h��r�Ѧ��W�A���Z0깤-�#�2���_0}W��m	�X]Ygnv[�[��6O+����jV��Z*�1հ������Ϸr��
�ˋmN�U+6�[�d�C��GZ�6FzC8��5�y|���+uOL���C�=����SY2{��w�S/=�--}tv�2�|������U'q�ĕ��p�͚9�fv82�ƛ����7p�Ǜ�R���vRU�P<F�-L0`�Z�l���f��uV��(I'�ͫu�,0)��J�Z�b5��X+�]���}�as��/q���{۪n��k�O���<�����4�{��q�N�l�:�O�Q5�u�g�:��X�U�_�ĝK��_��Pϩ�S�x�$���uX�� _�'ePv��''˖}��KM��n/�+�>W���X��O(�)��k�q�X7q7S/��������3��b��3�Jf~���Y<���b��1�W𸤃����7�|Ka{7nϑ�הR��'�4�V�k�ZN�8v�H��������ac#���HN����3��R0���W+���$oq�J-�8�D�:��X�T�+��A�.=���%�����|.^9?��s��E�RU���^���o��G9ylXi�b%����4�������[0�e���/e�SFM�&��#��v�S�:q��ZbJ'��N���l2T���Yb��,�ek�XwQ�����M,*��j,3�Ӧ
��w��{ZU"P���f��	Fە0	��GB�nr9wI����~�J���������C�(gT��h���L�2n��S#B�8��KKx�A���@���V�69�W��$Y�Li�G�gR�e�9TU-	��$4q?��I�&>�Mi�vC���v�:�l*�w�=fk'I0�ȑC�1��<lv�Z�6���OWW�l���:/f���/`��T��!Y�����l�6�v�M76K�=�U�¨5�d���AN�����&w�=��R���vPK��"�B�X6�����n�=�X*���3�	�.+�+;�m��x}l�-�x���vE��+01�B���<�kI��Zm0�\]STyU_��X�����H��[7'���]�u�fx����a/mј�ղ�����m&���&j���Vs`!F�rP��Z��)�\�{�+)�����a��M�X��ŗ&���o>x��H��]M,�+;;����6��7�������𱸕�ҍ1�ҕ��� tuv�O}c~������Կ�&is�mi��6Z�&�2�=؆?�B�R�8%!���r�?���X�/����h�a2��FP����
fI�m��2'Gz8=܋�Qfek�j�B��dqy�'�B-j������8+�T��@�Ze)�����0M� u�7� �,��VCk� �=�ZC���S،>��k��d{Q����b�D�T*ff痘�ϲ�Sb'�P����f�P�j���Gw���]E
�u"A����t$�x�F֗K|��Wd�9~�ɯ�=\�q��c���D}|s�*���&Q7��0���cj5å�H�4� #���e�����T�}r�[6'n��e���O�`b��� &�W�a��R�,�L�1�_}�v>�x���k��y�JU�c��AC�v�mzb.��v��*����9m즳��Y������c#=x]~2y�aj 8Up�M\n7׮�T��Q
35)|5�b"߷]�����NJi���?�	���ic{�|1C,桷����8�����S�{<��eu�D�a�!�`�,iׁ��#���<N�TH�U��ʅ��t$B���lr��EVV���/?%�sc�ϸ� ���Ͽ����M>���(e�:�I�����08���b;�Cpp��6:��^e���'��_�ds�!���FW���ї)Z�0�;	v�)X��V�*��bNq���X�d5bs
h���U�f S�`r�q��RI^>���G[؜�����Q����j����_�̥ˋ\�q�X,�[�9X^_bssSm<�=���� �i���wI����^��A/����El�2��6S���q��wo�aeu����G�}����<y���P
�������n�Ny'�XO2��Ó�k�
N�_��B��P���r�K�(��2^G��_=ʱ�	��V��ϗy���9s��J.��WDi�;�\����p��GO��+�i�M��<�����mO�R��t�U�Vd��W����o��~0�=����y6�@6U��>J��iL�6|m]X�^�����ȧ0�r�|V*�:l�`1�ݿ��.�q!7
�����'�[������tCIr�vrŜ�^���l��⫫H�o���'����B��;������'�,���WW�d	��buS����ۭԌE������aΟ������k�Cw_��0Ϗ����E�H��1w���=�:�e5N����I�ߴ1	%V�C�(�VT��*�BJ��::��'���W.��F����X��Y���ns��eN=�߽�Z���Ɏ�e���6���R��V�*����Cg4���s��S�/S��I����ao7ɢ�T�q<�\�6"��z�z�4쒽Jc��T��qX,�����O�[�ke@&�����s����&����(o�g��2��+���Ù3�x<���G�������!����xBfoG�p2D�>�2�/��L��OH�d�����f��V�ͤ�{��ty�~J����+�_"�����ޣ'dkuں:U����j��`�Xfv9����B�ɣ����U�h�mF�^�y(Q�J���̫F���X^����8�;�u�qx��ځ�
�%�ݻ"x��	�pl����0�C�5    IDAT�{9CV�u�a�U���%n_��*��FN!-����K���j?b�H=T�zM:;�J��@��v�r����)5>W���\CV��{-MΝ�-�`an��=�6*UlfGGGɖL|s�fW��9|(����\F{�ŉP,5tq��U�?>��R9SɊD�?]�I[Pr�s�s'���p�����={�Q԰	ͭ��l���y8a#�s�sd7Wbe��v�L2[$WP�^�!K��D+~"�[�E��� 3@̿�b>�M�n���[�}.^{鰺�$�+�6��Կ���ݹ��Չ�ÚI��J:�M�ޤ �Y�A��BG�K����������-ʠtX6��l��9E��%�W0B�%��D����$���Vp�8=J j��Iҩ2�FCͩ�z�,���&�Q'�q��o����)�|e�TYZ�bne�@(̉�12����  �|7#�Hw �삜?RdK��HI��KY���2Ջ��u0<�arb���=��z�YXak7���Q�x��!v��[�긹�O�,@'��|���鄖6����`����Vq�w��H�t(�w�~$�y����[�Ddqfs�y11��08@O�����S�apv��d^{;%fdƂ���%��_��f	';S �%��U*��ȼ9z����'�<z��믯`0�0�&[�Ff���M$��jn�����.N��*�kewS��b�'�f�_N
G4`:�'/�v�H��|�W�����6��&����ڑ"p��\��%7���㓟�����<���3�m]�d�,-�����A���xf��"�&wx1����.��#�Q�Ӳ��z	��H�ֈ�"��"�����Nfp ��n$�i��ŋl,-�~JBzŪU��Ԛ6S�p�2�F����Zc����$�~��\�6�v�N��U����4j�������K�?)�/h�W0ג�;$yMl��V�N��;>�+Ԏ��W�<��<��.]~~��)E�^��:MC�fӥ �6�$�f3�*dg��A{ȏ�R��a�6�*d�eb-ƞm1�d���.^;�������ryE�
�	r����x0��gk�j6��I�G�����L��˥�&�5��7O���ʥ�Z���ɂLwutjǑ�#��ed{����S�[l��[ݘ\J��V!�5�:�\N��[�H3���t�9��i������>��c�-�����s��z�s��S����-�cn����0�����+�Υ׼�~�r��."� ��<�s���.�r���&z�h�q��~lN�Z"�*�f�����e��	W~�B�M���n�҅2G�B���夔�`��Ź��bK.W�K&� �A$�P+����_\������z+�In��Q�8�ZE=��#C��Wo�íenޞ�l�Snةʆ�f��ljv�"��R��/�~t���?���=v���V<^����X�&�a-Az;�S�Z�3�|���$�Z�y�/�P����-��BQ�nB(n�
���9��;}��~�H5����A���_��S��l������[VVW���1<�P�[�b�M�Q���Z��I�pv�*>�����b�>gc�#���0�A�Q�J���(���&����q8�Y��:Q���D��N�R#�Ҋ�m"���^�����k8�	r��R�W�pr0F�i����^F�rm`5��>���F,d�ıa�5�Zh��X2������<c��z[�v�-v�V�Z�u[X)$15
���)^>�a���|s���!�';�|}�����P���>A����(=�1��a%�9��FQk��fW(d� Yr
'�H��>+���t(;vd���4�/&9}lD��r�IF6٢�p���=���Q^�0D)#�ty%�Z=!��S���f���W])��#�v2v�vWg�גܽ�����3s���+��F�9�3�C����u���B�eaT�I^�����.�U�ll�X�]do}E��p�����)�~�$/�p���1V�j��,?��{��s�NM�s������$bf2{M*E�Օ~N�o��d����
`B\.E)�2Z�;��9̍��%�~>z����"��?�'F����_���x�+��Ӵ:���n��&�K'x��a����XكGϲ��*4� �U���Ea�葉 ��w���.�B���(!��'�(����+�?��WB�о'v���?2�ۯ�P�jj�(=�v�m�4:���NzV{�a6������L޺D���/꣧��\��z2C���­�`?�D76��S�)J����r8��XP��R�Se���&�d�L���*��O��aNv�Me��3����a�Ci{{���G�7����fXO�-����X����5����q��s+����wd�`�L_]j��&j����u�y�n9���5�1�=�~�ʍ;XM�8=��@����19\T�� ��Qds�@�P���( C�A�ue)m7�u�Hm/�1f������Q�?bgk��C}�t�a7�)	��!=�F��{D:��̠P��H�R1��@T�h]�A3�J�~Y|�+�����Dg1ʂ�Y��/�aڏ�L��~�-1}nd�x����B5'��&��6[B��05����>5	u����=ʩc=����kG�PG E��]���baM!p�Q72$Tp�7t8�z%2%��{̯lS��jG2�F��b��׳Mh��2�B�sG86`nz���G��������jf�h��0���4�����굓,Xܨ0���V2����e��Q�_��M8�b�faK��--�
�y��1���s���F,h��R����{$�!��%B�Z��apfq_��à(�e�u%ڰTܺ|�+�����e����I��C-n���D���;M�(��,���-k[���n�(��IlV�P����5�R���,���S���Gz4;;���`m;��P����FI��y:6Ffo�é����N��az>���֐Ȓ]ħ�A摪~��{���Jp�P���3��YN�>�3���
[;�^�Ek,HW{H��{�;���)v�%�uY��l�<�d3m%�{q@�]F� ������evn�J����!�^�27tepb���U���i�QW�vϊz�b~�����IU���`FDV���!��h�q�vcsı��جL�:n���J&�I$���W1)7��s�v?5Qvl6-��V�T�Ҩi��H_[� {"������=�'���o.?!��p���;y�d���
��J�R904D��>�ݝ��u���6����>%
H]����y�������c�������Η�q�>�����N:Z��t{io�(2x~A���_�P���O�)������U<��j�]n��b��x�3������W����������vK�wU{�d�_(󻋗)�����?? �d�G�$��f�/�>d[�לA�0�"S}W;�F����U�O?����f~	KS(�e�5�A��g�ǝ��Pզܬ���ϋM.��ޤ�;A�Rfie��g ����5�]5���6Ǉ:x�|�nK�|{]?�ZS�e��}���<����_~C<�W�8C�h���P�<i�A*��w��O~�:㓻�xo�L�D��T<������4S/e�4R�,E~��I:C|��_koӯ��Vw�����L�L�^����VbA;^� V����39���fZ��v�┥U&�	�B��6Q���K{=��k/�ഘ����4�̯~��A��Y&����T��[y1�H:��_��XȡT��:��W������1����f]���F:q|.7ۋ�Lܽ���.@%��~�;��c�P�Q<�.\��v�UD�U�]Uɋ�0A����v�)|����N$��\����o�2ȫ�;���+�L,P7������{�=�_h㋋�xo��##���a6�fy��>n�C	��z�p�ϑ�g�?���S�]����Pk�0(/�@e�f(g�e��*Gz�����wM>��{�����/���.>�����`GH���C��s��Xfq��AB�jS	x�jX�fݖˢcwc��� o�6��i����*|��x,fB�A��\U�v�\�������%�]��!�ӒAz͞1�����CS�=R6����M����Oh��Yxv�FeM	��X-�g��:q�pE[5WlV��'{b�;܅Gd!��t����~��g�3����Kw)Z�,6R[�t�<���k�������)�z��r���mV�rJ,ͧ6	��.���0�7L��}��x劇�s��h�iE�MV)�mR��8Jn-�9|���`s�������)Vӿx�{����;8�A����Yhg���Xԣ����&��:C��"�ݬjh����4�RW+����g:���i|n�B�R.�G��k��
}��w/\�;c3|��f��C)G��$�brXx��滛��* �V)aj����R���1v���eW��5�����8�>�:G�a����)ԅ����(�QN+��̈[�#H��2(HL�,�Ԧ����[�����\�m�G,�}V�N��TԪ�fw��\�����QMk�Q�k�i��i��j�s����9���tI:m%��T;v]����"~�Z�zr�ў�9��i���_j��_���T���ቂ2����m�1�&�avy�&l|}3ͣ�KHgw�.}u6��zMO���GW2Kv�8�pܢZ �˨:4<ة�kC��U��Tw������/����A�}�$��T&��S��~�L����I*V�A��i� �/���#=l�Ns�d��u��Cݺ|�M�39�@�ہ��VO6O�pk��|�
fC	��L[�E��+j���Vf��$�[��F16�<�cu#M��VG���F��82��CW����/Ϫ����GL,.�Խ�י ��H6�ӊ�L��]���;گl�0Y|�-a�R�U4F,�@��K�V�g��4s��-��ۼ���N.^��J2����%]ng���:b"�vB-n�f�ϫ�=["W�k^Y "�`�Z+�� J�(�e��M���r|A7+��{��e���fEʲ�s8�皛�n� ���1�ٯ.KuQ���,%�\�д���x���ne��4�;����4���S�TZ|	:F_&�;J���-�R<�ٱ\j��G���c�5H���	�����}�lF�6K<y!�k��#$���Xq���*��%�k�^��*O�V�-DvK�Ӫ�0����^�Z�[H�W��Y!��a�
-�}���w[�F�.���M�z��R����O8�̹cl%��xo���v���Bw�y@���������3�����U�k�!��o��2hO�d�˹�Rd�!#��D����26��z+NC���уDBA��֥@C��W-L-��dr�bӢ D�5���w�Nl��.`���^���a�KO���T�^�~������r��N"��8Y�^����JI���9��5�^$�52�WK���*�BUI�cimIK$�]������B~���"Z+�,<Lf��&�`��̓�,�'1Z���A�$PG�0$�HY�7���FԹ������,�N'�31���i�F�V��U�ĭ7v�M��b���,�kiv�U��d��t6�j[�u%ϊ}6�p�h{��KX�&��� )�=���aq���%������g����P��wra������L�����T������,!��6�V�� 6��݀�!Xܚn
��2�XP�`��7����� �x�%`Y���C�v6���3�d �!c��ёs����<~���.���𘩉I�%�yZ�Ue��A��Y���e���z���ӭ&��j�]Ν��wZY�]��o/��o����w��y�`�/��e"�����3���e/]�ɋmfR�x`�j������I��֤�!c�\f_����8�#m�v���OW�Z���}�	a��t5�ec;��w�P����ާ=槚�W����W4�WW��3�#�؊Ů��u�h�������lL=��&��2���
%Lj<�jg����b�؃q�;)5��J���-�oR0�*��b�Z��~vwRT���ӹ	����u��2>�D_�U������"7n�Ӱ�+/��po�v�Y͂�6�ٯ��=���<z&��6���܂���J���&`zc�w_=ʉ�(��k�,������(��.�S�\A��*�����JW�6)�Ţ����-n=Zԃ���&���SR]��:7+�??wjT�G����Ň�Kg{�rI@JM��*���o�����m~��h�y������h��k�X�4���5&̍*]�~�x~�+B�������u�x�TKt��'[֢�'
Y�H;�(a9Ȉ%[�����6�B�bɄ��n4S�lr�P��_�cmn�L� A�с�e!�(���ջ:D��^^�$�=^�bߩ��
��%Ц�R�o�>ԇX0�KU��Q��C�l��?C5���_��
g���fjz�O~�7�����3f���])E�����u�t�hZ��,���@2��8<!�R��#�2!�9����Ŕ@a��X��[k��ıѣ�V�.;~�6�k���"�^<�o���8r�];TE��d���O�XNRs)�
)�����0�I�����ǩ�����,V*8���������n����y~��q��<x[����f�e�X	MZ�^�u��K��ϧ0ٝ��u
�5�{����zzh�E�x=�E9�6s��.w�N�H�Ar]6kyZb!��jǡI.������SR�v�_ʺ��Z�MA2�|�#���aA�����M���ͧd�&����
G"��F�����vH�j��^Ђⵌ�3BV�i��9��JA��V�̾Bb,��(t�I��8�K[̉�-e���
��M���[�Db�z�4~K�̈́���*��ӫ|{k[�M3 u��22�Ӌ�Pg���E�;s<��=��tw����;H��%�C��X"]؃��֤9����ʩM��>��m��N�,ý��?���Z���8�'�0:c�k5�|U3+�pl����6�6��%�<x^��{/�K}���2��<���od��6���]�r����X<T�亡͸��B��(�����[�x,\�t�����ӿ�g������.n��r�� �!3bpK���E��a�)�,V%)P�\��(�)ݑ���I�x�;X����dum�֨��?z�D�B����0)(h||��?����~>|��@����V��O,�~R)�%���Zh5�n%�:ǥ?���=��u�����F*����%so�f_'Vw�Hk��̆Ýu�1r,/,R��h�L�29����`+�--��x06�JR�,��)�J�]uZ"nB>'��=V�fg�G��Y����S��j���t ����D�<�.����4��-h�^�՚tVZt!g0	 L�Y{XY޹p����~G�����D:۸q��+���^7�f��m]"������3����@���9�<�&y*�A��j�z%�è�u�����뢯�Sm�����
��s�Z�_y�f)�O�^�63�M�(��PB�,��J��T�<��w������崓�!V7�G^!�}��Տ'!��=��6����Xy��1[��L&V�v�K)��ڹ��YLf�o�� P��Ψ��e7��j����].v2F~�;A&[:�A��F_'�s��i���I�C�7J<~2MF�I�O��H\��ׅ�I-��Uڢ.�y����ץ�A��SgN�+x46���2���VZ#1�v��o�;����jR��6&�C-��תj8mV-��5c��L�F�FI(�6�:s����4H;���줸{�BeΜ8���!%�$���O�Qj�hJִ~�)�jiWe�楋\��R�^�f����t�1�����"�?L�����0�
4
;ĥ�'Jg�R�N�\"�`w�d��\\�gmc�TN��$�V$�0���ݏ�`%��R+V��d�oerq���eLv���(a�,Ge�|]9���٥M����+W��,�]�)[S!_�1V+���z�S>�^��}���������i*#�z�Z�������b{\��f�������nN�3àt��4�(�� և�jT�]��R�du;��
    IDAT:=Ү�a��ʟ�z\LON+A���O+��i!ʵ:��;̮%��+Kv�#S&�n�0������-���&�v���e6�q��}N���z%�`c{/O2]��4�̈�`H�fs����=�w��Z^�n5��d����ݏ��ҵ1^LO�h���[gz'��s��K����Z�|��]�y�bVW��FȺL6���}~�� ������ѣ�����8��:d��E��!����}�����V��T���v�NJ߮[W��^�B�4j+���P��=�`O�'��SJm��H4��Bb�N�L����?C�T��_�GO"HM3u�[�-�յ163���aPzC�e�Љ�`mv��W�&*�`��a��_�'����i��v����A[��΄��6'n��l-v-lϕ*��n���gbv]��2�Si����p<N<�a���f(W�����\����3Zt�02�JKT6n
��U�8B/{2���b��U�9)�=�1�����01V�\8�ǻ�uq����^�ܛ�=}�G��{8��Q�&���9{z��!����M��7O�H�¤���/�X"�-)G&��Ǚ�O����m5����e3���o���P4�������^��>���v����״��4*9a�t'S㫫�Y��h:�F����2=����������h$���Tc�3��s�ġZ����)9��f�Ç:HD���"A�����ګ�����K2�x�T����W$��V��3��c}QH�jN,��2�b��d�[��Ӵ��+���t%���&�K�*�����u�>�|�糛��)�e�`��Ⱥ�LB�$y��c�q��Gwǹ|�*��!�G��'����Y��+f���xLF�5x<]�Ǉ�JX�~Rr�uЊA�˫%=hHF�c���:C��A�XP;��Sg=�,�A@	Vl.��=O����ɡ�.�"�rY�%��o����.-�Fy�t�ũf�,�0�l���"�S�h�0X�n�s�%�.l�<�vl����y�ֈ��_��1��漴�V�P������«�|ue�+x}~�=z�"^n/Dh�j+)�<��di/�Z*M��e�7Bo[�����D�bA2����ؓ����k\�6R�r(օ<,�&���-%i�:�D������/�M���oii��ŗ7XYY������5n"�k23[���yf����09b
�k�!��ZE�9��Z:Ȥs-��R�J4�%
j�J��K��MB~?C���	�iiwr���.]�ؑ!>|��FMa@r��z|v��� w���i��d��i�t�����[ӌ��-}]�{ڹr�&�K�_�AS����~�&#��+���W�i���g_r��"�Պؐ]T*F�q�9s�O~�
Ϧ��x�1&{��E4��o�5d�#�a7��.�.��U�L�oh���u����������j&�V�<�]`};G^({F'u�k���Wz?�B2�a��I��f�O�L[�ʝ�<�{���x�/q��,�IZ:z<�� 
,/�x�t�g�Y��&�N,7):e���*Qt�lo�j�`Oǆډ���Ki�����ΡC��w+/"�P��ċm.~��v<
 �V���M���{�����
(a�ְ(i�c�+@F
����`��M�C�Ht�H�<���a�����mi�+�d��k������<����_�*�[�9����,n����`�h/��/11���VQ����v�n���M�N��sm�r�?�ere� ��9�������p{%3jf}s�����u�6YBI���t=�d:�����ND!P�vn����Y�����+=�ȉa^̥�����E�Ha�v�E#�X-��1��˪В���FtQ"�q��!�x�뵃� ��ΪE�}�si��
�p@�Z=}jK�ܙ���\�~U��o����%W/�B]��p������Ă��Ct��c�aP�������2�4�0��a0�}��-�;&�Ѩg	,�=݇�i������Ea�Z�Q+�R��5��sp�\ܸ���-������(~�I��F��,�(��g��Y�)P(V�l���ЮYY��eQڪ�6)Ujds��(�"h�h�I��R}%�{�=6���u����x&n��[ۻ�>�N��ٙE2���:[��<��^�H�rte+EZ��ޓ&��U�j�벪����Ш�U��J��mF*�:ۛ[:DD&���'����*���Kj�~����z(�~oT����O'���j^��R�Ζ��&?~�5�u\�f�w��G����Ib�iڃZ��0��ki�87Do<@!�K*S�Xr�@*��%�t'&s���q�6��u׊��\"A�H���PkǊ���F�ōm�|J�6s�ۦ�U�$���5m,�%����)�d�7��Xk����I�R"�r�l/V���ׅ�]��s
�|�b�]�\����q�����V��n��N�)�"��X�^�x�S]�L4���/&�461�ϞO�b�ji�<�A�oGF�{
 ���	f�f����@��\*%��ԩ�z�Ϭ&)[dkxk�L���_��j�G�h|��R��d(io֡�v
��K�KN��+���Z�)aȹ��71lT�U�3����t�H���C�{>�y�kzW��s�ӓ&`�`0��$R���qyw].W����c��U>G{���:��L� D�� �s�s��y��P,Y�"8�o��������;�I\{ɺ���jw���<L��T�-�ۦd�8Ct,^�+���W~G2�$cH`'���Ŏ���fp j������?��x��/��F�/��B�Tӌ��		���Gfg��$����R����Y^Ok�f��u�m�v�/y��=#gZ���V�Მ�	��$�q[M�����ru�]|�J����3r�����D�T�*��ڽlej|t�6;��&�:I��P�Uv�VI�/l���֩���g��e`�y������I�Q"���Y	���TS-��l���m�00ЫEħ_]e}�H�g��~{��h���A���/���z�q��\����{��-�<;5��v_�HOT���i���Vy�L��"�鈈I�Fb�7�P*�A�������,�O���� 1��[�X^���W���esm���/�V���АN�v�yVv[�z��P�x�_Q�BUo�LQ��V�*e�./��p%��ӔF���/=��hH���jUCa���ӧd����߽�S�".��ʀ��	�.����|��'DE@"��5�M���[~½�_���{:�U�1��t�~<���N�fp�G�-=�f����f�K��t�ZI J�+�KD�_���1w]�-,��v�x,�ŞdJz]f���\��̓�<�Z�n���M���`_W�K0$!�������=�����u��T� ���[���������ɭ=���?3w�(/��,K�{|�ѧ:)=46��� �}��.�.�̯$��d��|	�?�Ml�&H�M��B۬�h�
%��YR9�l�Z��"�O�:�̔�N� S�b��l�?��s�ܹ�?��.�g���Jzh�yR3���ۻ����tD4��n�w9J(��֤��[fg���`{(����Z�5!��$p��/<;�3'c2i6W�(��7�jK�l�LM��&�/��`iW���0��>��!+�4J���e}}���}��5|���.��OO0���i��X]����Juv��Her1�'8��g3���P�B�8(�������!������9��M���+�}�����E�O�;6�7d![�p�a�+�����	��R��J�w�U+ �&A��%B-�ñ�ӣ��E�G�x��h����z����Cj?G$`����8rl�ǋ�\�r���N���0ʹ��Ul�nw����t�NC�3�x6&G�4�P��jz�zv��_��h�������M#�3>��̳��Q��#��N��M^~�O���F.�K�VSj��"�'�m/�X��!������0� ϝᅣ�HYyR���[\�w�J�K��&�jj��_y��'=77
ܼy�{��U��l�6OX�魮�n�~'���-���*���R
�[�}F<���߿����Q^8��̍h	���P	��f���-�6y���':B��a�]ԛ�_����yc#4G��V
Ν}��A'�L[���\e6S,�Yb����@`|4�-n]�α�i�}눒�e�-��m_}���ן`�T,���B,f�'@v��෬�������	z=d�Y�>�ע�����3L��o�K�"�Z���<G��\�8���OH�E����R�	�}�(��n>�d�O65�]TO�`8�Ő�D�L6�O�Zag/M�m%[�k��b|0J"b��i���&;�;�kP���آ�?�#@�-��d��UE��Ů���������T-��_~�@_?g_:M*����tlf�:�p�SIګ�#�l����׭������Mo�V��u��Frۤ�o��ɈX�ԯڨ6)���n�P��b�_@`a�|�ͅ_k���W��H��A�(�6�k\�1O�n�͠F[Y�4Z�ƅ/d�+��Sh*gh��1����#��~:��n���A�'���Kմh����NBݴ�v�)+|��m�f}�G�9yl�h�,q�l��Xy���m��T[6l�>:f3sӃLO�TvߨuXYZ��cɚk�B��
�;E\匆��"���ںT2��CV^y�0!�P�/���</�y���{;el���d�9��\\����&�|YC�E. ΈM�pX5�Ӱtp"U��`t�@�B����H��$(���'t�X��ބ�Z�������sx\�]-�jq8XZ�qw~���Lf*��2%�0���s�����[�.�-�2V����>N�#�\A���z��r��g��VkJ2͔J��ץ����ex8���Ϩ�����7P.J$Y�pP6�u��"����
C*uV7ˬll+��U/�,2��؎P� ��h�)4X�Ω��ْX27V�35k��U��Zad�,����	z�ܾ�P��s��`������I�PH���۔�I"�dx�����~��X�/fC��J4�m�a1)4�%�բH�x�N
ٔF2����u8th����ʕ������%?z����6���Z�a��?����4u�W�A���M�����wk]��Ͷ[3�K�������15����Jluj*��j:�����nR3tG��X�%\�:3C���z�´��IB���7����{��x�-�A/��/����Hm��[Rܹ�D�#/YY+�\��񑥊���:?{�$����o�������P���c7I��fx A_����>0�/��3��ga9K�f�l�j�d��_�:��UV�	����҄vU��ȟ���'<�j]%j�����/Կ���cr8��=��^��>�p���5�݄M�"�#�1��쭬���5�[?4��])B Wt����q�c�lV��*G��r�T?�����ͺ���Ri%_����y��3<��a��xĥk�0<}4&l�k�h���h��HX��v,���i.li�n�J^I�x�I<��Ѐ/�t��L�;�iֶ+j�n[%T�[�?�F�ŌE2-�L����STr6���L�T����S*�����hV�LM�37'q�v+�&��
M�-l���crH���ӣ/YG�hi(�v���P��6�h��j6�)T:�G"U9�@�S�McR��usm����ý�?U��p��-���ˬe���=��f�Е��Da�������_��_�N� �/���'	�G0<����z���ek�k�/����i4r]��������/�!u��_��I���.R�����e�/���$n�����"�<������:�JIX��#�&�W��
pw~��t�V�_[��6j���e2l75��>z����yB�C��W���r��������70۬�L�26ѧ1+�j���:7�mq��c��6�p�/H�T�0\
h7�*s�v��b�A�ced0���^�T���G!�'��#tk��tY��/p��5������STs����^V����7�qj��8ê�n��ڽ,߾Fik���:�=��X1Ə�D�5��7@01�H�n�����>O�ef�K�� �/u�$]
�Ս�+{ܑ@��!k�M%�O�� �m�b�wj{c���-
�6{�Y�[c���QFabwiQ�tIK�%��O)�m��F�jע�R��a8�ʕW���4sؚ)~rz����(z�_�;���y��S*�쉆0�p)���u��$%������c����\k�K��"�����|$���Ã��iVJ���������?˭�5�?X��N)�@��x�\!O>��+��⭗�0f�E�|H賛���|��J� f#x0i5uR����;�wW锶�����;2ç�^�mq��������cwӛ�hDO��㕗Npt:Do�D��E~5án}Ju�4$�J|��y�u�xp;����T��O$����d/�c+�fk7�]�nS�PB�Qz<fʅ�e�b�݌�M�yw��š~���h�����s5K���w�`j<��j���G���=���	�M���%��|�t�� u�/���-�$��M�jj����p��N�����w�\����ƽh���)�Ǉ��hQ�w�CV,W�}t�m��691;ͻoNbt�;(Х�އ�{M>��m�[s��0Hۤ��}�����͠��e��4�D�J����$�y��QB�������i��T*{���ҳxhѮ�)�tZf�TT�p[�6��5�8����Lf�����8.��j�����S)�7�����}Q�����11*�?C7��L���y��VI�vPJk���d��+��|���`n71L]:�"��.�&�>sHp�~�)�J��Ͽ�QO�Bā?�X5���ay9��v�������u޵�����2��2�gtث����zm��um�VS\�zW������J"ﰶ�����嗞"����G���_���B<�в8H�]�����~��-QY���l�F_��ٳ�'�k3�
�鑼�n� �qh<�RVSˢQh�)Ǎ�dwvj�Ryҹ"+{�RO["�7�7"��W�~�|�|�H�Pes�@�P�_oD6�a_@ϯL:E:�&[�j�� ��Gf�c5Dafh�d2jor]*�-z�^~q�h�����9��O����(��~���핸�x���<Y�vx�:}4��"��C�tY��$�+Y�e�.3�Ì��{��B�z����D�nc=^ҦP����[dݰ�����g^8��k�\���b���2ϝG�T�����J�9�7�Q����h�b��h�/M����1�G0���/�ҭttx��1�N��ׯ�)<�up�&�;>G:o��O���n53<dr<��/�� �+��AL��~��M�x���8� ���C�ur��f<&3e
Qˈ�Y�/�r��P�Xf�vۺ�p�-<��,�1;�k<y<�L��Kj?����H��!�x�
u�2u����M����	�ũK5�w��&[G=�E"ږw�A_̋�핕$����n���M\nC#��r>:U���R���%���J�mԫ��ʲGd�O�R��n��	rE(�gS�;�[�nr�?D�� ��Uݰ䵜{�i����g癿��GH�5��.�R���+��������M6���Ӹ�S�ejprz���_ī�Y�m#[����V760��D��nI#�8���;�N��~����;�RE/$�r�y�fS4�����)b����ʜz�.\��wW���o���S��߲��$ޛ`zj�xo@���L���47��[��q��D�vZ �Xh��!T��Z�F�@0�PY�����٣T,1�?��`L�����~;՚�_���SI���+JhHE��V7���^��N��͠�q9�t�u���k%�k���W�y|���kE&*Mr{h���/�8B��k7�QgV@0g����U�>�T�k��Ю��*�x�Y��Mq��#�����ɇ���X/#�b=^��y�������](8:�:~d��q/^�d �ؗ�|����l�l�>� ˝�V]5��I    IDAT#Bd�Эwp۬t�i�}F�ӿ?��+���l�l���/��|銂1��Ɖ����M<Y,��7WȔ��ZV�U3�`\O��H�,�	y�$6�T���9L�q���������p�G�J�q�<DBfƢ$�n�&\�x���M�y�,��!�D(E���k���'߱�n`�F�	G�a+e����x�,=��%���PV��P]Cs��<�?>���Q�F�U◿xE7^��3R����!�UY�z�Ll�Zx�܋#.>��e67�*o���0sa6 &@ٿ�t���R��$�I-Rr�6U��D�r�̎X����lﲸ��N���V��м�A��N&�Y��l�L�ۑkP0�M��MEx��g�9l��7bgw���{���8k+���8v��O��u?̓�m��2U������v��j��x�*a��@�*�x���lb$N4Ҥ\���נi2��Kr��#��:�ljz�ƉD{�u������K<{dL�r2���P����K�`�UY�Ä�Y�ҭUT&���er�����%�2Q�Q&O������W�r�ˆ��(�i�i֓D}6��#�z�ģR�^��,��Pi�iv=���T�g�Ici�p�;���9qx�����m36���)���@*�%�����yu{��׋�a���9��8�1�b����n*@�Ӥp���.�_;�������99������?2w����!�xp�\�����K,��8�؜����I����VK�0��堙m��L$��7Fȥ�l���l��.w��v1}�0���qO�p�;&O����P��/=7N�c���:]C��[�ϟ^� OX��L�6��-�`v{*;\���C=?>ǟ��5��P����)���fMv�P�o	�pBA�Hȧ�l��^����6���B���)�bj�@P�A����������������x9�>3�e5��{�<3;�Po��C�x�f�.��,�����}2��*g$Id�2Dj<@�a�6!GW���^?���0{e~��_1;{�7�>��m�������;��(�vu�%_O������o6���V��.�c�;3B�ҥ]m`�:4D^�q�L�)՚�{bT4{o�J���j�pʍN!�R?��O�������	w;|v����M&�Un\,�x���}��࿰r������)���E�����:��0�ѧ	�M�
'���ѥ\Ibjd9<c�7�P,��c�|}̀��$����-5�:��@^_��x�M_<L8$>��r���D�~���VZ}�B6�������`��5�dq5G��e7#q������(K�O$��F�l|-uU��nN=?G0$���,>x�駞grl�![3�����iP�plIޥ"�E�]�'b���2�m]��f�[��Ru�"wo\�]�hą�����$=�����L��ԬB�Y�U��'¼rf�X�J3פ��`u�l����UJM3&�O�y���6ܸ�w.K3��H���A�����gIL��e���0�D�^���Ӽ[�+<>��3�зK�n�V7�ht0ۤ��k�Q��j�"��^�]k�H(@,�WO���R�ٵ�͉s;����05�E����d;Y��b�t�����h���F�&�dQ]H~a�j~����K/�?�amu��?��ϼ���0�6���
	u7��VAs��V`6�;,�z��ؙ\n�R}�l�+�����a37Yz�F!+�]B==j��c��beeC�l����iPʧ��|��Ѩ�@%�Č�a��r��w�u�Ց����;���]��L6�͠��V
���aw�3}�ޙ���$	b��8(���	&�k%�	jnk�4���N۩�F��]��L����s(�1w��-���lo�J�����Vʲ�2Ɔ#����mVJ�
{�;�3B�ΫOXR��fP$������e�%��j9����ȑ	��loo2��>�H�XH ~���j�NM��{9����?�b�`sʠ��1!܋J�^)�p4���A�����z�r�#nL� �{i���E�^>��`�K1����228��������,^`yNB�~�*$X'&�H"��Q�l��_�EFiK#$�
f�z�^}��&C\��2�O��Cɗ��z|.���Ϝ�(��am#M��T�ީ�q"�?��,�[ZTV+6��g�]lN~��s���HC� ��R�E*Se~e��+B�-���	�j\�BqJ�d�H���a� �}~��1N��s��>���8~�)�z��V�)d�zㄣ�M�l�;�ָy���к|X�ʺ�p��PxDr�5w�6J8���fd(H8��.���loq���;)�;���X�f�8�.��}��ef&z�4�T�ELV{�&_\|�v�E�*�A�����`h �����]R��|@����z��j��-��ї�}����PnU	,��wgq�M��-V4���qax܂��i�R/V�z�>��EJ-�8x���cV<���a{{���m}ን�;��|F/<?�܄����n���M�wv��Iҵ�(7%O����KY�
�l���Sm�s�U��(�X��_�����?�Å��Ώ�ab,N1�!�
{If��qw���}Zy▘���0[��C@/m�6�zVj��12����`�|>Ob���Cl�'���9��H���2Q�molҩ��Ż瘛�^�R*�.߲����cY���B�lc�˧Z`����/���n�[�.�ɭj��N>�>���<�,�� ]�Jue�Y��N2<�Cj�f-���j�M�7���Sp�-�6�|��5
�����	^xF�D�/b��^�޽Gl�n�����av�)�#���##L�,�g'���Z�J�E����`2T�f&�2m)-��y��6�.9c�m%����s��6>���ܹy���>����f�޾ ��K�I��YXO��kbwpx�J0wC�Q$7Q|�]�)y�J�e��x���q����.����r��#'��dam�[w�S���s �`8D>��Y/���^��#1���B/��\�����-�gh8"T�B��tZ75>���;�x|�2���TE�M����0��9:�aZ���q�����+r�rv�f1#��.��$��W<�݇+4D��㟠&�!	��%����w��D�Nz�.�=^8{��-*�R�Ƒ�C��dw6H�o��e(V��c>���|?�����@����[D�r� ��d9�s�=^���c�<\����.����r��(�l�'Y.]�C�ڡa�cs�U��j�|�q�*w��P6^ߨ������ł����:�X��tx�4�?}��X/�@���_��q�P,Kw">�ռd���x8:�O8b�p�x���OC�n�M�I�z!����('7h�������u�����o�]����1bCc�,�o�&���a�]��T�u�/��+!6�����.�m�Z�f�FyS)�^���'���Qz��s�s��C��6G�>��mf��-�K�rY�z�;�sg�!_���/�.J~����fPH�M!�f�$9;e
�U�>�"O��ۇ��˯9y����d?c��J����-�0��ІK&�6o��I��;�ݐl�NS��-[e�<s|�#S��>��H_�p@�Y�d��~���~���9<Ya7��p�4���v�m�(���|.z#~�!�a��v��/s��c�UA���,?[G�D#�=�7����e��y>2I(�{����O�醇�z����@��ǠR�an��g�Z%�q�Ar(�D�L�ɷ��*r?[Eb�D��n����,Q�&UN)C�ہ����zHeZ���r�D-��>��� /�_|_�=n�w�J�M�XD�%���� s�M�|qٻT˻x|&�?5�Ҿ�/]f��c~����LFջ�������,m&1Y"X��62d�����=�M�v;�[�v�D���싧Tr()��rA%v�;*��� 10B�n���e�	csR�U�C���k���(рA_�.��+�m�����&�[e�RۉL�V�s��V�������G��7u��=�૞�_�2�)��t�z4�3�MS��Y���q�j��U��n�J!���!6��F���0�:����{�8\y(gh��D�ް�VI�Z%��
�_� ��{����Z�T���M9O�Ro��ϩoQ�I3�w�y��F�<�,oq��8s�u�~��%���Q*�+TiXC��]C�z[��T�� ��G/��0��ܨ�nDJ�D�˪�2�U�����������n�KT$&N;Ւ�Ao��xԭ�C�ۊ��V[\���0��9u&l�����g��D��~hk8%��!<{���	��{�����&F'O��Qot��M8���%��4�C�N���-���j%6.iz�!|����	B�c�l�l��1{�2�L�H�K<�1$�D��4�7�KQ�EvS%�u�X��H�jْ�P��Z�ˌ�'졐Kr��m�z{946�q�#*�
�k��gJJ��T��`�;E���&>]�S�4�@+�� ���&L��s�n��4�����;�?f/�cmm��TZ�|_�ͪ֫S�C����V凌fS�]Rc�J-�4�\T2&�ď��n��&��Z�����1�Q`x �3OO�u�*��t���ǎ!���L
���|��<�bS�˲v��abV\&��J�pQ�x�lo��8lr������vN?3�Hܭ�£�<y��L��f�D�!D�Q��NC�&m
�#f�`�n[+Ï^>ʋ�Ę���_��7��N����-2�.��l���eY���n6���K��dI���$G�Íf�)t��l�|:���ş4[5�'Ƶ���ý�Z��E��;���
�x�����G�^��dn{���ﱛ���Ҭ�eL`n3��U��Z�!��f���� g�-�b�е��Z��Ξa���e������G���65J�=>�B��A�U�T����O6�co7OS��L>�&���/M��I0�R�q�T`w7C��d?����:&SW7��q	����^2�'S����by�H�fְR�Cr% �K����tҭ�vuj���¡W�_������-�:1��'�G�n�Y`q5E�l�lђ`i����l6���� ��Ȝ�{:���ԸD�r��M���rE%��`-����.9�!C�E�R��0����r|ʫ�r���� _7�O�k�������[+06�K��e{i^=�[���ɮ�A�p�=A���D����i�j�	��!��Xp��T�B4��`��v���&ٗ�]���Ta�*񘗰۬�X$��i�ff7��T�si��L�m ��C�����8�����+�O�P`a���L=��mN��J(��.�!�S��t�v�k�ޛ�����Ͼ����x��י�W������}��~��N���ï��-	&�n��r9T�*����*�z���{��q/�\��o�Mo��͆�f���@�{�VX\Z��p(�TH�R�����'xz.NP�����������rG�zΰfE9,��S�h6X�{��ߓZ�Gu�1�nRe�x{�:)��m�4�J\�ʴ=�C�)�H��H�k��{<v�>�S�#��^���V�{\}�AW���0�!�F�vpI��=�|�q�j�����C�9u��;�������^�d6�Vr�l�N��f'�#�DSY.�2vd+����VG7ŻϏ��l��?��{N���Rfo�\��yL7n��ͣ+�`%��f����Ĳ���R�[� �1��f�����s)>�������/�.��T���x��īo�˥oﰳ_����thTF.���0�)g)��������� -��W��*+IV�D7>8���`��}��=�u���$z�<��)%��c�	�;�7� p)��(+]qzr�����I$�����v1[�"��d�y�N��<J���H�C#A%�;�Q�ar��I2� Wn���y6�Y&�N���ab�.�B�r����O�,R�-�ӯg�@���x�p9XCB��v��W��J��񹳜<꧔5���}�̑9=1>=�\�D�q/d�[����b����d���S1���uK$ �8�^:=���O?�-�r���8���{ܺy�ՕM���5�~�E.��_^�
+���nџH�v�V)ha+R�P��ȡݚ�n���4�qP|J3(�`<Dj�!?�k7�%vr���v�<Z�`����0}3������ø��Y"N�j��BjC�ð�d:K����S���T���mp@"��ܬЬ�(ŋ��:�ģ�Q(7�����v8y���"VR�y�w��T�X�f�&���U��/�OM0��9u	9��Q�P�>��v���-�;�`��Wo��K���p8�rc�G��$+E�j57NO�Z���p�[$j�P�ݦ��n�JGb�ZFz8~d�w�	z�	�(2d�wt&�~��X�vK,��Ab��M�m�i���B�nΌDq�lDz��L��I��q�s��Z����f0����;���)Z�0��hLr봪�DC.����n6��ɦ�j	
�:��m`&[$����X1$S��%�1��W<�]�fJ�[�|^��e��B���<��b���Z�q���L�z�B�T#W�`qx1ec�d�nզB$�"9�vk湳'��s��6��>`z��KV�����
]�˛��-n���fC �"ض��� ����ÊW��T
���!V���J,ջTth����cb�äsn�y�/Sk����-��ڤ��X�X�M4⣷?��~��wWF$�WU�"���F�K�����4���F�'B���=N��	Z/6O���(<���n���������,7t�W*7�H�!v$ɐv��m�;'�!�.�C�/��i�r:�#���t�1;��C}$bnJ���W�l_6���_��;�&�-���n�R����ܙV'�"9�[��CQ�ޔ�ߥK��ܔJHE��xa���e�y���&�����Q��d9K�d3w4�'Q"}QU�4+e*��Z�2�,�ZK�pLrᝬo�j\�ԏ�#��H��#��h��f�h�+9	��a����l]"B�}��6-?�Db�����S-�����E�L"�q�l�i"��+��%2�� �w�������ġ�~���֬�|&�3��!+�*&!��x���@�K$��bi�e���m�ʓ�}lV�A��JW�S&�����d7u3h����s��Bk���W����?~�5�d�+�v���Ww4��&���d�"�i�8YlR��$FE��
�N��ǎ���S�Vxx��v�r��=L����/�P���JX�lp*6	p5��S����f@���fֶj|����m�f����h�u���	���&{���I���A3hifSy��w����L?���m�1٭�تiT����ϥ�����^!O�ۤ�K#�^�+�~�%��b���8��{p{���Yb�>��j|��%��
�>r�$2Q��DX����v�f�_�CWaM�;���D�iR���U�f��l��Osh4̽��|����?��ᙠN��ֲ\���p�lɌ+4�^ĦE���|�\>i��"��Y������j���O^�F�X�iS����0fCe�A42zH�MRH��he!>��x�f�~fF"�z��\
���'�x�����= ���v����`s���]`��Um�Vٺ�1����S��e�"92������@��A��Y-�l�Z���]�%�a��TkE���Z�ve����
199E_\��n�Q/���r��-\;�a��6���b��+�!��$ur�nR��qy´�I�v�o Q�r�z*�mb~+?{�&F���ܽ��_��g��y�ٮr��"�W�)�ۘ�A���p��^�ճH�bW6K�Bȴ��Ь���gh�R�,iF�sg������o�< �3�p���X����lP-�:��D��v�v��_-���el��N�dj'����8�F���wX�u��G7h�/�%��"�̝��ѭR�o��Vswzo����4�ܽ���O��W�p��Ų��F:ob7������ϋ�I�U彷g�&�:�Iߛv�M�� �������/H�J9��969�Oޜ#�Y����g}/I2�e������'aRoCCj�x݂�.R(�27�O�c��    IDAT<l���U���[!Y�����*�����d
c�sڢ�d�Z�yJΖŤ�u�%y�6
�u��oЮ����	����/<�ɓG���7LL��2����K����\�6��v�3��["��z��+-�]�]� 3�\I��H�2m5q�,L��+���Kt�i�,����LO0w�0��'���!�r�4"������o񭷞gj�P��?�ꏌ���'�X��ag;/�W��ek[
��z���|��	�J� �D�;�Eb!��(��/���T:U��-^�o�<��fA=��/�vc�r˪��8d�)>���U�.f%�J~Zr�1C=���$�1+�n����u
�*ņ��7�[I��ZꕱH�/����B
�)�4p���JFX=�K������?�L�&x��K�Ǹ}�>A����.��+g�7�e~i�é��J�����j�j@`u�J�*�D��u5�ٖ�A��:��)���_�ƍ�������f��U��o�\�cD�Ȏ���"��p�)���u�̎�qd���B���o2<6̑�	kn�ͺ��M�y����2Q*�g���C�"�m4���J�HW%j;;.~uU�D��8��{��BV�9�|��;�&
53��]�3I����ެ����2L�{T��LOr��"!��߮����&�uH �j�\V/���C� �=���Y�6,V���j��B�۪�2�*��p��i�������І��s��tkk�#GN��囸}}X]aV��J{�i���!g�dz��)��I�[O<B�k׼3�]��g�z��	@�^��ןq���9m�c��78�Df^�o�):��@P=Y��N��é�L������y� {橓�M�Tz+�2X\α�'w��R6�s'g��樵��}.�,��w	�������N����[k2����~ݘJ�`��iYڬlWY��P�8i�PF�G�K�z��j70KLC�����N���Y�qsS���_Xk�E�%�fS3���2I�"�*6m�Zm٘��+>RQ��	x��KY�cf��{�*�ˋDa��Ǳf��
��8󋋌O!_lq��<�3@�-?�]�����l햆n����z���%jMQ��8��б�6Z\��c����h$�lk�����
�9Flj��3��ּn�݄���UN�w�Oע^�jU�TnU��5����N�����d�kX��-��-,R�SUFB����t��P����y]���zɧ3��)͝���l���B�����oE:-2Ύ�S)�!�J=֬eMpx�O����exx���8�B���4;�+E\�.w�ʴ�&���k�S�w��7��Y%O��׬����"VZ��IiS�oӅ�P��-�Vֵ1�X�V��D�]|�Br"��կ��]aQk.��m*u��`��������۰�fp�Vۅ��fP�("O�)��G�Q��y�.�x�*Mj�.����6/�h�KS7C)��Ho���N�'�/���b5"�|��fJ�&V�bz�v-K��K,��0th�B�ɇ�γ��:	��Ay8Ҹ�HE.���;�S��~z�W���Y���S���Q,m�6w��,M��-����oR��W�?�$�������)ct�?�	*��Qj��^���#�൝,��Q-����N���wh7ۚ��i��8���+Z���5R��j����ft�cn��ZXcoe��'7��4��fZ�im��00s���	l�8�إި�|/�10��;�J�r�\Jmr:�XMt��dog@/�R.�Pخ��Z=��"��-|~/�p�C�3�e�|�ї�?��3$�v��{{;ry�W�f01<I�i0��R���˪r*ŻSۢ�,S�D���90��y��A/�����˼��7	��ܹ�ˣG��&�؜1�V�6�2e1wh�%���Е�,�[�U5�n%���_8���
�r��PH��2��O�L�����B��퇚m%r��K��rȠ�D�cclt�Pԣ�۫ww��x���אɠU�M��	܆��'���ے3�Y�b*�dL�!1��6��;�(�ȓ(�>$��|J���@�L&��$�[°]�^����Q�f�:r�Cf� �|m:�.n� �C�x�����M_�q�3v2�i=xH2� _�
ݝ@4F��dk�D�a�����ڨ+�K<Jd�6���#.��g��O��ٗ��T4q��"O�6u���hH������`�&P(s�wi��mEr�Ef'�Z�����9n_��£;�ł$b=9r�����K/���m��cSC|z��e-�tB�Ĳ۬(a�h׈<LNL�y�d�G�;JPlt�?���@/�z��[�Y�}�fp�i��`��z�0�Ä �z���ibn8�r���k+,,op��q�x���Z�]>����ة�|ui����zq�$���+O�����q8�n��T(U���?�G�M��;�S���N��c�\��<�h���A�����|�����ؽ=4�R!y_2��&�M�-��]�a;�5��i�ޝ�?\զCBy�s�hv%^D|j"=�jX$R�:h1�Kn���R`}�����>��W/��o�rY�䳌��vL���׿)����������f	�G)6 [*@r��ikԫ�M��Ȉ�D�Y%9me0736����.�)�������C����>��7I�w�\�E|�(��A�+�zI3�87L�d�Ƶ�<zp���O��b?�����Y66|��mj�u�8��{'4���>�<�RLR|�����~���N++8{b�ىA���;�����w�,�{��o��-�0�aW9�a�k�&�nO��y�&z�xٖ;0[ЉrSs�
hrPM�[�T�]G><q�tDEl�M�DH;(͠��
��>����L�������|�+?��n���9s�ȎvS�hi4��Ʈ�Ԗ�v���/�i�vv=���㵕�VK�Nj��͜3	���E�9�s�[�{ ���REI��q������sj����:;R�3�x�|�����|ksK��Bpz}�ժ�[�,.��XR/fX��6$(��Ü�����V!���,�_����z�
t���#��*��*��^�ES��mC��∶���D>����~���C3�Z���y�q�zeZT	V��p$*��;�x���|g2����b{uY�Y��e�I��������dk�v�.���$p�W���#���YDMhR:�Wh�J�Թ��Y�6����Q�V)�CmT��ut�+�W.-
��&$���h����XgQ�`�54�Ny���H�R��>6Dj֊p(db��ߙě����.bog�8���.a�673p�ܹ��d����[{h�<�s.�8({L-gy�΀CR6�|��M��y�a�諾Vp��g���G�m� ־� 1-�� ����ch�"�F�hk��Ak��ƫ��xt�����u�ȴT�<�]���>�Q�2�p�RMR_�}��QW�<��暄��N`��ɓ'1>݉�_� ���Su!��Aw[G'����%��� 4�����GK�+���%g�J`̠��"����F�n	=s����(���!ȅ���N���1�0u����T��L�\K���4���<�&��G�bwF9��(�g!��~d�yll���ɣXY��-6�x��$�$S(7��F���k:`6�����"�>�B_{'����_������404�1 �@dt
��Qh�8!f��t5a쯡���d	D��έ�M����]	��ا,��W���]�E�D��Eg������,QnM���6�$�^���˃�׉T2 �5e�����+ۢ ʕ"�uv�r�'���� TC�<U��i����`咂˗o"k���acs_�v!�씬2X�56d�8��ujdv�z(JJ�ݤ�t%��F16ԁ��'��lJc��P*�2*5��kP*�����M,�l�fF>�N��.�c���3+Bb��� J齌����v�L<�@i=����$`�=�S�FPe&yHx]n�u�P�,��MD�iIL�q#b n(�谍Z�-n��
�^�leD�ʗ��ܑD��mbnq�x��N"�)be�$�5�r�<��"��XX3����&�99m��+��,�Bq�*�,�ܛG��+q,-5���/��3�'z���Kln�a-�A�Ҕ�E��c�*�H�>(��5R��Lʴ�=���Oc{���Bw{���jǝ;�1<2�K��C�%�w����M]1X���E�� 
���a�H�Z���C�Z ��Z�/!�`���,k3/�~9��� ��*5�M6�(\GY�:O4��Jz�a�=����V(����hK�Dv�Hd�驖"����6��5XN/�{����è�ע�\�!���z}�t�LO���#���6lm䑣V;Þ��e����P�a���g�5���hYX�m�u�q�c"1�q}_]�����0x���\΄����K�����a��&�*�u^�uh��`�%�%�$c~�}c
������Ghoo������{�D�M:��������+�`�Dj��'�1Q�*��[U���a�	l��ckg_lΦ�ǰ��a57Vf�`��%l�g0���!u-�����>&�\yP�v��Jbt����,=fL����jM�~։ե=Y��"Z��>я�X.��@�%��ְ��F��������Ex|~$�N��\8{z~���[YT�/<C�b �[G�LF7
E��l4�"�N��P�������P;~��(|>�������������"�p�YN����< y��`'��Y<�y�1�_���^?��qܼr�n^BK<��'q��������<|�*R���!|��}�rv����/V+���zvq֫hR�;��RUvp6��Ɓ�iHY9�������p�66g�e�,}E����ׁ@��^Iu��"�W�EtF��V7V�cgk�Zm�=��|�Q�_���c�#��Ͼ��q��2��8|���'���_���~��Ʀ�lD�=�0~����U'������2��L�`���!�>��B����E�}sW:*��a�����M�)�(Ww��ҡE?C��:\�k�+i�Ӱb4LA�)-���.~|�FUJ���r;)�eߚ"2-n�{��=�_�q����������X���.�s�C����r�t��?L��:������I��b����\Fy�j���o�AŪ���K�
�p7����?��+���a\��"|���#gy�=|�T��m5P��P��ē{O��ǿ��@�8���066����������~���
O�H�y����}���M(|��Fq��h�7�ܖ���YA!�����8}Dz8y�9}N̯p����-��L�&paW/�9&�E&B�G�I�6??܋=.<��0<�.�?�EM��h2K�:�^C���E�ϓQ2�R��a��N���קё"c��W?�'���bxdP��X�o�=��O*������g��,��Ȝ4�`
���ԅ}�44jUa����:=fuM��a��ma�7���G��ջW����><�KC(� �K��C�Fb�R��L&l����XH���O�څ�XY\B�b!��?~����/>�P_&��D�}fQz�a?����z�;7o0m��60<:���vw�Kn#��#��.E٧�����kk�"'��N .7�q���(/��&���yoX���TSLtw��e?g[��H��C# ��TG���S�%51�=q��KV��9J1��n2���9k����XZ\�������K����W������сgsi��:!9�%���e�WM�>g+����8����z~?<��3X��օOq���P�2X�e �� _Z&^G��q���H���k�߽zrZ���[װ�N����c��xWo���S�����}&ɢd��'�0�ģ�k���E����!4!?N�~��a\�2��tNz��Q��<�#�-61��&��X�(H�#�y�ѿۨ4pS����}M�.2�ꎪۨ�Ϙ~m.��u��Θ�qٶI[(Jn�!L*��*<�+y85G�#� �e]�:�WV�K��M�_0,U8��=�Ѡ$�i�+�C:	Tq佨7X#����]�ȴ6�ͺQC{;��+_~�o��Y��ˠ;*�`l�0��cP�1xa��c0�����O�a�ˏ\6���Ud�)��EF���lVkw�<�]�~6/���Ǐ �6���-��d6�Ҧwh�˅�,�fF�5$UB[[L�`�"@̹`{����Je�3\�y&)p���J�>TH�:م�V+�&n޺/]����R��^Igoj*�UΝ��	hً��o{�K�[D�I�Vm�z:㘛y(�ߎT���ҷHf0_Ѱ��C��G���(���W��D`�X���P4*<+#�;��T�鱒��j������$�`8��� ꐞA�9(�<4>�#�1�<�o��� �P��S���E�4���#~^~�g_�F<�G�pW����o
��p�p��ff����h��I;�ws3��lٚ����E;� ���u���{$���f��Ïϝ���f�8��E�<aD�a��[�~$�U�+fgR�<Љ^��Z����!Rʜ��`T��'�}ϟ>��_}����~�Z�1\�|��gp��4� �&p��=�u�����TKD�*J ������EZ$���6�P˒��e��ç�ՙEl/�!=w��P&3��9�M-%؉��W��=$iiD�M�.�3��p������ho�����g�����B8���/$����֞��g�aѧ��
��-	��r�|#S(Ԛ���p9\b</���W��ԩ)�>_��x���ҊXٶp��*�i�8���h��d�1=Lid12��� \���זp������m0�;�z��:TY�1e�v��QJDK�^��/%�AUS� ���qܻ�+��q��4Rm��}�쮠b����� %�o�݅�9�J�==dN2�\��uT(O�z	'*��2��*��2�����epy�1�_���o��_d�����i��E��.JL���7Ўw��R/����?���o���d����,W�'n�x�B��z=��.7~��ؘ�ċ��Hu�	�����r��ν��-�������K���������q��mDZ��::�*4\����7���0 �"hK�4�%)�%sj�Jp4+�j�DD��[Of���C(܂��@ј���l��\��iGV��S�\, �a������ e|��I)`^|���*��`�@�`i��&��F�	���Ż�i�I�US�<�9���e��e��ʸ}A@w˳�3ܬ��qj��l��].��������"�q<��N������-���#�P.�b�݁w������/P�6������j�����o��:~��i�ⓗ��7�iM�����ν��(��s�Z[G�f"��#N���b	���E"Q���9DU�YMa�(�y�0��L�U%�����'>`���)�����?�����Y5e(��W�s��!D�9X����F��s	;HƉ�F��Z���F�\�VN�����z*����p����`��/�Ň�y���_��*2�
b���%3���Pe�+d\�Ʊ�Sk6�d�Q5Ļ'2�@u����s�Բ���|��?��- G_}y��Q�(���!����ŭ�X̋�q�CҘ{�H�X$�C����-����_���g�Vw���|!��J>�3����6�2e<�+k����@�X�K
���ebʙ��8w&�ʹ�L����<��G����`+�(���5���3Ђˡ�Z*J�[ރ���� f
�!��d!d��i��68 r��Î�nPi���[�v�b`sm�����D����3"3�w4�lőc]��V���+�.��7�B��e�\//���\V�V]�B~/�BN䢒�M+�Ak��hȋ���s��W���W�<`jj�����>�˷`9�H�Bj�<����>�RSI�s��+KK�k.������F!����	�#8��a<[����R]�9�^�f�����B�$p���3ݸ�0�o��	�ӍT2�T�/��9.�;�"v2�ث@@�    IDAT�Z�(�ۊ�C�ɦ��#�M	�b�!6�
Yk5C�)��K�l�+&S
)QT`���(��D�&Hc������ Q�d�+�|���>O���������ҁ��Nd�&�E�r������+�U��B�ߋK�%�~��$�N$�A%V�n�ƳB���p������#0�	����-HM���� o8���0Zj=��'&���C>��b��t�%��d��=x��|���㗿{���4�AVFE0=�+��b����Ƣ!��I�V��YI��E4ؐ|��7�v� 4@˿H��`k;�\YA���R����	�f@5��C]�������gUU�)�j���`69'R�Ԅ���[�P���Y��`;�+�e�!i����MKP_O;��ڐJ8���^����
1�x�d˫�x����PY����]�d�xSgA�����A����rn�RF[���2�a.�G�� <Q���. �U���^x�&=����Ir���@�W^`~�)��8-�J��-b'���o��Z���w ���}��@ GO���kWo˟]m�31�ہΎ$�&���de��bq�������@�Ȭӵ�E�?sU������OA:]��^N��ꬤ`��Fˑ.��R�F5��2-=�M��ǯI��*g	;�C#C�b��8UI���o#���	bi��b�۰����N^@U�Ee����X���L�`jv=���"�����P�Hu(�s�45����V!�8}�*��5��ӣho�q��sܽ}���p��3���VILr����]��o����݅��8��՗H��"
붵����N�����-���rb}u�-a|��7Eb�rq��hk�������-c'G9�S�{C�L��K�!٧R\�(������Gh4�$E4�����'rSz[L�$�
�`w!�(� �0�^Hܶ%�Ň�Bf/f�7&� -�Ϳ��Q���͇hi@����G�``���=Q`��aB���5�>�Pʄ+��%"gjT����HI����E���e�L��u�WC�A8bP���I8CI����~�v��;�z�!�?D!��d2���!��8>���5o�}�������b�mK����1X�<���3Yh��X5JH&c���?D���?��x��r{(e�q��$N�<���u��f�+��쒁o��@:S�$J�y�Q&�1�<x*b��L�Q7����_���&;I��7�L��>�Y��+��Ry(�@.j��",�,��(x��ia|+���e-//��14�����n�p��$�>�ƍ;O��J�%�0�b�d��)��ou���`��b���
�lHS���{�w����c<�vi�Dk�xT�%u��>�԰�:}CWkE���qLL���O/cuq�lGM�ܹ�1�r�޸���Hu�����X_�9[WO?�w���׏p��OIt���|�%ق?����|y���Q˯�O>x]���M�bq��u`y���wv13�%��N�_�C�R%ٌ�4�f!L�G��6,�_:����0��)�'��r�R�"�x%��m���Iw%I(k�38qx'��^)I���WE�1}�时D��;S���&<����M�.�٠��d�	�dd�i���4L�?������*��;d��s�^_<���`�������2�\��@ʅ}g�	���"C��cm��Gw����kx��	�83���wq��S��}�6�\��cØ�s�q�$l��<���K�ț���t��+���eԋ,��ʠ���@����v��!G�|V����`�����$�;׸h�J�ZY� ����hd�x����ˠf�dSnh{�����ëÖ�V
{�����]r��J����Dz��w��bfU�9�Y��\nTL2�.��
��D�ıY,K��,�w�~���eprhZ����_�������W�#ڒ^���o��w�� *#�2�`�������=LO���V�C
�y��(TU<y��_���qh|���Nas_����~w��L	�oFO"�������]�y���%�.nsו����n,?_���3	�)�T�T��������m�ưJg9(Z�	U#��aN��-=���.U�z�yr�aa���6�O�!�8#ʷyO�[T`��*�,�>���]����3[7�V�X[M�ڍ�Pt��
J5��-�d}�	��2C>3��%Ȑ���!	�|�(1�جZ�p��^�wű�:���;l=��LO���q����4�|�&,W-��"5t�H+|��~�7v����;�TE�d�ƛUu ��ڥ[x��kx�l������w%�ģ�qx�ǧ:P)r�e�3��n���*=�����W��8Qث#��E6�+}Ȼ�"��Ҫ�
BsS"�c��i3�NH�2ZCTQ��!8DP,դ΀�^ìHc2�RE9^9���5��x?�M��=��N�S��m$�aY(�x�l�+Kҋ��3���7�ԏ�vH ���:8O)�8���9s�L���$�ˠAuAUY��L�Z����3X�x��l��3xZ���G%@��H�C�!�����.������E��@����-<z:��}�r�5tt�%�=�-	�H����՝��H���X.����e]X�ɱxe2;�W*f17�FÁbMCS��8�&��%��2(_�m��Y̸ h�0��o4��̪Z���5lЙ����r�jk�d��)Ǖ�B���z����ku�*d=גJ_�i��u:<Z����Օ���As	���Yt�eA��D^����s�J�A�@�B�TD_{
z���>�%�?0�5S$�J�m�G��@��LJ�}�����ɧx����_"
cbdcí�|�6�>}���ɇ������#ll�0���3��x��&��L�dY*Վ��v���~�6jU[����z���XSS��ه��$@fec��Aw�E�]g�$�I��th��d�`�,I�+f��g7�"葟���]WC�$�K2�~�d�Ϗ )��KR2<�!�7��WE�F0��D�c�!֦)Xx�����
���lm��(�)��@��ux�f[�K�<0J�V jZ�e�n*���a5|H$z����i5u��nq�v66�^_���1|����z��c����34�;����ԭ&Ƈ��+�xx�n߸.�t�[�8}�>8�6��2�'3�{����E4����11�rl7��q��V��RpI��r���R�,O�2M��J��1�*��+��U���P�YP\,�w
�_�g��$�����4�~^L(����f����G��P*����~�b�(�I����ѱ	|{�	�-l@uǄ'�*���,(|8�P�RP{�`>+|	���Qf�R�����<�K�Z�@e�e����`z�=��#�5W8��B餅�v�����na��C�z�����?����-��?�����g���D����	���q��,�\@6�E8���0N�:���
~���Ez��тְ��dcc]��7��*(�
Xڴ��k`nqG���,=���P�	��U��ץ���C@A�e��t�f�������0TT����	����/���d����(.���ęm2�޿{W�\fd`h�ÏTG'�Fw�� �gPK؎V��$����v*k=�F���f��`P�M4ʦDj������ҳGxr�+���D���W�����2��`Kހt�T�<�����������s��\�:&���g��x�l���+���8��k���#�<[�egW?��qX�
>;�%��\VU��vN���/��+����О��-�����HD}���b�T��F�fW����B#�H�DU��iv)rn����^څjdm�����Q��Й��1���5�&L.A9#����np@�+��+���l!r��w������oo��o���@<Ն`�S�N��0����HZ�Q�!X��$Ҽ�,i�ޙ4ZɁ*}x�=K�6冒eQB��c��Sd�/�����[؞{�Zf	�m �F�<�����A(n'*�}����n�E�䏾�|���FkK+0r{����f	n��7�^~K����̑È��ٿ���+k�]����.�ǦP�UP�oat�aI&K�3��G�v.�g/��`� ���E|k.�.	<i6x����>4.�d޼����vP�`TM�����,dwN񮱃�Il�%�oBz6�-�d��L�ʓ�TB�������;7�#�M¨6�%���{E�\���`ʥ7�˳y�*M�F��F��u�:%��0���M��7/]D!�����k��9�I/���q��D�������뚖0%_��W���"R	/�'����8{�G��+������ۙ�k����l,� ���x�:s���kY̼\ƭ'ϰ��E{�����5	�ho ����r%���'�[ڂ��y��i�����in!j�eYՠj�e$$Ƭ��td�8�����rN��C"�Xg`KCRm����BH�U�E��:��zUd�i�/�F�Hƃ"��=���cc-�h8$�X��g���r
��4F��0������x��^�b)/f�C��y�U��0ԓ���S|����;P�M=<�����-)����:dF^Ej�C��(V�Zo��hG�!�W��vq���.�k�S�x6����4B����xu�I7&G{�ۮ��Ƹ����F�\U$��` ��
���RAd��
	fp(�Tܬ��=�Z����J�:H~����\���O�)a_^%ve��^aF��Iy/����%��<���@����&��|@��d+b� O��l��6d�T����VV��[�tQvh{����٪-���FY!�Y���m��s|�</<�7.�2���3����������A���u�%�ZN#t��1�"�K��``sc�L^�0>V���ȔLQe)�bF��C�=�C$�`ue��}�X\�7���p�YEG[=]�PP�����%���R5�I:9׹��0pŒ��)[:�Ls�����]ʣ�	�\)��LJ`[T,Ey��)��bH�L�C `���lY�Kyy%��F}�Yʗ`V��{���j/?
�����S%�HT��)A�:���$Ut�&��	3X-�'̠�~��-e���$���v�OEbpB�D	v�[�`��O���X�#h��bG�c"o�t��w��'��}0����ŠiXR�>��
�h&}Z��R�TkX^��΃YDb	?2�dTCn/�r� �Z�����M�d=8�Q1�a�����n��b�f�r^:E�Y�L�2H{=�$��?�>�h2��?�?�����^:��
s���J�=Bfg��k�g�������Õ�4�6v��d1$��4k�rf֖)�M�ly��u�8<�9���Z"����4� "�~TM'b�.�C'OL��/�g�gq��5xt�&���������_~��CSx��I\�4����֖��;�"��wocss.�_"�O?���N��on�����鑅l��gNu�R҅�(���,a3S�N���1T�@���#ɇ��j�y49�#L����aJ Nw��7�!]���f���I���B$�ˠ��4�d< �X�Y�D_g�sL����,���?	j(@��;��U��׶��lYWa�Xk`kQ��W�)E<5V"�N4�">��0�V�a����^ =wVzN�A�`��B���F��D:�Ju��5�2H�|�?9
��C>��J�bw"�z1;���?�ݽ����|��g�ˏ���ߊF���}�x���t��w�R*���F�½'�x�tN$�o�q�=��U����]d��X[ߖ�=�x�` �C'�}"�L �è��`�	V648�^)����$PY�TA��6p�#�J$�:��QI��&�yd�< ����W�ɣ�cwg[��������9.�ޥ�/���`YD69�����Z&��9d����'���T�ǧp(&\ä�:�<�wstb��C<��{l?��fy~��
c�]a�{���2���/~������n�rz ��U�1�SEk�E.�/.��WW.��~�^���>}�G�D���]O��4�˕�/Zh����(�����fW��(�v�0��=�jU<�����c;W@�Cf��=��텥ׇg�vA��wtydd�R-�K/�ӁZ�ۙ}�<1W�ebt.zИ,��`$ͿPF���A9�+��*�M���bb��=AT�%�B0#	a{��k7_ ���?Eհ����\^�$R�X�T�'�f�R*>����0�3ـY�GЭK�bT0s�.�����C�e�ܴd�3���>������B���E_e.������0L��.�r.EA�h�UG�D6[�ϟD8�����Fp��4Rq���(��kf�s�z��D0�,t�0=�.�J�@2��w`���ջi���}$;O�%��00�Q�/�	�GE�b}S�L��8�1�n���s:4AL١E�[�^��&��%���x�9�2�͡�V�٠L���/�3��J��fjH����0֗_����[����ɠ
�=����
J�&B�n�MT���UE�Z�ҭ�_\�&�FƄ����6_"��p�_#��bp���m�:G�u��L��>o���>o�oBm���Z1+�Gc�de�5Yr|'
�mxyѲ^�߂�I'3��������a���P�0������.�VҰ��4=��ǉ�Q�}���
v�Y�CA$R���%�wm+�\�W[�?e	y 8Ɨ�2 �)��
4�pI��&Y5.�0>ɪ:u.zM�|kuS�X���x2���R2��2����Va�˲���YQ����
�h]����^�wϽ��1���_��7�ރ/C��ˬᇦ��h�EF׬����+��+�e��z[�^z�����؟�/�Ʊ�"Gv7��x�ꮄ,�c'���R�
y�7�ȯ͡ի���B$� k��*�!�ˉ禒�b%F�"���ʹm�":�^�w#����n,m���j�E��Q��QޞJ0>؍���C|�Xada~is�[RG��bb�X�!�����L�f1��n+a��ل�ᑥѨ4��d �DVՔ�F��! ��B��dr���K�)��\f�����Z.!��	@�s���a���u������]d"M��UT��b/��v�9��v�:�|�2�{�&g-8��4�.�wn^8/2�M�D�������Z"o4�����'�R�����m�s�t�Ϭ����DBA��b�Z��1 �s���m-A�#~	�S�M��[bi`Ջ��|���b_w����{�/��̂��<�7�Lb�F^�
�Q��8����=U��A���Ʉl�³
����?sZ��3<O��?�mDyA&H�êW�rіB�����h�gU*H���KR���ۋ`�K���I��>cdm�r�"�+A*\�x�k�.�`?�6���_0@�0w����9������qX� \� �mII�Wk�H4��$�J����d��߯a{+��O��8rlX:�Y�N�@��"I�b���G���C���A���t���@$�xċ�ύ&�s9�vjbs�d���l�I�ڍZ�)��L;&�H�F�>i�Հa�d�����B~.�me����iw�Z���� �7�����BQepV���~'����!�r�\$�^��v[�(��ڱ�?���y`Ǭ�=�$��TV��Iv� с�Sw���=�|4.��Y��d۰��"�<^j�,z{Zp��1K+"׈EÒ&y�����9��h���2<���������á��3ľ'8�H(*���>ċ��8��+�&��6���V�v`��(U�؎2�n}!1=�)<vʙs.y����q9��g�E���Q�f�����	�s�,QdE ���>mL���M��
�S�d0�߁������$�%�z��2x>����]4uj��Rw����䌾� ��A�YTJ�� ��n5�>4�����T�9,?�Gza;`l� d�FV$��kQ��~��D�wю~4\n�2�$����Q$�^�pp;QG�,    IDAT��Y\�qs/�ݝ���C�]����e(L�,���a�#��G�QWk��4?����������j���3铃��e�5�LW��-� %.~���`��ךt�ymZ�H5�������%��E�?3>��9y�1uReb�"A|.8��/ȃ�@U/�Sy ��m��	U��ۡ�N����%����B[U<~4��L�p ���aT+�~7�.J����pѷ*v�P�ߠ��>�Uj͹�XDe�wu#�va��#<��9v�]G��	����u4~��}���~���ɠt�e��	��­:��R+��e��
[�M=}C�ݸ}g��5h���]8���t���i�[�RHL؋�x�|��,�����{�cRh^/W�gDT��{0�FF��BU��k�I���Sm�6��a/PL@+��"�B�ˬ�}`u͉��UY�حE��r*��/���e�fj�=M�@��H(ua�2�khV3H�D�՞����(�U��o�˸s���Juw��\���.�x^nDb��ɰ/��MU����3ڛ ;0�ffq~����>hF�o�����^x(!@h�3h�8�&_���AzU6�:UK����¶�ɛ�B
�9-�(��ZZZ16ކ;��x6�������u�]~��lI$/�|��@8�ޑ><��ģg�ƿr��a��|6��P�g����ś�S���Y�lf��<R3B��b� +q�fx<��U�����%%B�^4�72�����`
%e������Z��9t1�3,A�6��lfH��%d�Y.���(,���߃raM����y#�~��$$;��v
X��#��T�%�)#���C4H�P�Z7�TL���7���_"�������/>Bg��Rn�#�˙�'яxg?T��hH�tUY9��*����;dy!@�z1:ԅpЁ_��"����c���m0J��ԉ�VJ5�� [Pp��"�=s��~��oe��r�x�:�:������s����h�^T�S�����\��ɀ�a���"U3^��~��y�%�D�-;�Х�'h�^��n���>��+JU�-�)ﭢ��s8�3S)�E�H�T�΄�j�y���O΢�����r�<z���ц������s�/4aY�_g�b�S�=�QG-_�A����}��Y�����;��=�So����n��l5��<1���A��1h��@@�:�hF.�#�/s��� oQm�d���H�����B&[����-?{Z05L��S�����ҹ:��o`'�E�Z��p�'�X~����Y��s����f��Q�iv �I�H�&@�{�QJ	5f!i�7�
K��B�T��J�L�ځ��	;�о3!â0W$;��R)�X�A#�[��������m�y	�X�|��7}�l�y����s=E8چ��!�-�#Պr�(�&Y�E_�]�@u2��;:�\?�ͯ~�?.�Z��>�&�GN�=���qh:��}2`T
p;��#aG~�G���?z�[
8����l	�<����!L�&�a_�vZ��]E.�A[{:{[q��w�����	LO����"n�~�-+�0Z�h�l�܌ŕ5T�n��r2�*
��!ͥ�J��ù]�S��I�2҃�����hN��f�@j���d{�!����6<�Z)~~�JE�5d�	��	m5�N�������/��t�{b]���&��M��eQ�p>;	��kde�✃�,��2h������_�2�z:��\S�m���Ga��p"h�?����Cԣ��_s;��P*���k���Da�:�����B��f�T��1a��*�26�3X��E�rIe�ھ�8�!�$��P
� S(![lb=]�n�"i�&��ِ�bV	#����g|��<`�hq
�<��&{���B��E����n�0$��@"1ҡ�Q�a����:
�]�<�|AyV��,r�,��,AB� |~\n'�wK�f���Z�V�)ֳj� �3�6(X��a�t����%q�?7M5�h�Mx������T܃����׋ގ�a�ZX�½G���ˣ����x�0-K\0Gfwa����G__���қ�Ng����|�.���Tɨf���}:��cI}]����Sc�B�C<�� r�B�A�IY���V90D��K7�g�f	�ذK��
�֚��`�͜d����f��6��e+g�Y%�'C�kC[�-�*k6w���&�|x��@�!��4drpx�hh:
U�N'�+�{1�Ŗ���S�1<<�R&'����.>��3�73�j���+ah����B���-���~Ev��x]�=@"��5lG/��g'k�z�uYTsu�Ah�P�"���qazr �d%��i �]���.��XCK�E錬c���)y!����T�/��޳XZ���O¨�1��s8\�q���?;�̦Y�1�˃����`�l�
_���#R�5�Y�K��ms��P���ɵ�/%7I,��B��ށvTke�(���hu�ct��:�0�%�V|����M/Wަ*T�%��v��<�I�ف�σ��G���y�>�*2Q���>~�^�z��;�&��h�Y m�����.��qDn���PYx�|F�r�(`����o�U\:�]v:01܃��	f�f
x��V���x�H��.|�:�x�z{P7�'H�a7S���"W��8ES�r�DVI�!+.����L��	i�@�RF�a1��Xc;���5��o�gX��)+�wM'��'��a�߱��U< pĈe"ԔB�&⨖�H�=�hC��`g������Jpz���{v0R�	��Ah��n2z]��R�CYZU���(��\���ב�{�z~�
v��7���a�:'�� �: ϮrpI����\:ܪ��	h��`/<~�f��6p힉//=�Q��/��_��8n^��o�[�I�+���y����Z���/�xpdj^�_|����p �R��/p�;��o��w���ѳ5�t��|�Q�x����`P�R�BV%�Z��#��H�H!5x����]g�qy`P�E��J���g�!�^��Ծ(LL4�s�A̯�4Ɇ��Q&V�_��h'N�o?�,�>���(��/�l��݊t����dL�e��&�3�*��#�Q+�����n���<6��/��ۏ�;B>p������q4�ID"���F�5���`���FyZ1���	g��RKK��y�E��*�G�׿�Z�Z�ߋ?��ga�������D�����{K�/�?8'U��O_`mm?�ɏ����kl�f184 ���9;u�OOH(ף��P%R3x/��{���J�F�eŔ���O$�%�t��Q�TDv��m�Y`H<�al�HǄ�e��u���6( �v�	�a�/��Y�)�t�R�a�w������W�_��;���~'Ob�e�j��6�{�����θ:�A�����oX,!�c��{�������gw���Cv�F�B��܇�O"9t��q���#v0�YD�Z����[D�Ȣ�#��T
��"".<��������������`�*xx�jU�fT�d�8�������k�.�}�58�����K��zZ/�L���9B��싛���<�A��e�A���j�v����LJnҫ�V��V�Q^�H�9;q���bp_h�P�Ae�d�&(����*�iU�r7,�G�K��^;s-V�� �)�w��5��'����bՠ��¢y��\qy#��_����n��*�}u7�3��J}W:��3�nA����>��3C�3��r���Co��Ĝ�vk���QߋF=�)nY���E,��X_ߑ(��_;����\����4����e�7qtro�3�������s?v�CQ|��M,.�I�?+!
�"ƦF�����Klo����R�t�C�@)/i�Nk7Th���=Co);�������*"Մ��u;v��md�����xމj�*�A6$*dqaa�e��6��{ծ�2JY�zz�B3ϟ"�L`p�no5�)5��R�#�גBKV�g�)������V5�ͧ����k�@&j��B	&�?���	4Q�� -)�C��4J��ͼ$(Sr�eײ���&�� |!?�^�wL���et��0:Њ����b%���:j�K��ˍ<
�:���ו@n��}��^~��{���W0;���o�;��a�r�a��_��Sv������p�r��C���:?˪���!8*g�J���L���J��+uz~���ғY(0�ցF���#�7k�,�����N���%Hgv���-x<�P� e.��"Kh
�[C���j%�@{���e�o���G"��l���
���q;"�uìW����6[uY0�HӺ��?�L��p,)��O�=4���82��t�%����N��h4�F��X���O��K�%,dW�v�by�{E
���"b���>�0������I��r������|x�����l���F�?еvb����j_w��#�b��$��Z��LS�������]��X��ͺj���7��~I���Lץ�X)J���Z�IS\i�g�� ��<V���`��CX��<X��2���a$�_A�{
�XTb�����R�}xt&�P*�d�c�9� G��r����<�5e�8>���@W�p�t4P�6�����gsd�y�y2��� ��( �L{��G"9icG1������ﰱa��*+jVIQ4M��lW�]�U��P�齿�;繉f/���ꮪ@y���c��/������J�2f��pbz�ZI�p�;������!���58�q�%h��B���)g���)v�D�w��)�H�8��,�h��\< Y�k�顐f�)�F�P��b2*�է������{?��Qi���81s¨5�h�W����p��U����b�!�>H�K"��ub�C6\�ڤ�-�A�[����ǿDf���=3t^��f��+&f�ux��i�����(Ɇ�e3���z�X�vѾ(<� �%+�9J�������s�Gd��-y>ύ�&+�^;�߾��K2��o��ɉ�?\��;Q�7040�_�G���͇�x�y �%��,��:�0��r��$�P��65��͆T6�=Ly4�_|�0��Xs|�Qή�ݻ�M+,r�C���*�)���w��7�^����`T����ߜC���O�����py\��D����{�auxѶpG�	u��A~2/˨��W|jn���w�l޿���;h���v�l�!�N�=8{p������z9���ڭ�x�����h?"A^`,�������B��U�)&�>��zk��p��-(vJ�:�/����׿�������Ϟ����<��A�FMb�P/={N�?��9Ju,:=�c��%E�� u����=d�4
y�VoH��PEA,>���qBaЊ��5��q��B�f�	�B��M"�&\�C�7�ǃ���|�"m;>���t�h��xf/��?��ۨ�r����!�W����:'��_�XY������]�6��^��f�"�3'�T,���_#�� 31����xܘ�ǧ7�A��߿�����ܾ���e+I�ZEh�
f��8=?-4�x��r`7i���C<��@&�G��|>]�_{�<��:~���b�H��F!���t/=7�>x�?�gΝ�[o���V���-[���ˉ�œDu,?M��ҪL��'d��`��#�鰼f�zK�i�&[I�����n]�ez�lPF�Ɛׅjb�{UzS�/�I<1�ܘ����'x�[����6��ߜGf?���^{i�\?��Aq���W��{�q��.�zU����P(��a�Z���݁�D��5��������<�r*����g�`x��[��?�w0��e;�z��F���%�����p��R^]C�I�g�46����Tq��`8�7�6��\��[w
&�Q�e��m|��o
e�o��D�G�z��o��Wp�=p�������~G��_��ly�5wT�6J.�����E*�B!��3����FX,+~8\�������'OcQ:PZG$7� �����'�䁙��?�I�r��W6lF4�)l�[Ƿ�vk�x�7oca�����Qȵ��B8>�'I<�<��i�.SY@��$MxF������D���\��OQO��j��i��������~V�A�Dtp ���B^��~� "f>2����|�rG$�uTZvSN׮��I��X^^�n���EE�X�ԋc������>�y}�0�_�G6����,j*K�������w�������'P��n���1h]��h7Z(�(��r(@o���F�i6z�1��x.���sVH��zaV3)�������Aַ�2r����<��N]d��alm���4v��q���g/�!����-!]�cqdJ�r(�RZ�8h27������V�`vl�6��/�W��'��{��Z2�밙wG�>��'aF��@1�z�kYX9�x��&1w�;^||��X����1��rN�:5��A/��x��QI�m����DB�0>�����,Ν9+�o�D!���N����[ݥ����"(�jE�(�l�[͖����~b�Ά����[��k��E��jӅ)׃w��!z�@�w��ǫ�5�����z�V�&:tsSO�3g&���ll�{��� ���uw/'nz)}�vX�#�����
3h $����mY��������������]Hz�JMr��d;$��e������R޺�P�PnTN/���)��f��l�.:�h$�b�$�m�!G|n�Y���h7o.!���js�ER���ܼ�摚en�Sn��/*׶DQK��+&����VU����i$WP��9����|�~�4%k���Q�E"��fx���B�
�73��~�3'g���Z@!�£G+�wo	�i�z��H�R|A��µِ�764���m5d�391�Z��ͥ'8\YFv���U����U��R% �'�7�<�#�p�`�]hq�h�@�x�Q�S���
�K��������5L�����
�}�%^ݎ����©�����pݯ nI
���7��_���o������:�ѥ����vyQ�d��o��u�#>�׿��*c��B	iM|o�ۅ�f�+�JY�3��4�A�4:��
���(�)��^�ڱ�0�As�b6��/7�����&�@�&�e��-)�iL?uz!�*4'�"�(N,LH�|�5���ֶ������ �r`�͠���NcC	Nl>����
�G��[ރ��6�V�9�"B�3 s�	۰9��kA� ͨ�D���brn���h��w�p��2j�&�G���˳(g�x�DdrK�h6k����W�/��7�wB��O����a
��~ ]����QeptϿ�<��6��YB�9<�$t��*�fvo0��l �"���.6�<Zf�X�9�!7ii�Ւ\�/7����֝R���![�k����nC�Q��㓜���:���;;��� >|��8<<���g��DbY�;pwy�n�m��c��d0z��¨�e�|rf�z�^����q����`P�o6����p�B"�?.Q:,L;��'b8ra�v��V�����n�	8� [�8�Fs:��Q/WDn{��,F.C<^/�Wￏ@$�7��<B�[������G�x�ճ���d��w?��o����
~��Uܻ�_xH�I-J�5`����aok�LڔqQ��!���c�L�Z�`cSH����w��j�@ՠOI�{��˼�`��g���BE��^��-�0^z�A��C����:B^��W�uhB������%�������������n%�9#htmMa�kR2;⩱Y;�L������Cv{�Q���o��1;;���]��Ep�$Zz?b���@��*!����a��.�*��'k�;�c/U@2_@�῍�������kx�ٳX�!u��^*����e3���_��9�V\��P�N����
�g�Xy��x4�j    IDAT����W��,"}:��HI��FYbǆF�E<! v8t�OIEl�X��}�|�vQ�'�i�|����I��26ņj�.�E޷�F�K��fP�ާ\Wn����Ú�p;4T�I4�I���.��å1MÕ+O�w�ĉ������?����<�>4:T�u�k�if��2�m6�;1�B�h����c��Mx�V�>uB@b<���>�zmg}#���X��o �t[�<*����{��o��Tfr�K%\��,qZ�zI<��+(Y���o�y������ZՊL�զ`tb_J`g������=!���k��Sp�!�C��n˽ 0@Ͽr��	�NF��Q���n��
�js�0ii���BK���A1_PF��F�ސ�[F��XB8��t�B96e���p@�5)榿����D�z�a0k'���,�jEi"���0�C�V�
����_?�j.���q���� ~�����=�󯾅��ŵ����f�[bO���f�U���6�6#�U� ���{C��r�yC���îw`m�pr:�3SN���2�$ַ��{�l�"���y��:P5ܒ�ڮd���sSPu�E������qra�^T�����y��0���>��p��&����p����d
�?���RŇ\������-�L��$ҩ��<j�x[1��144 M'���Y�v�F�6�jRK�:��r�#
����&�CB� �:�p��t��.?����p��}8=�-f��~{逨�/0�[do�Xm	��Y�K3h�4����d6��]��BZpE�ZD��)�Bai��"�l�nv+�g��x\�Z��D9�2�L��L�(l�V�h�6�O����/}��	�^XT�[��3	��GKH��܅�B�us��>T���g����|�k7VP�v�9	�bq���KH��ȤR2����f��Ej=<8�H$,��QmS#��Y�=�藛��y�o���3h39��d��Q�,ɡ�>�9����\���^��ѡa���*]X5�bG�*MF����9�娞'�R-u$�"�O��ӨV-p9B��ьJ �􀹬C�AS���Dl  fkN���d���C���8�0���'���4�Q]+�-�+�x���}ׯ�ɑA���Eܻ���?�N�_�+��O�>���)<Z�ǽG[�h.�f���}���y�u��'X��!& �7.���d2,�)���fQy�p��hr5k���s֋��6s�+t�5���cf{XTN���Q�+ϟ����O>�DB0���0=w�lu��O���t
�D�k��b��M�N�'أc#hR޵����X�5���u��bH�=F�~�ѓ�T��J�sJ�����D@��/.'T�>�jI�J�j`0����g���*�~��"**��"����`}��\��X8�W^y~�?����w��<�j�MS��k��oy>?��u�j|w�cZc(B���F�PE9�G1�F������vm�x�P~�n��VE�v��=��q3�;�h���=ڡ�
6�l)A���ÍZ��v�.^��^:	�2����F���?�.�n�y����*N\�|�+ �k�KE#.2Q�_j@�����=���dߒf�q�(�ܰ�,b��N�^39�9���C��Eħ`2E"�C���Dm����� T�'��dWd��Sx��Q��gWp��x�q�]����������Zu|���� �������w��cD�C�9��:J#��o��tłO�ߑ�!�&�W�P��P�NYG�D�)RYՆIB��p�����4�4�:�Uא&�l�7BfS��f���ܗ��\�"m��rOSX)��bI�B�x�9��&~����A��_|G���?����!>8�����mB2��eH��&�B��$ںM,L�J3�t�c�,����-Թ4*f�;���3p�@�&�����W�֩���a�z!
�bC���ǫ˸s�!�.sUt5��apvO������m����8����:��/ށ��óϝC�j���:��:T��Zu��p�� �e�y���
E�J��&�u�}3���R��b6�|:)�C���d��/�9a����^�Bu� ]���A̝>���B�Ր��z�:$VR6C�|�l{�&�P���܉���T�ڜA7�RZ�m`z����"��$���ӧx�ͯanޏ���gWP�2F6�r�����^����d/�NOAi7p���Q:X�X��G��h��x�OD(�M���E���p�Z<��D�q�=VT�������]��A��g �� �>n�s���p��!���^����w����P,��G�zU����V��'�
��^D�lÇ~���5����}�s��,�@8ff��X�t�v�RU>w�wQ)WQ�`��$�1�rj� 21��`C��P�vd�Y�Nv�K������f�0��F�����oV+�	�"9�����S�����a�s���Ed�6���-����("/��NQ��"�����ǋѾ0�k�s݄�gÙ�&QVe3��gWn��:���3p����t�h����^:��ςR�"tߕ�M<��B�RE��I�lw(P5]2]+��(�O��Qx\<~��Ǘn ї���C��T,?:�����O8:2�s��vYq�nW>�}�q\|n�\K��8:�"�ƚG��ckk;�{"��8]��w�&U���Q�C���FB������Z=�=B����Ti�d�oo6����j/��l�L�I'$����N�k3���g��������H������X�+AqFPo�kXe�B�8��F�K���͠E�JlCd�"N\��	B�����D���8;�ϡ�Xhb� ���-l��Hٮ��ۏ��A�a��F���Q���L?A;*���Ȕ�B������F5�Q���u��x���D:�E| �G�����è�,�g�b�{��6�H'�����$M5���dC��;��{�ĉs���"×;��+4����&�w�1��M�S�Y�r��M��Z^0>������aN8��Cp����ӻHl2(���f������4�M̰,����������4���RIP�G��E�8%�_��0����b �c�_�}��V�k9a6��:RGd�y>7Z8�~�9��
z)w�n�QD�����^���ʥ���81;��q����׎���&����E��(��G�p�*GO$e+$�y�o��n��ڢ�b��"�n/F&'0П���5I��i%�Bd��v]'{��q�����^Md�(���c�6}�N�&$��UKczr�l��ރ*���<L�P�� ����F �a�$����n���x#�:�A'^/�V��{X��F2�����N-���|��1nݾ�H<.�ݰ�����P�X��C'�����_{��W���6��gΝ��Qܾ��K[��.ɬ��V��5N�X&s���a�J�G�!^[�&�� ��?���Q���k\:��������$N�͵�J�� �ZmB(����]/�'�͗/�YM�g�����9|�{o���x������`?���\�U�������F��,H���$�ssi	��K�n>��^����g�u�D�a$�^Bdh� ���5x���t[1���熡5д����cu=�t��j���1o�����7�;����jS������&p��4._^����p��"Μ����>���d2�˅g/�`x,��r���]�4/�:��:��2B��,��,
�,�e�Y�	��A�VT3i	�w��&"Q�]N�#&�'zD�/�U�̔����r3HL��XI#�Ǵ&�2媔q4jY���<N/$���)�b}I��_|�����������~���ܶ�ҋHx����3H�#8�#����?��{��E��mt�l$��ق�cd��!48%JvF�%�h �#�bb0���J�b�,75�k�m���� ���t[�;X^ZC�@*U���������XY���?��l��|�%�-�cuk�]}��Q��|�'iA���w�peoX�e66_@�%u�n絬劰0���b�bN��G��74��@�h��b��%��ǛA��)�G���ph���6�T�w�f�it�-d�D��*�pjfo�F�X���N5�����t����u�翾,&G��Q��I�xHxcA�mK�4�%,]���7q�z���]�L��+���9���<}���Щ�0ְ0�@ȉ����DP���M�~���|9�{BE��Ѩ�����-瑯�EW�ՠЫ`SE�@�f�!�MC���N�j�|4��?dU���Q���A0��?st$���F^�N�)A�5�F~�̭�k���C>���ɗ_F0�f�TQ`c��b-�S���i��`�������9/�u���W��3˓��n��t[E8T3�^�bxtã�2�|�v ���X��kr�����f���:=1k��k��jj��&>��_#1���S'����A�Dt�,j�������䖱��K����-�4�\"VF�V��Q[[G8�I�������i��V-���fԉ��2��m!�Y��l� ���i�	�!�^>R)+,J�-�t�둖+dF�$9E.O�z6�����`M�%e�r	iN�s9�K�#a�.̡���v%�Gl���*X~�ώ�R�Ոp'�.@�G����D�
�^U2��2��D*����.t5/�z�{�L�'�^���l6�>�V��3��|/��yiU݉f��O�^g���L���V��F�y�fqq!���F�A�Mllo���
��*-�])>yY�!x1���`zjX�2)�>����cC����F%K���f=$�ԋL����U�qٺ�Q��{��aC,�@����ڦ�#�����5����4k5��!ux�|>�����LNOI���25���C��-?�Sle\*ĶȇU��$��˒�=}Q�0����[����Bn+ba] J+�O1=1�s/�ѱ��q�i@s�M��A�!�Mf/��:l&(��d���Vq�T�(�?B3�0�xm_z0$ٸ����]$*"~�5�Мvt���(�����
b�̶`�D��)�hW�sx�����N��|�n�R�O��ز�'���Z�j��ZN��B1'C�3�L�
K�#�Z�|�LV@t<C�|O��6�r$w��"}_�b|�N�:�p$�j�DgSQ!lnܿ��~ݓ����o����7}�&i��8P*�y�D[��dTx>�������ZǇv״uȗ`3(9�T�uЮ7e3�e3����;?��݁�R��j�G_�Љ���!�����ۡ��S'85���&�[�m�n>�,D�헨�Y;ZTRd����0=����kWQ,W11Տ�A6w�x�xS���#Cܾz��U���}����B�����[(������%���wS�DpX���?MW`4�]�!��;O�dX3:5���Y!K�������?��h_lq����8� ��Ͼ�Q�'���|�m��<��B��ţ�=l����y�\��˛A �O��T�v��p� ���s�"�!dw!�J�g&��>��J-�%S��9J��_� 
�o���Vw�<F��A��C ��H?.>;���2~����կ����+��c}kGt�fqr������S�ڄC�e��'V`,h�.�rr0W�9�z�!���r��r�����I(1��"%I�j)B��҅���l"L�(�\s�v�BOD��""7%�N���Ƌ�11�D�`��>.��g�"W�㵯|��%���U讐��'�ꋮM���3u;U	\�G�Q���2֖�Y #�H0�6��Sh��A-��PboD�N��a��O��R�hT;x��+�k�V*H�(�)1q��y��}�5$E���ǅ�a�?5��q���ί?
����04����;X_�����ċ�O!����}v^�o�qJp�_^G�j��`���z��{�J��P4x<()�<�%޸L*�J*%򦁱q���N��@t~ �zLJJ��8�5�Ԭ�L;��#-��P6�M��4�<{~S�
-ocwo��pbqo����o?�'Џ6����
���*(8������ ��ܕh���t	i�$�����;���$l^�Ik�8?�g� �è6������+H&�8�VвjP�~(v�V;TG �b�n/<���!\��Íw01����0��~m	��%�F�����1�����p��L�Laf6�d���O��cS�H�J�ԀSw�V�p� ��{5PٔXhVvEE!�A��C�R]E��(F���
�P�4���5�!�5=��q3hN���l��/��L��/"O{'��QA��,�<���i�4�ܺu�|Ϝ����(޽������ѱðy�X�&�D!c���f������"�_��˟�h�Z��6C"a`�":��yX=qx�������Y��(�����D�.L��adȇ�~d�6,�&Q�4�_���҆�U����)��(��Ţ�!�e��k��u!xZXl�&yg|e�E?nlI-m�+2�f�+	��$Y�QHge�F��zb�)���|qk`H�f�6������6b3���'�8,H���"�ΦO�S�_���_�󺈗B���F>'��05ޏ��>�]���{����5�J�z�72�L��z�
��'�/^n)�f��A4j���hd��p֥���O��ں��sh�D�O���&��,�jZ��D̏ٙQ��Hp���]l�p��D:_��Va��O�CaNU��\����+�Mt���GS��g�,�V�ue#],�ѵ4a�HNT�k���5���'���N��ZG{�gr�;����{D�&���NpJC������pD�Xx�#C��5yVo���fP P���X�v�{|���N�P��bfď7_C�o��8�O3��Mb?U��n	�3�.�-�.u������f�2ѰӍ�X��DK�<���8c��8�B�z�6���,S��������Rn�C����� �}p��1m�j�̓.6��:D�a`�l�#�L	5��͍v�;=�h�n��t���H�X�X�=�Jz�M/$�GM�8��ޫ��Yt:0�H�`���iD�̙�|>��o�m�$�->���5��I��c�_XD��V݆.�!B��mS�{��E�����qn.�����U��*S�H�=l�������K���u#�M	���	f
W[��:�3�FY(�6��$����AU�e�!4{�l�P���l\�&��lݒ�rH���K��"�`�c�j�v7V�H��V��^�(�cts���H6� ���J�6��b[�.��RQ����r�i�6�D^�-s������M!	�dɆ��s�#m���"E�6�|'��sϚ��<��{�׉�G@\�-��f^�����Pt��4}n���+hT��5�#����Z��E<�0��5(΄�ﵹY-�Uf�̜nJ�gG_3X3�A���]����2x������D���� ��|&ͼIOe�\�lͲ�V9��;*{Ld�̎Tl��*�}P�a}-#g�ۣC�;�s+d6u�XS�?*��T��hX@i�6K%R�R+�������A*'
H��	M���33��y���@�L������]��m�/.bqqQ�ѵ�y�x�Vcq���׆l:�6i��w�P,��
�%����B����11G�
<~�D�X�as�q/��߻-�.� 4-���%\��%p���
����c�?},�r��D��r���$��r>����	9��[�}62�C��[_?�͍n�y�B�,S�@ ���f�����������ų'�[�w�ƣǛp����\��h�K�<��E�D�w=��mB��Z���EtdL��~Bk�@!Ma�b⦙��ۏ�f�������    IDAT6e2f���ň�3��� �4��=3��~�Ho�^F�Q��3���u��m��֞E���6��L�:�
T�������O�`ei6��u��E�Hh��p'0��B3p��I��#r૯� ��
xk{�G�8̦�����Q�VK��A��D�NZ���n`b�'O�����'�ބ���`jG���T~9��b�
u$�2�_E�Y6C�W	}��b��69Lx���e�Ie���K�P�KL�E��R."�J��L�e�adj��QtU�����ה� n L̺H6�_�b69t�Z��߀a�]�e�JTu1����������_x�4��O>;��N��(��c3�^�-4Bw�mct4�f��۸�=���[��E�A���E�g���?�Bb�9\x�$Μ����5p��֗�P.[�-ա��fΘ��eqªLV#���D"�x<���2�7�$�ٞ[��(��!������*����1�R�S�2������;�B�^mC#�6�9�P���t á;a1l�r�Y��F$�J�\ȡ�*��OL����d��ޛ_l)��y?�$H#�{ 2�[��d�/��F^'q�Ex5+
�]X�y��3�*��nW0=;�7���v���B��A��F�����m��L"t�03�v)'4��בZ��N�^�r	]̓����as��	��D4�����ͺ��a��G�bv8�Ɂ���h$��H6��~��t��4�v�z-<��fB�P����,P*��鋶�P$�^w�II5鼝&T;���܇DxG����R6��Kq�Z���ͬG~������d�nW�AG����C����i�9ƙ����l2��@D@?l���M���j�勍!�C�d	ab��TT]daC��t���k:4�RY>����I��}8J�dS���o�&�)��-�řɉ/��fv��:.�����Ν?���S�5/��R������E��z ��"���ln��x4���~L�1��	{G+�����NN20�ހ����@��}�
��/��v��
I�D�;�Y��f�p�5�^,�&��P.#�� aa����E+�R����])�|.B.����ޑ\(� ����ud�)ln��{xpn��=�ύl��j�xz�o���S��5�i��bka�����4�n�[���ih���>�s8D �'����^B��#�?�B�)�]Z*��X�FK��B&b�����~p��Ɖ�	y6�=�����x��cpj�x��+4j)6��r%-T`��A<��p܇��C�q��*�U�ߛy��,�j0(����x>����>�`7�"e�ճh������7�nŧ�a4����9�����B����ysU��lp N�
Z35[�B�����$��VQ��1>1�S����[`p�;~N6�v��rCx�!��G�~-�>����Pԍ�'|y������~���Gk[��o)A�����_cFB7���ώ��Z���{o�l�z��*�j����� ���!Kp��ƌ�"#/��
P/Ʀ�kw�_�1��w����ZKI]��s���u6Je������ݡ����;	�2���fCj,�����dq�������ʵ
V��e�Bp�z.3��׾K&YŌ$08(���`�+��
���Wސp���O�I��y�{ǒ_�Y�*���Ɖ[D��:Ej3�(���C��0��=���8��gU����nw�����0Q��kr9"~���j����n���:0���<���������^�*��9:�yt�=v�]ny/��n9�i�`�����%�xm�[sBry���Yb[�x�(W
hw����w�<kn��A��� �ы'�d��>]�������o0Ű������5��|e,�g�͆J�"v���5ܻu[��^|	��%�Yb8z^�c�ŗ���!d�%D�{��Tihj!�^��ׁn�@�:���B��V�
�/�l����3���v� �1 x\!y��#`q~c�^DwW�������R�<r���+	�:�U� �ɡ/@<N����Q���y��װ�W@��0L�2|Y����NTd�K�(�J��u�V�-kZ>�� �>����$���q ���+�b� �[�+�^�gf�ED:Bc.��z[0$��Ň��L�
����A�:������ �G<~��<D�j��>�~�}>��[�X�|�S�O�����m�T`�F��%V6n-&>�c�h���� j�vVV��t	���d6�����\�<|C^|�9�.K�Q�!��.�c6=@(�;H�^	G�$Z�s�?*��`']E�e��Ⴕ^r�+�PK�Ҕ	I�R��ۢ���*��u�I������Z,����t��FЊ�"�wwkV�#`\�
7���%|�	��ւ~���-��̜>��)�x�zr_�~�M��S�Es����)͕kH�������Y���@��!}Nؑ��hB&j�e�H�i>T�izP���0 Yd�Z��~|l.E�ӻ7�����o<@��4�:v��FN#>w��(��>)�Ӆ#x�:����8���8ൻѨk"?9*䰾�B*WC���Pա۽\�	R���M�Kt@���n�!XB4҇f��CL��6��e�>��rmЪA1���H��pin�}a��ll�������	*�P�z��f��n#M���\V>�?��G1���_K3�#��"�'�Ȇ�l�!|�!�.1J��}��D�6�u�b>�k��ɸ#�~D�A�F��=��ak/�\���'����gn{a�{��X���Q*��DK\Av�>����|V�H������͠;<$�),|-�pI�8�q4���"[��J�>Ն�߇r����9؂a�wk	^6�VjŊ`�Y�tm�Ț�	FxO �9�1쪊R!#C%b��v�@DH���^jU*Qg$K׊h_֮�էk(���� ���b��`�<�iJx5	z���m��c�?��'`�C�ͭ�r�ڑ�9� I�aCH�/�q3�kK9�<dE�d�%�Q��%�V15��,��'������F|�G
���W/�0��O"���cu��ب�E�d�;�-�����It�U\��!���*.������	��p��FK���"�JH k��Q��!4m@�Q���Р?��9��M�y]"q��:�>�>Z�X_/#U0�0\|�M8<~�6;���A�VE1�B$�MX��@�E~�[��@��ۘJI�m&܃�'z��@	s���f�!)AV}1!�juy�I��m�]k1��*�kW��������181�j��|�r�c��/Yx_��aD�h-zrC)N9�5���f��p���N��'���Ǘ1>4&s؏������G�����4g��٠f��"+���^�艱A������-��_�Ui`fzT,)^6̓�nn�i�����|}}���CT,�l+Yt�����m�t�z�F01> ����6JM;5tm�\mH�e��F�`��݂j%�퀡�Z�q�:��N��# �?		�`09=��`E��yv�B��*�{�����&�3��^��ml<^�'��o�
g�ы�2%��@6��Z�ms��]C6������˼զ٘S���Y���H��BzOb[�(%�1A�o�g�t7��dV{�*cF(��˼3�����͠��+>�f/`��Et���B}��r��.�:FA�Gv�j
U���J�l~�V��Qˎd�
����lg3�J����N��Q�㕚�ҤQ��b�v�YG.�6����6U	��W���Q:���-�N�����b`2%��|]�&ՖuN�Q��;�P��p�X<9/��cb����X.���?;���P�3��S=�a9�����4jE��6^ya�j�߅K�I��x14>"�KW�#W�e��ˊe�̍:�̖�ӎe�l���_�Fn����Q��������pFⰸ�����u@��`k���2��k�,F���p#���v���V���+Uܸ��@L�Z5k�ì�U����S�ux.��&A��
�nn�%�J;r6̘;n���l�F�x3~J�F/B����F�!1,�7x�}��g�]Y���<^{��?��?�^_l{���f�g4餼o�Ql��RB<���X?bAZ�Z0�6I'Ȥ���ϋ�@wxQn�w d�o��.׷��8:]'�Z n�V결�
891����ɦ�Po�q�n`k7�t��t��\���ۇz�0���Clv�zE��5��y�����\��E�P�Λ�66]n�R��j�x?����j����U���N�i(:�B��]\oom��jcӓ�/V�}�K�kA~���9�w1;s�.�>��0,��i�ը����a�b0��p�.o���&��y�K-�+T�:���L;|���D�l"$��fI&"�#�g��_����H��E7�ku�fN��g�����O��@b�.o@��f�*�5\-����T��06��mw���rG�q��˪�b-*:�X��YzDO6��L�g����bĀ�F��TN��Þ23D����I~���5	���"sQ,6(U$u�|2�UY���������K�4q���C�{�E��d�Ȑf�t�J� 2M�o3��ҺL3U�.�un�k�4�A�|���߂JM����W�{PB�͜�jm�|p
C����FL�-�����`��U<��!��ѥܷŘEK��y.� �ۏ����k�O%g��!ҹܪaݎ�A�gs���Pn2���[����iT=��i���{�xd�#�B��-D���,0+�N��Y�}��ʦ �������lQ���z�E�G�"��h�@�Af�8=�4�hyZ�jv��T���KaΉ���6��۰|8��Ey(P
�&B�}m��dp�,|���Ќ��]�-��:t,��T4Х��R�p̉����[��Ć��R]Xz|����3@	Aq���"ٴ+����Q�uca����y�Z�㛟�ΥwP���
�A��c�!6s��Yh�~�#�p��0�5��64�$���W�5y6�<nXy�Jen�
EX)����� 20[W���͂��5�
�ү������h~!�5��kB��D��s@�.��]���{����E��ФLE	��x�R�P�O�5p�v]Q�27Z��Ф\���ӕ'�L�b���.��x6a�����a�Ҽ�x�{L�c>p{�J�X���w�E��|�+�����{�3��e�wp�B��4���o���4>�|}S�Q�V�I�W�LU���d3x�ӏa�@���{􅂸x�,~�ޯт����h(Q(�a�ϝ*`�SC�Q��a��E7$��e>���<:�2���4=g $�uz����$3Z�+>�q�pL��N]��3��-J�j��T�H$�<��q{|�Pkp�-���GOeH
F̢�Ͱ�{Ly(�"��	����f��f}c�l�Ϝ���8��(V�Q�f^�ـp���x#aN�9?�=?�<�;��K��|�6��߽�ͧ۸}�R{I�ZTd���_�
5�|�s@�K��@�H�����zS6�q_ ��C�%�����o^BWi���YyV�dӽ�r��Vcs�Y�+�����)�/}۩�t���#��v��N�,��F�"���_��D��CuŐ�5`Uu�Q�����F #Ђ�ֆ��E�i5���̩���;6�Bl��@#��R_/|^�ܷ7o߃/��!�P��&�����^)�|���b>�'���L<}�f���i���r3q,=�K圥��	6l��l@���X:-d~��yd����_"
Ȧyh`�X�����6�����$��@��<���ݳc�Pu\��%~�=�ݬd��A�X@�Cs`�Ah�0��#и�i�N���[�SU�<�9�H�٩}h���4��nh����8��j��p�f��m¨��p���m�]��ؔ��3)��v]1nϋ�Ԫ���vA�:���ÔԱTB�>��H��@��.a:sPY/і����������k��y �Z��<n������	�R�r3���Y�v�Vo�<�B���n�U+���04:���9�j�so�ӄ��h���"%�˔���Xk-����Ӟg�
f��:�R�DF1<���8�.'?<~�v�_s>�]T�Uhv^���
��z����������:��Z�}۬v4����Rf�m�S�&r�q�U��ծ��#
����z��D�am�x�)��e�Z1&��\�Ԛ�W��䖗6{>s�6�q��e�-���2�<��3?���m��shJY��N�@�Zn����2��Rp�S�����
@���#�T���%$2�M�q��raFK8`9n��Q(J ����	O�AoI[&v�C���� z�A�����C,=�A���f����rx,�T��IEb�H}L�P�J��7����~���1�SB��vɣ����!)8^JH���P�i<(����݁�talj��#(�k�O��1�Nr�w��,�}u������ H�	4�jn�N7�w���w���M��E��#i4F��(� h��h ��������̻��j�]�
	4�2��y�󸑐M�W��n�p5a*A��"��$(q�2S�%k���̍���A��^�����`}c�no���:�m�=9�+����f�Iۗ� 011b7��7��x�����v3�Ӽ�F�_�Rc>q��i(��ȑ� �zQï5�f��W��j�D���H�#H���M@	��7?���GhJA����ÿI��ii�H�cǦ�k�&��>�J�!� 7��`8��!���=�H(�Ã=�+e8����E|q��6��ӑ�9)f����x"6<@���ϝ�>����[)���m�'�l�4B6�����`7����Y6,�5���8����X�7���rx#�Ncx$��7�q��,�=9��c7�br{�a!4�岤�Zn}��>}�͛�Y2{� d�c�0|�I�½H���@���@�TG�c�=�Ы.�JӒ�I"�``d�� ��ź��}^n�}4�6L�-�����Cp[MN�M�5���zpXfPwP�-ʅ�� -#Q)\�B2�D�ya~oO �0�\vn��B���*E�Ѐ�,���!����'����o�Yg���n�d�H)��q�M� �&>,̴�?��#��85;�g���O�펆h"&��3� ՗���7���{"�U\Q��=K|�N�y��S��5���C\y�5�W�²����܀� 5s��i��9�3Ò�J�?�AK�'N��b1�[6�nh-1 �8^�Lo~r����	Ra�� ��N[E4@�o���E4����Vږz�8����Ö޾v��Q�T����r��#��W$/�%^h<���f�L��M:?y�(��͖(,��OO`dnR"&xV��F��E��Q3x��M͠d���Y
�^{;����;'[Ln�n_C�Z�!�/��3��U\��:�,��<�UK��K��9j����wѩl�?�������${�,~���hY-<U��)���9�B��q� f���%Vu�E���k�s�z�]�K���[���'���CL�+A�����OH��|�p\�LLP.�����u��h ���S�&�ߺ-J��/$aʞ�%�{��-�m�����Xy�R�됭?sP-����-�lnbtn����(6j�g� 9�Mȏ~̟��=�J�aI�`������p�I�ˋw�����ڀ���o��X�s�������Mf�/���������v��l8���Zkx����+B�vp�،�_N_�/߄���=���I�=F�wah5���:�Ѡ�M����y�h�7��P�ʳ����ZD4=�N�#��./7J�v[���Vqp�D��!�7��C���n�*	Qeć[6حf�`L�ن�`�H�ˏ>�/�R#PWmË�B�i{�u�I䦢����2��
f�prZT_�{>�%�u� ��P8 �    IDAT=���[D@�4d�b��3m�	K���_?�x����x_d��-
����^@$���\�I8���.��%�	����sc�p�5|��+����D�nIK�$�7w��G`��2Z"; �����`�ߍx�	���b!�����`m�����Z˻�]qt\.�Պ,@X�ph�	���F��
�:�7ܑ��G�FM�(�x�0��X8~|N���l�X�#M!�Kð����2뼨xBe�!E�gxG��<;�Y�I�g��rHmt����x������&i���#@����!�G⶯
{�B�٢�����2��Z����'����&
{[��+(WjFc8��� *@տ>�xI�����W�����	�D�7����6������'��Y���ޠ�D{�O`p�,ܩL�T�xNY,�� �[�AnC٤�j��Z.�d�m>>x�!�,z<�U�H�IV�|l�x�[��	�s��j������ᒖ�'�^W~ئ��Zeݬ�p��������s�!�!7��"�Д�a���t}���Q��[��.r����!���~���@_}v_e��d�f7�:�N��sC(���O�N��&�c~xp
�}(u,�[��[�gЍr� ��O�$�Xr>BHL�G�"���-i9����D.��P܏`4�H<�x:�|����:�&2�x(S"���h � 1�mA���L6>Y|X��\�x�)��*7%c�:NuMC�P�,:�*���M��ȩ
Tn-��c!��J��L_/�O�@Vf��Bɂ:�$���C �~.)!"3/�BhA荡5�S�x���1'o�@�|�g�x�G�Ï�?����v�H�ĠKb���TI���_m+�<��I3XX���gcN��n3H�nrC'/ ���+H`N�&� Vzf���݀֩�g�M���wK��Ufd
�V����ɤ�����w����.�A9 I����[N)��s�l)�"(U
px5��З�����dE"Z#�L�v3H��6Z�|���d�-���踻�(��g��{��֥k�f3(�_����ۏ�A��fВ@z[6��LD�!h�\��Ǉ��y��O�FB�=zg��Z��p὏��Tg�G�����0�?�_s�U�~jb��{���#ܹ��4��p@B	]���;}NJ���$�J%(5tq�T���g�)]���>�X�Y	�����g�=`ða��Y:-$dR�����&6[�8
J�J%	/V�OqX�T�pz���B�{�:�ai&��܇�i�	��`��b���qkpt8E$Vپ�����?9������k&���r��b�_k9��O�$	�$�&<���N�`v(�?��P&�}C8("K�ԣO 76��g$��ɻK
v���v�pj�Y8����Ѩ`������먯^'�Xr�,��0ҳg����Ό N��V����^��3�چ}��`��
Z-&�X�\o"�C������4/���F�EXFErI������S�pki���c�ܑ��e2P����eG4t�}}��O!_���oa'_�/�����H�B#iV���?D�G�NR�	(�vY�?�֗��{��0<?���1�� �ł��E��m�\���gY��fP���E���^��2:풀��y�F]�}cG�ݴ����)��1|~�>�u�`Z���@X~�Lx��D�6���}j~C��CoO_��9��믊b���h(I�ӓ�g���E����Ĺ�"�!0&��e�L�aœ�6�Ai#��W�"���Ќ~�V�!�nh��ӏ�{��x��'�v������ܞ�\�t�plA� �+븿�O(&Y�T���,ݗ��Y�.2�S��l�q��ZT|�m��	a{�|��~,�:!9��F���&�v�͎�HG?>��zx��pAJ#%h�ZE��܄�N��������m�n�� ~��;���G]3�;4j[DK��ڭ��HØ�Cc���_a��%��&�$���No W�߅a:���i{��ݫ@W�N�����%\h�-�%vE�7��Ѳ����h�P�N�/�HX]���v'�C�C�>��qٲ.�_Ez`J���1�j��l�1��"�!��E���b'�5�f#c�p9���#F%y�ŤȻTI�:<�U$����X][C�Z���4Ʀ�d���Վ���$X�P��� 7���e�� M���ڔ�F��g�YG�v���><u~�R+�����F���?�<tŅ7?�"x~r%n�j��7�I�L�77��0��;����0�p�`�H�t����kg��0B�� H�m=�?�@����F�p�'كkK��zo�;"*š�p@k�Ѫ�ћ�c~d~K���{u�^��z�l���5�yss�H$bX�j���]T�l�}>?��b�f��!@?!k�.X�Ӷ�g��С�{�������>�}vY�"��w����"z�Lm{}��Տ��fFp�ڭ��A7��C$#^�����0��7H+n�{�!��f	_\ݐf��U��:D�j��w�e3�� ��R�t�@+�i���;���#��!�A1���<H�z]v�4���c_;{�]�BQ�n���t�A ���&�%l��#�:��r_�U�Rf�A��B��"�D�%rܖ�D:���ѡoז���Iu	�����?�~`h��&����|GXK��W�B!���/\����Q_֧Gu�A�~�W�R��1�v���@�C����n,߹�Ra_ 2UE"և���0�߼�ÿ�&�P3�X��D�3e��a�XS�j�m1E���ʉFCd0�]�˴�� ���~���}R�8Y�T�^kJ �Xut؊����D2��6O�k]�{[mH��	��*��œ���j�TdAd����޸�iH�7A�բ���K$,����ّU7�,b�}N�l���/?��s%�E�P.6%��t�%�Ѳ��VGC�m���O�k�k��#ʕC��B���O=���
~���\K�O�R,6&陔HR^�ϧ`|r��!6����x��0+�p6v���jlH=	iO|����9�!�< [��S�x��X���֚*�P�k2��%�qcm�İP#��vtT�&�+���l5%��~�I��h5��L���;J�Ϳj��h$M��ȉ��Alon��/�J凼��?�ܥ�g��ES�!�274,p9�����o}�8�ӧd�V�I3�FI�_¾�S�H&�sy��wir�)�l�t���h`j2�S�r���8�ٖ�$_(��	��o�$^}�2�{�e��,�ٍ�)��U��(�����g���;h��g�� i�J��Ә<�<<�������c��Ӷ���*,:X�q�k	�QW�pdOU�H�����$�0��C�>���T�T����-�+M��s��y`�U��Ihlm�W(#I�9~bt�F����i�25v���C,�-�����i�t�� O�mnm!���Xn �Ϟ�F�K�d�<�V��i3(~�DE^l@�4[Pt�C=���,��ݻ˒iX�UQ(�0�<������o�P7�v��������=8��\��A����=\y�h�݂SQ1<����LO}�H� �`b�p�[�Kx��0~�����],.�� ����2J�jib��ܳ����t�8�ILO�a$G�K]��>��`�h���k�-���5��<rb
�cY^�B��;��ఈ�=1�dڍO�x�K�Wt�L �����5�Z��;bH0�*i�~`��{*J<ei�����c|n�#9�H��V��6F�r���4������������EF���7�
�Y�6ٗ:��ia�����V�|���-���v��Tp3x-���Go�����'���?C_oO>�~��K�7�?�����&ѓ�m;������k8,����yd���{����!���޿�2�jAC>�
 >F�h�k���t`u��E�6�ЗN��NI�x"J����!^'�G�h������PF��a:=�v��JY�89ܰ���������8�@�,��5Y*P�s��${3B�㠔�ko( 4;z�D>��H��wI��]1���*��n�@��7e�yb~3CH��py�r�|zm�\�ŗ芟j����Lu(���AL�K��k���X_�� 07;�f�$͠�µ�{P5/b}�;�h� ܱ��y�������p�K�o�!J���`El�Q<D�TX4���G?��0G,��W�(�d��	@�X�q��.V6�t�8����������;wn�����
��[��v 78��ܸq._:�zW�P�G�	���<5B�X79]���D�^���$�"w�;I�}�4d@x�y�Q<�~H��0����H7��tb�O��6<f��z�8\r�P[���P
_,���u8|1i;:eѶ��5�����f�S�(��!=��E'��'J�E�7�
�8;���A|����؁�`�x�q�Q+b�?��g���m�|�A{�f��D�����:�H�#)�x�>�V��Mʳ}X�F7�6��2Wr���u�-����ߢ�6�el;p��w��^�wۮc�9Gpɫ6۰�����n�;��o��`��(%�6E�h#F�Hr��l��m�����!���V��ZH%���EX��{�H ��-��0P��p��%T�%�R�?�r3H�(�.���-���Oq�5n� ���˙�Y�Ƙ3x�tV��P2"��.��ٱ,�G���بX���*<x�#	ll�psq�Ek�:Z�)2jn�S�4�������K� �t�|T�Q-G�7��ON�XV�?��F�&�ܑi�����ʘ��k����%6��l۔�*
��>����ϝ{�c�6q��ǯKA�~|�!�j�؅�#mr0ρM��Y�@_s�=y,lnn�^��ȭ�?���Q��-ܽ��om��E-�7ЃX| ^wT����Pږa��A��< b�����0y)�*
ɷc�(Is��zh4C["#�%Vii0�~��dp)�J�-�SU�x��I���X���a@;M�A����%����-�,Ł�UH<3mx�u$ؖ[���uT�8{�`@�A�!�L���A�ĉ��O�)�'6�T��>C>Ny��v�4K8{j3�	ܺ����E���á�~��ME��?����h<��|	�P�+�<���t����O���?��;�Z��<s�6w�09}��e�&G0x���%��#h��H�<x��z�n�}N�v8�����9�7�Ku��
J���������K�vG��i�O�̿��>����������b=��>�kyAE�ca1�?���	V�X^߂eҼ�iy0�?�C�\��`~�r*c/��� ���<��I���j�����g��f�!@5��ɐIjL"͠}�8Ln��A�-9�IǤ׆�(�YD,f�{�:�l4���U��� _G0���*M\���	�.(�C8/]�!씐Y���_Qp�Ӌ�u�-4�o�-;��ϑ+w�$��?�`z�p\
0n��a<���>>��bJl%a|_xh�M��r��O���II��B�zK��*�R�C�#��&���ͭ��11�w;��۔l)1�z{��csr��\Z�iz059�v�������2	-$<��['v�%6/�� �Pdr�������&�=�/�A�w6ׇ��-���B�˞A���5���ҡK�rkx��i<q����[��F��prc����x��[�/��X>x|)��r�H��ӡA1��`���������"����D�WV`z��?~��Y����"����Y��'ό��oM��׮�7~	_<�h��R~>�C$�>�����p����?�9�����89��I�R�Huk�\SLQ��֥ܹ{�f�%�>B؄4T���R�熇�up����PW��������ʇ�e��O �p"-�V�*2y9S� ��@�Q��f��1�d�"��gL?�dwq���e��6����g�e�J���#��3�Ã��Ѭ�1ؗFOO�� ��\F�a��d4�/��|E<�,�x�?:O�(�zSB��x�����>\x�)��g��jǅ�P5"����J��7�U�������O@�,�џ�	���@8�`4�m�Y(�g���c'1>5��~�]�@(��� Ο�@�a4e��:��KՖ�_~�@�bC}=x����3OV�"��W�ࠆb���j����vA"H&�NBqs�t�f[���pHŜ<N��#�#nJ�)x)��jX�\���F''d��-}��Xm�y���_���P��r�~Y���V�K�n����6���p�.�e��c)�jZ�gK��d���@o��L�ǔG��D9az�j~]r�o}�Pȁ��I�k%��Caܺ� �:MMc|�b}C�F#䈡�8��H?��n~��K]"m��E�A���v~�q��3��������
�$�0>2��)���9 ��ͼW|P�T�:^y��	&&06���I?�6
�����]�
������g76�R�x`N2�
a��
��QJߕT��|OigpH3��ױc�H$�l����?��3̾�ymI�9��Bx�.�/A'�8H��J��B*BO:)97��Vwq��ڌ��F�F!>r����Y}���U3�fW&J�`W&�t�Az�<�=
��`"�T�9���!��ӏ����wp��M(����������*�͎��'���竸���@2+Ъ3�F`M��foD��1L���j�׶�q�11�C,����\;��4g��VP���?,��"�N��6��Y���i�M=�J��r_���$�	�|oZK/���D(���_���#���>]��T
4�2�>G~�"�]�ⶊ�����i"P�V�:�sh@��=���v��!�H6R�A�
.z)�gp,���2ї~��^�;%�$L�t$�@����f��+�X�Vĩ�Q���xX���h�+�kJgI�����U1�0���|�����CH�IroK���0E:�!k�[K��?,"�at�.�. n�� �G(�X_���VW9�	[D�ȶ��F���$��Ѓ�f�-�*�B���?��V������Ϛ�_��3/�U�ֶ��]fYr0�\Ӏׁr�>��D���KAq���j��庆[7WP�4��F�2�o�g���YDcY�̜��,"����O t���F?�N3oֶF��<�x����a9�v@;��D�K6MSB���FM�������jc��57���(���jΜ<.�;�`c��b^�XB�"�{��
��B��V��0�����I�q[�mi� nnn!_.�L4����+�Q3(n7gО�PkM�;�%���"�FN���I�-Q=��Po�x�z3>���`w��B�&�7��Pj�x�O�d�/;�p=�|�I/�N>�����w��x[w� �vFu��>fM�Δ�������?_b�T/���g��A��:K��RؗK�
�Ę^�VM���.�'sP� ��G��������8�1�B��GA����Y�*u||y�{U��E��{�M1s��)V+*2���As:���Uܽ���G��;�b����}�P��?��� Y��D���{�ࣟ�4]�/%���ّ����[����&�ךA�'c�x�tKc"���G�����a<sn#Cit:>�<��Z���2V���O��^�*��jN�Sw���MO���勸���h���b-�^WJ�<&}��q��18`�p|$��|k�&�u[�g)��g��|jI�~{��.�û��`!���Q*�h�T��cb�;�U\����ͪ\t�$�CaP�&굦��ff&S�G�.bo��'�!��������dH�ZT�A�0ܬ�^��?;��^�\�a�(tߩ�Y�
@��/3�{/bK�5�(�YN	���x�N�
W��jx��󘞊#�C7�������M���Cw���@[�L��P���v���S+�֥�q�����^D�m �	c��]����x��y(�^S9��I�-7+{Ҡ��oM���~���.D)	���i-`�����~{y�+���    IDAT�7����E�x��t�;pu(�������T�@�f(%ϼA�Sq���2��%Aµf�D-6��(\����Q<�bok:ɘNB��h;)EV��
� ���JG<l,8k�
żd��3p�	1�A��Z[�.�D7_�����IQd�H9�E5J�ٌ���#X]�����hue���`(���8<�4J��lR4���>�З�	gK�S�p��l+��p|0������p.��_�:��������gQn��C0�EoO�Z�e��{������?�+t��$����j{�H-��{09�����p�4aЇi�X�y��2ҩ$jM�Y��zPl��nS���]���ʉH$������SZ���%U ����=�z�
��H���l9\st`������t�������B�QÉ�'�ӛ��7JBy�PN&�G�� �Y�}%C|8OŁϭHo��������v�`� �;���T��;4�Xv�;E�� ��l.�a�7+��Ø�Q��K?�s�ݸ�PX�<��j.O �p��wqX���bl�2�#�q���(`j(���4n^-���߂'����D�m.#��o?ԏ��۷��x��&��G*A��*��Z��e
�B��@�#ؖl�XԋP@��<����K"���p$�\��МP-/��A�'�5����8����"�Od��x()5�B����A+c��f-�񢾲B���YM��]x>�]:�#�s�!^sm?T�0T��S��@n�Y�K@!,PBՃ�jh[nx���墠C���lZl�̿�XC�P����?�(:a6���}�L4J����&��Z�{�~��|�`X��~���U\8
�O��һ˸�q�p�W6�n��^�����N����0c�,��)~LF�Lt��n���e0C5���z��D�˃{˻�d"fÕD3�A������!|6xщb��"Q���S]����z�~0o��n����~Y������ͧ�i��D��1K�\�G�t g�6]���Ը�	�_���ix��}.}49��s����f� ��V]ȫ؞���<���N�"�H ��]����8fg��u{Wn܁/����z�`z������p�7K������Hd������s0n���{��/_���~	�T
s�`��ӎ�Q:h�.�����+��Tqy���8ܷ]�*�~mnm �� sCȂ�����-,�Y���S'��e�����9��.�k�k�/��r��Z0L؜ЄUԪ��ʫ��BH'"pz��P��_��֡�s�����d���O"MfF�t����$D���c�?��;�N���ށHrl�'�m����q�򧫸��	YN���b�V=�Kibjz}�(V6��bq��"A/f�����^zR)d�!�kU�^.��p�b������	�0E$_��1l�_��V^D������M9x���WJ���O�֡��n�$�h7V�+�������v��v��9K�N����,o w�'&1;=N���2��ꋟ�ǽ�}��=�p:�J��A���l7��4OH3������fp�L6�=8�:.z��v�Db�O�@2ӏ`(�R� ��(~��>�����K�@�F�`nTJp[U<������/~�6jm?��Me1?����n�d3�Z�����o�s�[�8>?��g�3��S.j�_���eayӉ��WQc�?��l?��W�[j�D�-���L$���%yL����ad��D&-�{�#y���������g���-�sr�(�ΖHx����9	�Ѡ�K/��018Ћ����s�{wy+�h�-D�}P�Cʋ��-�(nSD:�6f&p��7?z�5nw�T���B����g���4�z]d������K�r����h�uz]��U�.<��gq�o����h;�);ulO�����@S4�ǭ!��@����z���C1��Nb~>O�2Q��!>�j�0CUu�W���^C�������;8�+�͠��5�(8����&1���u��n�v�'�ۆ�x6���a���<S5�B�{\6����1��4QJ@<~�-��o�MxMJ��t��Z���=��I��������P�����yC	t�li:��G��{z),��8�p�z	�.��k������#����C+<H/�Gdh�H�԰l�(׶�2r1��}J��/~|�k[h&`t�
�����yLL���]���]	�?(�kU8Z��kH�;r���aDX\�c�a��!�/���v~CQ}=1ds�t�� ���8(5��%�p��j)��M���J���y��FeHH�����V�V0t�m�	��7e�â��/�ۢ��K(���B��3�
��H���r�'y���f}����vZ���U;�|w[;�6:������kK�$��Tc@��$�w� �����a��/�Ay�.�������������������P�HCz`�h���Q��s�=������*�y�m��9�E��A"���`���Y(>'��'o��3�܍Z���	�u��nyV���l�Z�@���&�Lf��Ы��hD��D?bQ���~��Q(6Pk��)ӭ :?�����/���6�l�}��)II���ͦ�+7�Ğ����p�=�`�?� �P���b3(�D���ʦD���I����_I�hM�X �Fzc���=�l��HW)��Tk�t�����^���U�Z.�	X��V�v~��lJ���@�V�����k#Q0?7�j9/�5_8�Æ���:�~�ΝFvp�HT$��z#�~���Q*x��w��hhN4M�xXrJ�'���Ǳy��nAU�h�T٨�U���Y"cA����MPmꘝ>)�Zm��.45��D<F8F���Ak��T�g�x����M�K�⿖�NJ��o
)Z�����
��VK������������Y8"P>�ݕO�φl�9��;d�DI�ls@Gzs��Y��O�ؠK�w�>,�7(~M��(���U��a	�ᨁ1L�!�̛/㓷~���f�C�PX�ޙ'��=#��;�F����ji=q���	�ܿ}kk�0�D�D�A�C!�%�������~�PT��!���X�X^/mE��R���(a�<9cdl Ѩ"��q
E;�U�9��׻^8�l�Q�kP���k�&X_�y�]�Ɯ�&��-߿Ã٘�9u�Lz� #B����L��t�"�`Zy�_�3�Q	ܜu�΍F���n�K�-<u~c
֗�0���x�K(�jH�d�pGpg� �7�2��f��f�c᭟���)�������Ǒ����<e�)�!$c)��tE�L�p�t��vp��kpBP-�XY�dXmL���sc�y��+�/"�"�� ��%��ahp�f�HO��J%7��-C��n�`ӷK�l��� 4�%y�_��QM�ZAtͬ)�l��A7���c��f���I�66e��d177����}�N�.T������� �a�("ރT�QQŦ��Dsbr<���ă�%y>�䒷Jw�G2��˂��%�}�� t��f0���[�?�DfÏp$#��ry�9<�\��
V��$�cpMJɤ�V��\_
�<�u|��=�[9�Ûɉ�IL���t�j��ۂ�A�Q"��w/�����'óO?���G�|V
|�IւK���Z	W�˚:Nȋ����fCE,����� 'c4�I԰�x-��������h���p{i���M.ģ(�n������.�ͬ|���Qкl �~W^���(�«hr�d2=�FCrH�mW�`�@.1T<��ɛrh�0�P%evz
��>Vo\���8\a6��ڗ�yN	,��'G|CǞ�?>�X�_df�V�����<�k����_A]3�蛄j0�K�V/a0�ŋ/~����'x�]G�'���4F�,X�L��:pXl"�?D,��?���]T*u��%����L���7�}-���G��n0���D7�Z���JDC�0$���_"��Mu��G��4�����B<�F ��U�?��Y��|�9[G;^66��h<��Q�m�-E*'�=ql�@k���X} ����&Ք��<<,���a�K�4{S���+Pv3tu7��Dm���?'�D]}�?��4��`�&��Ȕ���o=�>��_��B�8��8��"��k�!ח�o��X�,���o��K���cr�#)�Jf�k�L�d�@7=X}�/����B$̢��j� %��Q�pX��J�m�`���� zzr`�pw�\.�s��b��'�v���6UEm�\���i� $�ߋh*��]��b�k��P�D�P� <�������Z���w�b�@(��8����� ;>���~S��(U�s�_I�X��F��sf��.�Z���B'����J��W�#�d3x�үp��7Q߹�xЁ��!\�~]��=�g쟆#�E8=�H���M8�C���9<z&�fӍ���������l��G��:���Wqk����84���8fGb�E0��@��Z����Nww�X�ϣ�nc ���Q�� �Qj 5�	x,Qp��䱹[��ϗBGU03>C3$߮ʘ�!�j��-H	ga`�Whq�) �(ҽ��jP9�l�M������mK��2S���C��z��\����T�h��x��y,޺��;�0Л�������kp��-?{���*,�z�@ D�;��US���$�N'>��[�n��Xڅ���08:�o|�9�ŏUu`���(�>��f08>w�%ۀ��5,L���1<݁��=T�B�ˤR�!W+�����
�=�Y�805���`cģ̣���֞��w7d�Y(֡7��a~>�����mi��V�;�x��b_ �M�O�J��������3/�Pn�I��XR��M��U�f��bh|�9���$
�(,�s����t�����tXгi�J���<1�A%ٔy�uX���^�����:������̣g��Zp�\��h��>�n�l�E��i���i�&�>��2�U��_�֮~oĉcs�(�K��G�qG��W���`p���$��˩<�s���~�ILNx��U��f�����T=��O ���?����\�0j�2�~'�)R	�|�Ss��mck�  �P�q-���)R�&��Q���V�����BՀ;�����`�p��w�i:�m]d�Ҏ�lA�����u�*U�P��N�0::b�@Is��#�zGRQ���g�Az��'�D<D>d��{���
!�^��
���?�`������������폢�t�ҵm�:�m�^Ɠy�$0F�hm̍�4ыo�����t�De�8�7$V����1<{�/w8�doV�A�,@�o��L���y�֙�ɡ,�?g���n\_��

`�hV�0��t.��dH�-ry&J���X}�&�b��Fs��M����V?��;L��kw��;ww�F�b��I���/�Q.U��'@5)��׈�Fd�����ζ|���X���o��qs)y�]�������q�(�V5���ʻWX\RvT��av�G	�k��f����H̛�k��c{߁?�+�)&މ�� U�Ġ�dΠDK�w�$M��n�@�I6�'�K���H�3HECPK�I���s��W����6M�l�M$�)d1�O���������\@���SC��4����Mz�c=p�=R%��'�w|V�ݸR�ն4��X�lti�cv����"����c��X���Ee!�E)w�����@nٞ�( %�Vbw����I��C��ٵ;٠J��#䒮��L����)$c
v��awk5֌�n_�h���&ʦ��>.�\P1�
��z��-%�F,5��@"> 4�rq��.\8�[�oJ ����M��B�Y@�y���#��w������k��
�e��J��7�$!�kuӂ���)ae����]�<.��a�ʢ�&e��_1���x�5]ҟ��?B�TA�X���R���� ��J^=xva�˳R+�T/#��"���|��'���	�@�HF SkR�8Ŷ���^�m��A�^�̙*�N���B"�����(y�C/_	A(яZK��Y�P��X����H��-��s�)w�E�� +7n`��-�h{�^�s=�(��1�{��(B��N*5�V��?<�FIŻﾇ̓<Lo�: 7"~�i<{�,�+����@$�Z/����jBo2�: �]=�f�@�DFt�ZC�`a��PF� ����^��b��Df ��#!�T3=i�����ڂp�6�����-�Յ!��r�"2�X2�`�Zhg��C(m���Y<�f��JU�q+u�������n���� �5���f�|�k�ڣQl߯bo{Gp�+k�r��M��n��RM��qsjlh=����AmV%ckana�����������M���U3���9��Sl'a�����l"u�^|�Z/����Ē�4�dn�-Sc����z�[��G/�͌��!��6��[�RL��|����My�8e��V%���� H'�PK��W�0�z	T[&"�4b���[�h[�ŧ�d^$��8�`�N�/�6j���EA*;�l.��+���M�j��~f|�I��b����]"��,���4���yaZR��������M���wp���A��0��
���a*Qɗc�eE�`��e�q��q��}���\���V�ʄ06܏ϯ]���g���
� ��`<�z��X$�jy>��c��89ۇ��E@HT��}V�gw�P��)���J�nෞ{g��t}:���7+�$�!;>_:����;X��3����x�q\~{_|��-WZ-�FGq��	ܸ��.~�'�l�W_��L/.%��s�peny����k~�^��ƣ�7��X����	U�����T�sY���ͥ|~r��C�����>��.6�^+­hh���QT��2��G173���Id����/ރf`:���'>76���ETS�˥||a���Ko�	���Ѥo�ßc0׃�}�;�����%��3@ ���#HPb~`I$Ԧ�D6�w.��XN�6���Z�ºvkwWvP�(�T��؟
��^|��*8sJ�h�`��F�P�_}t7o����<���9��.|r�c���7FJd�@�\x
�;^�Ż���0�U�	ƤX�Jfo�P�'�	��ݢ��$[���4Qm4��L'��&e][.�d��'�E`�)6"]�I�u��2,�JH&;��ԁXȏ��Be�>�����L<��'�ch�Ghw��/�n�ҍ�I���	�2�!1P*�x�S�t�0ޟ��*�fp���f�2x+�˳�8�t��KmlWu�Ϣp�T��Co�`�����\f�}�)�ӡ��#y�/_��;�E{a�
��<���N��h;z�qm��(U�P\~�m��x���g�f�p�mËJ�;�[2�M�z�.^(���7?��!��q!!��I�wP�@��6��}�U�d!+���x��$3TB�G 	�2����v?E��p�(��IB����P���?eod��Is��aW�+Kr��c07���,|!7��x��+�a�u't�Ў��-�!�z��ύ�����荗q��vxnTd�I�(�=�?����0I��1${��T�(�
80�M`r(�$�N����tK5l԰�_Fä2$,�>��O�C-ְ�z��G8�h[dr�[˸u�6&���̓s�����5�E��e��<N����f��ܓ�Z�� )���8���j�?�'[3F�4hgI~�FC��T:�LO)J�='pF�]N��Bd�υ_"�J��%O�����iȈ�U���e�$��<�@��M�att=�8��w���}o��wٱ �u�p�y���x���W~��ŴI�WL!82����qY!��n"�r~��O=6��T�;����"��5�h��8Q?�M|~e�*N��>x=:�R.��C�����0��L엫X+V���	f@    IDAT��ɦS�K���i5�C*&���'5��H<J8���yC���_�������1H-���\eT�H&�L&�����K;���v��ݼ�Pi��O�7�Va�9�ݍ�n:���{,��D��K�qx��E8d��5�K+h�N[A����5�/�w,�)��~�r�Hf&` �` �p�t���?>w���-��s�d�V� ���ӏ���^��.}��p�Wb��-(�*bnz>��Ń��
����8�(,��V5�^��p���96Mll��)=)T�'IL>1��R��rɈb���	JS�G�$�#�fNCCk��QŴ�G�	dQC��I3������'� @�.NĹ�M�Q��r@>�:�yn��|���|�	�^`{�����е*�6����F$݇O�.#_f`mH�حf��_��bH��waf���C�޼)�`��fpW�A۲�a8S�;q��8���N��~�<r��6v�q�h���Hg3��pbj >oo��.._��@�Or!zр&�-f�$�QD#q��jX^�G�n�ɝ� ��L��i���*��N�>��Ԅ�Q���4��������&�TVV���M��@hxC
4�F)q5�H3;;;q�a?��pww�D����ȋER�h ���h��F{��M�����͆(M���D��������!g&���i�VF�(Z�$V�RM�[���cK�L4�@ H�"�#H(�ͻ��laHGАF��r��:52�`�.V*�k���<9Ȟ>q���mt��l�9 %RQx46w:�yo�[5��J8�T��d�*��R�~x�2Qn]}w.���)?d������㔉N��J�����΢0­[�q��]�H�`D�f��F1��;��o"�3���ۛ��0QH#͂W�+Y���N��^��ZÐa�z��0S0){2�5"�?���kX�mH����"�� �ʠ��%9��W�C���Æj;R�bu�n�c�T�w=�}�4j"�b�=U<2���i�b�����I�nd�1��(~M�cv�q���}0���ҙ~,�{ 	�#Ã����ǞƠ����g�������ȷ9Z�.��+@ג��'��Y������KoB�x��B#����U���G�=�@fP��Ѥ���є��C^ɐ����D��Ś�b��V��B�Ƴh����,|��S�i^������%���|����%���W.���N��sO������Տ�{M�K��`|�F�'07���s�д(T~��`0/&ɍ-�pY��� �a�r�pJ���v۶P7��.J�-7ǲ�a%l��C�#����)̮x��ve��t�Ky8��l�a���g�86;��\���zK�+�;sK(V:(������Vq{�(Ϣ������������sw
A�����L_{��䥗�h8�M��'T@0s�� B)/�^AV�MX��SA�D��,au���.�j��^I7�D�R���U�:<�o�0��~�~��W�1���WS���'��מ��ˋx�W����������ro����mx�.zgϞß��g��������i	8Nv/j~Y����S0�6�~�^(a��~Y}�߇H4(%����.$�RN��r!��)M~�9��w?%<��c��i������1��h����x��vkM�)RXj v[�F�{�aU���s:�
���P�^������ �afj�k��Ұ���3ت�X.7�;:���q$�p�L tP����H���`x �H̋������@������$�_�O����_8�^��O�`oo�ݒ�k ���g���l�u�b	�O����.\����n�0�R�]�������^�����Q���K%D�[����(V��3�_�y�槺+�0l��.���.H��00��	�\zK��'�8���I���w��$��M5���a��p�*<�⚍��z�)�a���cjx����v�W����¦e2,)(ݕ�RS�B����qh��~E��Oa�<���jf�Hr�N���Qt�iQ�drY�C���;ْ��1��`" �[U����>�6:jm% �^ޭd�'s��sc�^��ӫ��M��br� ffGp���|�����+_:��k�B���7qrtb'�a�Q^��v���Qʑ5.�}�M.YL��&�Gד�h�dYD%�l�DAJL��V���y$:)-峓�B@Jǥ��kܰ�j�=�M��Kfҧp���bA&��H�HF��z�(����[D��F�T�0Y��/>���?G��Y��k2��?�>x�{p�;���3*R�@8���$�� �;$�/O"�M�"��40���Y�CAD�E>�0��3��ba��[����[��J�v�T�!�II/YVN���P0�f������j"�N��	�"�)#6L�ga����0=	\�� ��vb��B#�ķ�%)=��C��YW�D��[*�^k��#�fS@TZCE�M��~�P~.�O�p�?�l;�2��]�^f�v�F�!^�L��*j�Dh3��� 2)����e��_�7���q�.�ؽ�����w��G�C��Ǡ�{����S�q�Pwo.bsc��%?�514���h/,ۇ��#���,��Ѡ��BS��XZ U���J	;u�l��&�E����� ����إ�n�v���R���5X�&�]��*���`�F���V�~/�����%3H��I�#�	]�����|A^2d��-�AY��N��&I8�C�<!q���	�2��(�ܒI�Z(��6���ġ���l�1�����p�*~���4�C	׭^)eOP�,I�#)fc���`���^0؉��������O3h�A���@O
�OL�'���R,�����A�R�o��O�[1�����T/��ġ�tx���v	C���q��h�-�<9�g�<�����EX�h��#�[W��;��j���2r0�_G�l8uVӐ��p�6A�.�'?<ȘJJ�����cW���qb![�Jb\���|	(����s0H��M%ㆉB#A�OU����Z%T6Vjš#S80�/���k{�p�:<J]v��`��@F�3 Á�-n��-�x��u�}�!3�|h��7�l�Oc������|����7�&F�zq�l���U��/����m�����Ml7��I�Զ19�ų''�69h�\�Π'���ǟ���OnK��ӧq�� �2*�t����uL�LI	r�e����`�ȮJB���R��t��vwE��׈7�,�co#�|6�j�y�p���z��ݣ��D�K��BcW��<�\�}��l�zzW��Z)ۦ{9@����ׄW�Euw���88=-�0�ob��ƫo����6��h�$t�}�]��Q���!�?w����>���}�ͣ�7��|�oހ�0?���q�����kM�ͺH�T�Byg�QC &`6��&V���	%�D�PciX^?j�"R>�N��Y�[	�^���L��B�ͷ����%2�)8{�&
���`AE�f�n�{]\�x��/AUY��i=�Y��A���~�@�)�4au(m4�2|�Z�r$ð�b���Je�(B��J�E���幐g̾2�e����tf��n!=�_&E۲�����9���R�����ޝ9��"v+%L�E�o�K(W)��Cr�d@Y[��x��>7{p�F��*��e̎�������B����~�ӟK Sv���A$�"��7
؊�`Psӣ�u��a�ќTP�%I�>�1Y����E{�jQ��EuwG�{��q��Ž{�� �C���h<��W޸�� �I��٣80G�f�|�,�����_���R]%*���ʺ%ޣb!ʝT�%II��Ro4��I�O��r:(����P��R�C��w%؋=���;Obe��?g�"!s%Nn��)�j���PW�SG'q�hA��:��ݟ���2��,�������W����ഽE�Ƞ�}�
�z��X%��4����KKa��m���b�	��L�@�o�d���eڸ�m����24��}�Jյ��+�v��:+���x�(&�¸v���>����ҹA<��Sȧ�����j����,�L��,��(	8'�Co��ð�;��+C��||���L2)��5�2�R�ϥ�T21��/rE�,��6�օ�j�ӻ`P��%��'�]b��[C|�m�4I3t}���pN���Sg�xɘ�'��19G������6����*��$?�q�m� ������x=b��Z-�.��͟J���`��9��F���F�.�d��А���H���BH�W�+���a�j�V��qaY�X��<�SG�Л�AEK~.�	�u�,�?��Sϙ�==���	����0o��Oo.`u��p�#j�H  �[�O�;�F�w�%�cf��?�|0�l�b�l�a5D>J�%2�@^ד�e���R�3���S����}%`���W�3�� ��1ԟ�'r2�@��c��=,,��������3)��+���ź�$sV�s9Ľ^�����4i=�m0�CH��Q�z���#�$�H����2a�� �c!�FX�`�n{MK[{(�mX��3/dRa�?=���U���v�	��"�����r�r{�K�Ҏp����Vp��'�	�I�{��gJ�`na+[5�,�HE#�8|b��G�!j���6B�B���B"+� %�~R� %���-�+�,�+�����A����o�� �ʽ��UlR�/�����#lKGq>B"�B ��:�\�Wt�JM�k|��ܽ����Le�`�o3���0��|jB� B�(mah(�ٙƆ�d3N_�7x�39icc��q����b�*t<���rPJ9�I��&�����oH���� O0�ۃ��	<QR�&��Ds��{��Ϯ=D8JY{�BH���l6m�-���o��+ۮ��uBm�Tc!)��#� �!��H�"�n��݀���P�t�z�ە�� A!���m��(I'e�z����L������X���o���[������u�kІ�ޝ�#�瑑aTw��x�`���Ơf�1:�E��c��`�^n���2�`�'��B�t�4mK��l���t'�.�`ԝw-|㋧q�` ����A���Jҧ�~����?~;{%<y�4����'���������B�Z�7��_bdr/��,-���s�xCh�LIǣߓϋ���p�v[�Ɇc��|��MO�V:󷻊$�Q�J���
�As���R4�2�3�"w���p �H�W���H��{:fFz�M����u$����M씚"F�����K~�\)*�O	�>�L�K%ĭ�����Dc��ܗ��P�D���`�p@0x��Yn6`�u��q��(�R.W��*V�Ml�oc��M/@��0����O#�Zx��èVd�(�`__y����������[�x��q���_��'��P*�������;��˿��;����}Jf3٬l'yY��Ш�D��.~��j��Wb��e��P [�Е`~��)�uSS�}��-��8�P2&`Е>���앤D�!=�>�mD4#/f��0:܏T�)�&�q��]�T[�;j��x��_��������E���-�9<�N}�}���@��MDI�z��P�{d� �C���O"�7�쵗��&�8��e$�L���?�B"�G<�E���&7��`y��HF�C^�����'�0w�[S�|rs����U7O�aT6���ME00Џ����j&�v*"]T�q���d{],2I���ǭ
�&�ݔ\����p��A��S�lJ�8d|�[(��3,`P��]t[�1Wu�ݿ\�/��]��X����߰���hb|$��f# �cl�P�{8���Sh�
��?@��B�ĥ��![0!3�߇`�ȁ	��\x嗰�k8<�����ӗ��:��?F�2щ�$Gщ�0q�L�!�/Ǭ�:���A>GOoF����̣�T��ha�;:
�'�����[�y��f16���5(,�oz��~r��x�2���҅�?PƆ����"��˸3�5�������@g��,b��!��I�����rA�x$����Ck
L�΄Qz�\^^: �Ś��� ~�O]`�{����#�����u:M�=B�[�M?��� B��Ȫ�G�X({�ݗ.bm����	.�]0�DQ�ݎx�	;���������1;3���X�h ���M;M}c���|����X���[�b�y-��*B1?�a>����l�M~~����u��M��'��iD4 ���!���Tnc��:n?���F}IL��bj"�$6�f��7�V�p��N �	����Zt�rA�+��c\01�n#��"���6t�yŃ�߁�etS&��������qr&�|�u�a�bQ���w2=P�Q�6Csj�h�r1|�� ^>������pqId����l�]dx�_�Xt���bR(2 3�>�𭟊gP�>3�%$1=7s�3g�hj(�T&-`�m�ڎ�l�{ʠУsKb�Qiӱ���ƃGk�T[���P��֚ ������tSB�hy�Yj`�ؐ����&� F�
P:�[��dWo���d�L��"���T _ص�V�b�bT��|F�UN8��xz�ky|2��]K��땚Ȣ��xP
LFR���>A 覩���m �7������^IY�6�Oѓd"%?cLy�,��$������kR�D����ϩ`�(kM�d㪊_=�-7ׂ��.e��P8p��ax	�!d�QXV��"�v��i!�(�Q֮S���g��2h���iפ���(���$w�e9"��B(�ū�XZݔnީ�a�#�x�����,��f�Ľ�5���g%�Z�ay�dj"#JPN���2��<[����|%�WC��p$�xnJƽ����[ 7��s0�ߪ#���,W����i����)�px�Wj���n-��=���Z!-�����4����L�sf�`0�#��	��)X*n@U-�f�N#c��;�O��f���dYfX�
Zz����7O��Uį_}]4��H��"N�{O=w��|p�#c��o��"�{�=1�2����_��t��6����#��9;j(�S6uߎ���-~�k��
>�}	Ҩ_�	|!j�ݤJIēm8�i/����,݂uw`q�cf��"�@2�4u�P��{16�Go΋\&�?�v�.��-����H����I)=�;;��0�:wۋ�
D���?�Pn�� �>������L2�4Z���b�(4��ȈȮ� ���=�l:��6^��1�����A��dM��+���������G?� @��ߋC�#�#�Z[��4��b������nɃ�߾�����׏���fZJ�X�-)��������m�u�÷��y5�����o��l���}Ώ쭼4�Q�L_������d2Zi;��W/c��8���c�/"a��%ܼ}���P�M�N�{g�	ş�W�3HP [;�N(�+801
:�n\~s�^Gc�2�ңƢh m�$Ǝ��@TL�9�����pZ�"g��=��2Yt�Ѝ�	�E,�'��R��`�ķ�y}�8.��:�;�2�Ӈ�q��$�����h4M<��9�̤p��#��KHe�h�6�j�G�0�ڛ7��U��on��
�bQ$cL9UD�ɮ$awn�U�do�����Jʣ����-e��cCN%�&Zjb�8ǿ�~M��(�(p����P/<3���$T)����".~�V�w%���a�hB��a�����������6UǙ#�Щmc��q��7PY��D*�\*����,<z ��Y$
������9��cJ�p_҇s''05֋P�F$�Fk�bo64�����Qly��ɡ^Z@:� ��U5%��ģi����,�Ry�
K��ɱ-���:�߼��aI���    IDAT�����B�3��"KK*%��R�-��W�0��)���ϯd{y��8;GY�3l��aEY��Z�a2���zg\�@0HO�,��+�ͳ�_������;h���X�?��lN$�'q��q�	�ӏ��ehP�a�����w�:�?UGL�۬���o�[�� ~��7��)|������Zґ�$GU�b��I�z���L4*���<4ҏ���8=.��/�n�[m���{%\�<��]�Xp����G�HF�vP.ՐI��[����*;F�嫅��ư�� �������0��v�sC��
h������2>��'|�Z�CA�Yx�i���=e�`�uX�	ʜTQ"(ZP�IwIF��/a�=��hy?�I@��=����g`�u�:P���"^^����=��{��B�\���K�L&�ٓ��$
���<6J-�C	��8�W`�L��HU�hV�Io���~��� N9��G��h0�6�����������H�� ��@��]�Y�jW1��K_^�`�$�(Yߣ�k�������x��o0.����5���"^�S!IO$cO���(V�cy�o�|����HD}_*6�f�5��F�=���(��0XYK�屼�)��:>��
ZR M��]��E>&�2�r��l��d��M<�Γ���%D28�p�E)Wl��U�x5Y������nGG4 ��^�PG���X4�\>.g��D�/�X:��v��V�my�#0mw��Z���Z6f�����]f��}�zE&�`��iz�X�}0�h��bg��cj"�l2"L��<:��T��x��������/�����'X5�������5\؎_�_�` �h�P��y�b~,=\@q{˕�2�e$I���㏠e�\���E&zf�կ"���ԶR�����]��9I�"�����RP��E.��nO��A��2���7�3��6�Km߃F��E4�l�z��G�ƞT�|4�|=�D�)D��qm�<�����$�R�@��%�ٜFf��pȲw��̘��`��C(8�h��pф�\�6�/t�@�t��D�o7�� P5;h����Z]���� ��\����З�!�G�-��m�!ִ��2MCX�h؏`@E>A*�ř#v�j���vՆ%a9F��E���������5\Tш�I�-a��T�]O�):k(���0��������w.�gJR��-܅���!��V�H�� P�m��:�bd�=��Q��q��0Л�O���-�*�w��	�3o�h�|#Cju)�h��`�K��#�,ů>��"���s���@_ />?�Z��g7$�t��xp���'F�����U����WO���cuqM��� }��
H����-���ˈ����kF]{ׁ_�#�����C�ѫ�����#����	�ᕁ���Tz���!��V����~��>d!�:>F�J�G��C"��ܢX��ML����s02H�(��x�`W?��b�@�omDѲ���;�%�h��ɨ���b:��#r���>Tv���`��ơ� �x#�t�^F��tt%hv�XD"ҙv`�-��~�h1!�b)4L���av4�#���gЬ��f�=5��G+5|v����F��☙�h!
���A�g-��tekD�6:�- �JJO�T|V������/ʗ�uv���y��p������j-ă�y���R�-(�K�?f&3��<2Y6�My�2$m���C8r ���F����jZ8���~\��"��j 	�s#|咥�сm3�ԋ���p\���}�:�����UC ����1:���
��ӁÓ�c�YZ�
�b��HҺ�M��6p7U��c���h�.$q��F���**���K+Z{U�>Z�����D�<R�ɑS$b�7�ꚉ;�x�h�zu��Q� =��HW��i�Zb\�
M���24:���\�|!�A��F�����p-Bi%��G\�=�_��JP��#A	�5:��a����|Ӆ�J*|�cJ�Wo���0�,�s�x�G���(7�~5à��������+�L�����4��8n޹�i"<zP<���I��#p�~����Boԃ�<}��,>*���#T�ϐ�cb���0���|���.^���o��=�Ó>�mw�[���- {u}uÁI�K�n�'���g�`T<��+o�ֶ��3_���n�A�e�T�%ЀɊT�L�U��`pp$���9U�l@���ځ�k���/_(���z��lK'#=�HtU��2ݒ���U�G���A	��@Ě�ڞ���/��Y&������-��AO�4��P,�kδ@Z�.%�<�)a&3xtfz��ne3Ca��W�+"�0��o��/��f�Bz���(��Y�NA��]�Kr�x���Y���^����v��tT1><���~ln[��_|�n 	C�`�?��|m
��\�)`p}mO�1<��H��p,��fq��4��]ܹ����5YޱD~e���ݪ ��?�@�,�պl�#Z A�/���&:�:|j����с?���7�����*�"��w$q�M�2����ś��+��|���E&�S�B�]��h/�F���hK_��w$�O��a�b0�|V���;tS�j�J��b2�(��£��?�§�!�����ܽ};�;�=�ڢ��X;����H��"�Lɠ�t�;uL�pd��d M�ʵ��a��� �"����ks�XXۓ�	�c��q��(�6p��g(n��LBǋ�B��4�͇ٙL�+5��l�Q��痪�b�@�R�&a���!I�&!Z��d1�X��<���:톨��@ ��B2GqltM��+ �U.��F����|J��&~5JC9�����׫~�=��
��{�	�A�-����2�V~��Ԏ���ah|w��خ���/�x�tb"*Af�0�#3���$TQE[�`L����i�̞�7> ��H�ӈF5T�џ���d�~8� ;�E4Mh	�t�Λ� �[w���eh����>��,���*Œ�;��^���"�̉l"*�M:D���R�)���v6ٳ`݁AFR�Coو����&����zVt�� "!M��I�"�~lι���Ax�Ԥ�y��t�h�Ć[��9�˒Fz^���ʙ}���v�x$!Ϫ���j	ɐɨ_����h���HZ<�YV�R��93ȳ�6.3���>3x��!3خ����LAa���Ao8�X҇l6��.a6a͋�B��
X�����``������ ���"4�C�T}ՑOE�����M譖+�6m��' ��ؗˊU��� L� ^Q4�ݪ7Q*�c)h����7����J ,�b8��:	_�0��>�ss�$�m�BU^�M��+�dk���=����qJF��k��� g_���P��㔪*���~�y]O8��9.�px*	�Ϗ>Z�f����M`0����֐͌�7���@�/\���<R��l�ͺl=*:M�좉�qY��Ъ/aj8�C���/�x��.E�P�7ń}��6-v��B&����ҿ��ʏ�vw��V���]4mv�1�' �ަ�����8��hn�8��7}�vͳ|�:�*~�ϸqW��4>Go�'/�k�u7��`�����d(��҉}0H9�>$3��Xxtd��c�$)��]�aT�4Md�4�)�w�>��?���ÓU��P����ɣ���퇏��ut˫�� �����<@&�3�2��
�i,��~=� f��0<C$i��MY]�-2ֺ��K���Q1[�;u��}�M ��Ь1��M��,l+��]X]/T͇T:��^�2� ��o��Jv�5�[J��' ̭K,�bUǱ�0$��󣌁��_�-��v�ے72R��gGYQ��P6,�,�<��KP����2��A���b0��c"�l�U|m(�<�
2,�̦%���(�����l��O��ąd�����e��1%�lj|J����Ž˿B�2�}�M�����0:��)(~�A�dmX��8M��^M��H2�<�&�juc������Rﰦ"F���l:��
��P��Ф�Pm��mX�ޕ�V�!��t"��ޑJ��Ν ���S*²�+	#͢ive{�� ]ϸ��v�x����t׃�'�eJ(�D�_���L����M ��j�}���&��U�����dTMC�$c�A$�)C�<m���n��v���B8ƾ` #S������w��K����B'D��s��eנ�l
�y���2�>x��
��Qܺs��AbjV�`8?�`z�e��U����$���'P�k���{�*6�H��j�4^��Wd��㟽��a�R�'�D6�br��f
�b��H�n�����?�Dq��|4���"��0�@<�h".��x��<��޿�	�6w$���w!�ͦ[�bªm�'�a Ǫ� �>z^L<Z-cq��x� :����\d�hB���^�ע�����`�����x�*r��63H0He�bס׷���sϜ��P�8vtӃ�߻�k�籼^C�w�O�=V5�xy��!m0��đ�ke���W$i���_����H6�?�η�������)�c� YE �sQ��������c���"~�և(58t�f�L���|�8z|��-,ms���c60;��h_
�}���t4t�W[�����*Y�҉ ��.
q?�>���,vJ-$2!T�.n�oоqoIz��%�»Đ
z�4	%��(��BȦ���Zf�b��F�������a��?��n^�+q������]���a�o�A.^���ѣ���*���hp��$�3�=�O����7���G�5X���"��K�\EC0��<���l���/�{W�B"�Ǚcp�Ƨ�\$H&�z�v3���	�&D�౫�	9���� �p�cV��K���@����q��*M�|��-��N��đ>�7�:uh�Pک��W��R	J ��FG:zgg�š��X��m$S��I�V:(�ml�TDʝ��po��|>���tR.�
Yi�Y6o�cդ���,���^���AGU�+\2p�q��$����gsE0�p�x�k�_�C_�xɰ�9F��Y�Ӭnc��B!�~iz��:x��,�X\RY�9X�*���S���ߎ�����ۿ�'���IL{j� �"RI���kH�+ύc��.�}�L��{��^��5+%������>Fӡ8
�YFO2��ǧ��GQ�e����mZ�[�{�@�r���'�AoO�����h~8^v�^ܜ_�.W��q�a�<���W�����16����F��r��b���z��4��98�_d����cfP����X5]7 �ɓ��r�RJ�˵�@�@uѵ�Hż8=ۇh��xԽ���U<x�%�$%�]��Try���۞A���`b���ʏ��t\0�aϠ��Y�8�He�A$>䲬!*"��brd ��4��pM4�-����$�����K�+������/H�E�XA�A.ͪ�E��G`�}0ht��ڦ���]�kuD�	��+�Pk������`������'	�����g�~Ϯ��r����y�����T��3TF*��5�;��o�U�.k_���'��z	�Ҏa=b�q��ⴡZUt�:�~�Q^xA�]k[�(��6w*(�������o��R&�����B�,�F��N_���if��խ����{��2�Ƒ�j�ۼ�� �3Q�kwPg�?(��N��K�
?l�!7^�lJ4}�r�O�����3��Ȝ�&�^A���� s,���2w`�X\L�Hӫ�p�d�;���	��,��e�24�ڒ��v;	,�P�%�6뷙An��3��B<؅�a5����{3n9��#�ar� O����*-��8L��7y1�ze�B��ۛGew�L�����AS5�N7%3��_�?=,��n0���Ρ�L����4BJ^%BLm"�<�И��u�{U��-$�Q�=9���nbcu�RC�Ξ=�x�ص�5�O2y��+�>�Qo�'����h`�ڒ6(�v7E�	$SK`n�u��~��r�ˋ��]~/8��&^�t�g����N�=N��Q�Z)u��2�r��v�gn��cf�}�RN�{�H�/R4��5ae8V)��e~}n��au�����3حظygQj���d���A�ʂ�)����8<��k�~����t���!�-��.�c=�42C�am���@!C��N�����0��bV�	��m;��mܙ[�f�O0
�߃S'"�P�\��[7$��%�u��^I���pR���'O�̩<n|���W>M;/��Q�7�LI㟓^3�' ào%���gJ!K�=�M�&A7q�d���4�hy��P�N����n�9�I��	�i�0���[J� JW�E��C�U+#Jr���C��VBS� �Q��]B ���C��
��U0֡��)�R%O�2O;�vuw���k�@}��.��`]�'�w܀j���Az��Vze玌�O_���+k���^AjhT"��(.�S/����w0=���~x	�K[H��R����Oq��#���<��bgk��H�y�_�ģG��K'q��'R��?�����x��w��W�SO���`~�������H�0�;L�u=G\�t�w�0=����>̌%��� �&ps���7����膅�pG��,�� ��ݔd%@��(q���Е��~0���O��� NÝO�Kb*����GӸ3_�k��hI(jZdZ�+Hj��ʶ)L��O;�R�?�)��e��L���_���;�m��noU�=�`jf��)���t[������G�������Z�g�HB�\�����9̎��?��o�6���p��i��`�L�c�/��;��I�νۈ&㘚���k�G�n �^��5,�}�?���8}z�^�����gO"�֋|�'W�0��a�4>ٜۦ�҅U�Ao:���$FGr� a�P��F��m���.*�J0.�.�`)-�I�ա�&8添%ap��u��K�bu}�T���afV}p�M���{�����D,�|.�'OIE�Ƿ6qwiź$UJ��3L�s�������׋��+����XJ��3��s�:V�Vб=�>�eT� *z��#�7�@"
�k�k�0���/��$je���K��������f��0t�2���o ��+�]C���$��F���s'ቓ3�u�����z:
�m�<j���
�a�Q��?��Wa-ܺ{�t�}#��y1�b��w�"ɡe��K��	rY������`����q����>ċ�rkk%�*ua,2d����Ŝ�r�*==n��3���#(C���XB ⑾Nz�j�:|E�Ԯ����A&A�+��@����p���n1|E���;�>��Oi�~5�8�0�2.��~&%�09y�ǟ��.�$d��Vc����	|��C\�����"�Sh���XE!������]^��%Tm ��ay��N/>{S�}Xz�0��x������KW�T��e��~�i�p�.��F{�����6>����jS��	ХYX�F:�k�Y��i�!��m;�l�-K���Ul�U�Q@7!I����\R��|ݴ����JI��?��[��y���`q��@�.M0=���*�;�(�?4$���*,�ak�v��&��\ ��#�����D&��/~G߁B0�RW�2��#�;p��!�`L$4�3A��M�]=9;�e�֭{�1$�39�vKl-�c����Bss����$���"�Ī"Y�&ʕ�-��E���� �DԇhPA&��s<,V�H��������:�&ߧ0l*�f������@-.�-x��$ϓ\a��x���\1��0HȂNgg�X!��Q�rRU���0x\5���>�ȯ�JA���9�F���|c�9	�d�%��Ž��Ԡ7���j\��� �f�����'Ȯ�Q������dZ��{����8q,'����&�ź���s�"aDR(�t\�8��q�}�    IDAT���¾�:3�t�����lNt���i�4����g����q�C�-W�����K��������ru>0��u��|�%�G���Fcf��;���Mj	t��$���Bb��/Ib�<��BdR,�g,)y�CQZ�*�K2��x��ze�c �7�����(b�\F0������{���ɗ��/,D2�A�[�������Lt���`��}f��/�WRPR#�:�����R�]7�"��㯜���.��^�"���\:�20ޗ���	lm��������8sb�9�@j��V��J��͝��w	�Xa����C�ȥ,�_��H�BL�u$~��u�Y��U�[i��< 6@ɿjHE�Y;�.zn�Ltڦ������ {R����`���@�j����"�l15Xp}�Q��:
�m�+�`��@ :|�����A�:V#y|�� �^�0�7������srX���i���q��/�?_d���a|��L�������+o��4Q}C6����=�;��cϊ�E�0+iq:����`f6��{+��[��v�&�̀��P!�������_]��ɦ>S��xrVC&���fQ��[���Oz{�^U�%L����TJGCo6&�,�4QnY�4�ޫb�hʶP��:L�s&�u�D;�~2�Mta�c���mp1�`m���bfׇp"�~y�/�����W��ԉ�^Õt���0�&|�`��	��z�j����8��.��d�}�(F�9u`�*�l���{�������~T��0-���' ��ƈ���b�p��[���"���1ؓ@@�`��m��f�g���^��R��!I/ocf8�?��,�{����:#��	xD&�F����D�y�y$����5<ZځLHEI����y|鹳"���F�||��N\��P$�zyKΣT*�/}�<��V��S��/�ͻm|��4�ޣй>�/�񢥛��$�}wgg�N��'��tQ�6���$~�����c�uT|�gW�Y�gw�WE��)��P���3����
 㳥�\>3m&��=��$����,a�m ���������
~���I�D<���'�~�'�q�n��u	��|�(:t�q����\w��=8w�ڵ*^��?�[�Ɖ�^��_!�_�_}�+x����ZDx`��h�)�'f��Fa��d7�/?�/�����mܟߒ��p���Ayo���8{`��?}�\��_]@�gz����"21���?��tvϦJ*X�>�t��D��ڰ�U���3�����fǃ��by���Os�Jq��ڣH 5zU+{����x��o�@���ހn�q����H�o��U�]��L$R��ѪU����Ij!�O��������7WV(o�d�1`djb��_�	����:)����������!lnmJ��ѓ�1t`
�^y���,���F��sd@8X������;x��G���x:�'N��ݛXZx$g����i�����;~��	�q��w�"�����q���/��K�=���z����wP/���|g��w��cl�
s����}���©ك�k�kC2F�
�ta�f���[����/?�H8�[w����	��,mm`����G�m�h��*~i4�Bf�ĀYG<��ԡ9�{-��=�vatlܺ���G��ʅ҃"%W<^�ًC2;Q��;������J��Rj'�!����97زdboG/c�?���ø}�
�V����=������pq�?��6�Ds��ɥ�3�\��vqpdTz?z�U���}(���F�gp�$��'���C.�HTA�����8�}r���g��2X�b�
����T,��q�h/��x��K�9
b��$kf�~<qx��� ���~k����llm�H�p4�!�p�`?�� ��U9�H^,,nb�X�O�QbK��Jɠ�2~\t��?<��G�����ޭE	i"�ɴ���),mVq���M>-�Y]�_mKҧ	�I�p�jp)!��\����\Ĺ2���C�u�,� 굲t��>>����O?����u��		!�eaz�0�����/`���k������� ��.~�����~����;���څ�f�O�`�0|��$��i��l_|z+M�����{N��z�|��2�4�z��q�T{�0E�U�!�O�Z�I�M"IZ��]ܝ���h�YED���ɣHēX[[�����^,�[�����*��~�����Ֆ�1���+m�dc�8?0�B$�|/ʕ��g�\�p7&��m�
�du�<-U�ST��D�/d�c�;��&}Ta�)A�.$��
G���L�c=�l4��E@c4B������X�,����vE]�0��&�z��L~f��c9$�)IM�e�x��H%|x������C�ؒ����B�j�ñSGq�N/^E<C���@O }i�a��,�}�y>�}b��}sčȑ`&EJ�)Yђ-��;�W�SS�b�/�w�o�Ŏk�;��r�F�(��  r��͡��O�>�g�|��լ�(Uqѧ�����y�#�z�ث��4�(U�(7[(ԉ$o!��1��bl ���hZ���a�Iq�nm���|�u�����b��6�d���=d�QdѦ������z�3��0�=�r��� ���Yn��ṜzP�F����6��f��40<�4�P}-?0���8F��-ö���Ǖk�(�����c�5]�fX��ԋs���*e=j���g�����fPM���c/�g0����P�$�����l�l�G���=f�f~���MN���1:����n��EѪ��m����y<�d����nB1U�!�=���se��1\�M�K�y
�j���bv~��C�\�������Tudb��B]�Q/������,��m~n�����z��.�A���E ��*}2^E�gg� t$��h�m�������|�k�h%�q�B����f-/2��>�@Ž�L�8��Ӹ����wq��D#p<������K��ے&_�ml�?x�ο��������ALy�G��T�z���Pn��˿���*�!4�����UX�]����
�9��;�?�\���n�iaXqr��􅗱���F����so�Z�xy	���U�M���/?���"Vַ�x�(�C~�Z���[�yoM�ĭ7��a�۳�g�-�4zؿ8��aL�hT{�)�Uܼ��>��fGC0���0˳��C>4��-n&<��s��~t�En���W$d����u��IK�׮#���N���X܅ը#�Lch(�j��ُ>��;p�(O��ʃ��4���-}�j��4Q4�����]�Vocx &���;�Eڙ>p��Pb��3h���]��m"m:x���7��v��*~��'hv�2�8<;���0�R�����޿��^�?,2�CYLO2����.
9����]��G���e�����Ӈ1>i"`:����;w١q��"��A�f@S�j�9%���H	o�c���Ҹ��.��7�ONЯb'�����?��g'������S��f�-��	O���-x*,L)�h��ꃷh��tJ���x_>�d�`�u�������{
N����#��������������Cdp���p=Q�)sm�!tmF���A7�8u� :�~���E����Q?���ۈg���Ͽ�_�y{�{LCr�<�I�&D�Q�m�f�˟;s�.>�õ<6�M�[M$�~<vd'����?���.\�iFe�p������P�uy��]�'7���z��|~ăA�x�i$Ṣ�࣋˨V(��.�K���W������k�����t�%��G�X�������%��D�|��/c��<^y�n.���JA�"�^+��'$��ٓV�{�!�a"��}��M৿�.�fN#��?{s�1|r��0��?�.���|3GN����-7a�"��N7���R��BX�ppf��.^������o#�	�S�q��ܻ{W�n��N#�T�MH3���H��."��_z
#�^���u��,����p-)�������t���P(�%N� ��3ӣ8z -��r�g�[[E��*X��V���l���� �22�)WZ��+c��ƭ�2�s�a�0�ӣ���ud��W�h׊кu<��"�/&�r�6�~r�@�C9ϼ�,�e�b��?�J��a�&��t��5������PӍ~� )�*=L$���~Y�t�2g�$���+�K���0><�VW�02:�z͂Gհp����ֻw��W��G�v\(�_�-0��BE���f��[��s�������B�̜�!BY��$��$�~��#F�cY,�+k.\�'�^ā���W�-�ʭ{�hYj<��>D� ̮��.�Ju���Mx-�D�:ff��̇F���^{�:r;��O}�_�GJ��*/tmƜ4����
8~hO�Lb�a�����q�NN���ceےf���x:�W���h7�b��5n�8'A�+�6JŃ�b�Qh9�mfQj����#(���8!�F�.n]�.C�p$��n�iwp�gK⽏��CU���*�Ty���s��i�q`f���g?�;������.i���8̱9-EdxJ��Ѱ��l����W�t {;=�}�=����N.���x����������QmIcl��M/���P�B�f"��Xk��jW)o�\�����8�֚0Ԡl���6v2Pi9
,�s���'ҖA��۩cd ���.7��PX3�DcihzW�l`m� ��65�<��d�'!�ŉTRfDR� ��O��.3��R����]���h��885,��k�?�n!'P�X,�T2���\�n.���"�o��7��¤x�X�O��L���E�%�os��f'��/��J�����P0Jp������&b���[�/۷���נ1Sů�Uނש�'O��S�q��2\�ãi@m���<n޾�n��^��6~���p��۲y<xt�����kx����K�� �q�����S?��PsidHA���&���Ғ�KW�Q�hPIT=y9��v�U���&@���$�L�ÆL��{�`��e��Ҧt�Ϝ>�Fu=�!���t��(�Ws���l�6��ա�d"C����2-�������a�n��{k3�K �Ly���3�h��H��n�?�����,���1�M/B�X��v�p��2���_���	���^�õ&���V��疰0��^zv�!Z���A�b*VsM���m����$� h�����u��A���ֽ-���awI��4�I(�ܭf�H�*�F8uj~�5�	Y��X�)0�qܹW�;�]F,5���р&���G~,h&e�]��U�7���	L�"ͽ�DY]�)	f+��Ş������W^����baBA�]����������͸D-��f0`(80?O��������|�Y��끻iFKx�b�0���f��?/�H����ן�F��o��wa3��GP�+:��&v7�����7����_��Yl�,Sԋ[��phz����cym�J���:�4���[X_݀��U+`zt �Ã8{��C���7�W����p��&V��p�04#���N�J�!�B�k�Y�ĉ�3x��Yl��$⁲��C89�ɹA���&μ��d�zD�Z	�D�Smf1�ZI4�H��1�#x�;�oJ_�1躰�m��8N�r�F���3x���pᣳ�Ld�$�)�8�����'�a-߀HAƤY��^S���D���s��vq���p��YT�obp(��b�2Q����㈎�F03#��L�^�
��G6�����?�z׋��e\�u~ ���`n*�{w����ZPUN����N=���qq��ml��thk�3��<��EB_1>���Lmo^������%(�_�c�GR�L���b�,�i��ן>��"���t_}y�������J�]�x�(N>5�;�m��W߅�5`�tI�d3�v�&U� ��&R��u(�y��,�K��VI",�4Qr�vM��÷^ƁEU�8��]����J�
���ZS�/~�t3+�v�D��2��#w�+�An�;�~��C;��#S��o#�	����4�[�����A72����P��A���]�c�G���EL�?��&�}r�J�f��_;�L��3g�q���-�@P��/��i/��j�����ΕD�S��3��"�S��!�̙��j���e�u��Z��=�3�(ך���],��|:�X��������ࢉ�v�����<:���(U=����+��H͠��ݡu��Ve�dL�56U>M�pT	���{��0�����JP}��0���:��K8}d/�p �� d�po������}n�(�Z?y�C��]������""�Z�E��D�����Qhv	?��_���g����Gq��%ܽ{N����(�:��4�SG�NBFe8E�I�[ñ�A=8�D��^���޹���-ɓ{��c8}�/����*>�|[>o��MN��g�Ѳ4tm/�r{��ʣ^s�ߵdh�pzm,���҈4l�ױ���z��[w�a�h��.S�S5[�>�Yghu����]��������L�/_��O���l��x1�o���g$F��3QkxaŢ�8�#t?l�֜P(*�T'qx΂�o�`���[��҈��`�$��i��M���"�]�127o����*F�����ū+X�a���W�P�~V�BO�4����7����3g�͠[���f0�	�fNbh�$<����̀�v���ccav�S��m��s������8|`?Bf�[���F�tZ �šc�����nk����U#p�|6ab>�CF�0M�<���l�z�=yM�J���$��I O_��ͶD���e�1:�S�1n����&�__�����I$�tcV��� M�˹*wh��M��ߨ��I#�D�!��~��oi�"������:n~=*굒�*=8�C�T�0��'���oݔzjv�0�������� �A�>��ᖞ͠���H��]���~�'rŜ��ţ2���"
#���"p�����e}};��ź�P�
[�?��ረ]���8��U�<S����N�M���ȡ\��R�����v5�.����L����j4���*�+T��[D��EGJ6i�Gq6=�Ni�淉hPé��zp��mܸ�1��&��0�;���1ܿ_���hXb�G����6��FxP����C	��4������]������E�?kE/J����d���m!�K�[�Q����sַ���S�8�_5�2�{�38;���2�)t@21�p8��e��Mॗf��T7ބm��3b���e��V18����?����~�O�i*h�xY���=��9([���C&K�p��
�\�&S�۪��g�����Ւ���r�.]/��RQ�D��K>'z���#R4�*cv��~jF���k˰)?�"u������u�c���j?P���M$$�1U^&6f�l���i���͠��`U�q���G���O~�R��T���f�061#E�;�_C���Ӡ�A�S'��.1�6�##��ܸ}��ۿ�t��$>��F�M�a튷�?��������;�q��*ڈ�g`5�rt&��30L?��ul�ڂV�UL�G�Njx�Ytm*e�\�`i5�\Œ\�V�F$�.��K&��cG� ��y��r�*��Q�R�����m���̗_~'��p杫8�m�!T*�`f�'�\�f����2������^�? �2�Y�^z1]�01���=�}�?ۿ�
�cK�!�S�zYHl�)�::��_����v�6�P�6q��8q�q���5llWD&J/R&z}-��ԯ��nZ$o��.]|���@}]��0��;|SG�Ff�����X�8%��7_B0��'?{+�yt�:t#?��-�F�嗞������~���2TB���O1�����)��h�]]���|�.`�\n�F�������bdl�G���u�l������\�    IDATðʩM�Z@B^U��)ǭ��|���SO���ŏq��E��&��&f��Mܺ��o��U�X!H�KB����N����C�q%�	�&��K(� �վϐ�n[�&�!���ZqW< ���.xK�oalt���\���9|�O����p��}����ҹ%���/��@���S��Ƈo��ų(=����6>��H-Cxx?��0��I(��Ȩ�J��J�3,�M�p��u�J�54�o����=nZ��F�Zh*��>4�-�+u8��p0)Dצ�Jq[�5d#R��X�Y��lbxd�4̂��S�P���D�R�"Cd#�Ht;����ի�-,N����i̎���W�c{s��ϞG���?��P�	8�	�� ��k�D�M�I�2��j�WBWU��M.e����F���Iz��9R(1����rq�S)�Űz
��t\�x_�_���@1=x��.~�懈�&�3C�Y������}@���Yt*E������ O�+�����◿�_���Vv�XD�2��,g����4���a7v�t�H`��n�y���E�M�B�3�\��*�]S�K>���'h5�X�ܓ���<+��BP�KE
�(Qn6-�e�N1�Ц@(�`(�J�.��Os���*D���$�I!_܀����3���� >����W���/=�����eܸ�*����Y��o�D������e�+Wp��J?2�rx�.QP�i�#/�P���Qb��]��-!�u�J���c��s<��w1>�A,��ֲ���;hv(�V����|�m�Wrf;�6��bvt �^���;���HeL�:�(��ʊ�������9MG83	-�'�y������8�\Ň�߹���mhJSS�e@���#Cl�̮5����?�Akk�(���Ыg�0������&,��d"�ᬉv����m�J�¨T;0Cixn}̊@�c�ު�04Ă!���\d�ԍ��~?:���F�{z(��G��l}��C<XZ������H�%Ǚw��/5P1_Ev`�.;�>�o�P/�#H�dv.�DKПρ����*����~�B���kWoʰwpd�l�<s;��ж�-f>$�����e }���_� P��6�`đ�=��ٓ@xj$�D&��c�yQ/��p�29r{9d�cp{!$�i�[5�9�� �^�І9g\x�QǟǧB����
�jK,l�I�o�u���$�rq@��l���z.�t��u�*�̓V9'�����eQ��8�lۧ��P�5p��-T%��R��PgM�A�c8�p��U���D*�JՏ�yy�3Hi"�**%ز�z���H�uL�����e�/��5�oL޻;K��p_ @���^$Ś�Ul���B�v���>z�GB����c,�4�cӲ���{6
#	ŵ8�0����ĵ�jm\�� ����<��qD"ln�p��vw�p������T����*�����v�����HЏ��ID�^��UQ(4�W�0M�����P� ,���GS����6�6�t_Wb�F�B�X����5�{#8��(Llag����ǜ?>#Z��TM?�!�bSF��}ʳ�MEūI�F[��zU��8<3���Ax�M!���lN�!����Ç�I���e�U;��f�Fo߰�H&jaz8��f0��F�g"E4�^n�d/�x� ���í[K��)�{h`d4�C'03;������[HQ�)��� �&L�e��B�+�lo�b�H�|�&7&��8�F2�D8�`y����T�+��3�i��$N)`[�6���S����'p��^��/�jp��Evp ��Ͽ�;����)S�tٺ�>���8y���,(6�eͭJ��o�2잗�]���O��ho��5ح62��.��j���q������WQ�9��Bq9H��3K	�ctt��.Vo\Gn��oo�A��3�''Ύ&�&�jTptn���#��aee\��õ-���G�GQ,tq��>��$9u�$Y��O���$9����2�e/��7v#��D������~j��J8��y$�i�0R���Kb}��f�BM�c�SG���V��*�s�}'O�q��u\���V.t��)��⳸v5�W~�+$�S��x��T��jn][��>N��!�_���h��K�k�L�_L�s:�0�Z�M�g�9��������$gp���8�4.�x�;�֥t�`V�����u9����Sp�4�/��:�%j��y;}��o�0&�< ?3�:�4�{8u� �������.\x�r�T`r2��KL��5�U�y�`z*�o}yv���^k�M�j.�7ȕ�h�[0B{�q��?=,�+�ZKK;��̣�p�/�%P;'4(�c��}�5C���#�j�x��#x��,.|t������f��7����N����8w�&�q�]Mzɨ��I��I��$��ϐ�p)Y����<@���B.;fd���F�ݨ"T��_9�����d}��{�y�.Y9��vj�|kYd�>#,� %w��sG�
}��g�ѩ�����{ps�è��\Y�����?�������	��1t��BG��|݆D0�C�R�aT�����A�'�P�D�$3F���"��5��ܴ+�\�oj�X�J�p[-d҉>�U�а�yr��I=���5r�I��E�Ve?K¹�s$"���������ÇQ�HE�C���	��}c�M!�bp $�𗮕p����5@�)�=� s�0�^Q��4	#�27M�!�_���º�'L�H��Ʀ&Q�6������EC�h�^t��@5x	2�������S}��+?Gq�N/f�����$���W����}�s�e�X���У	�h��4��[r^.e$����%���N�y�80�q��0<��j� ��FU�F�Q���^Wf :�S��k�Т�Wo�0ZM��%q:�KP�F�[%�z$QH^�ѓ��y�����k��{���(�KhT����B˲��S@��g�&�2Ȧ�H!���{�|������^�-�K`%D��*B�K2<��xd8��p���J�^O��u��!��Vc�bL��^K�����Ն����8R��`�ص:0]��<��ě?��>�:�1/.L��K�Q-�V�Fa�12}��>��8���xm���:t��ᕳ�gO�x�	㐄q.t��0P(�JN"J$��ݒ��_�cJ���j� ��y�Q��w4��L���v�{���>�/�V?v)FJ�mˆ�Oz���ľ����Yü����	��f���*��7�6�0F�ږ��H4 u����"�n���!n��8*�O��������#�IF=�B�x���
���h6BFWb��������ѨВ_;s�F�HͶ#l�>��+�=�lu���D��f��F����s'04wnxZ$�D&�T%���v�$�-�Hc���U-��l|$J�)��9�'�4��
�y$n����ph*l~��w�P��f����y2�Ѝ�9Ư?��^� ����d�R�M���� ��v�Z�]�!�aumf �D*���-���cTR4�D�#�#LX�iBӀ�<p{��VKh�=/�WZ������~��26X�v���V:���#��xȔf��#hƋ�@R�#�y/���p�����3�-�#�?��f�.͠�����->���r3�6�n�fЈCۇ��#�f0A(��ހ��N3���" ��Y���G�ڂaFepğ����\���R����PZ���Z+�r2\�TU��)-ou8������+7�<�:��H8
�`|\2���$��'��Uj�
��.��f"X������N���� b�v��Xz��e3L3��\�/w%��ǟ;$~c��J�|>�Q�KQ��;�GLH*�V~���<�TK{�7��H�(�t����"��7�V��[�|��/�ޣf�2�O��}Ϡ�q~ޟd��A�Ȱd��+yx����� 2aܻW��[+X��D$��s/���Tp��-��T����ez��a,L��-ܿ���ݢD�Ju�ǧ	c0���� r�5�,o`7W"O���d��4��=����-�P��40�����>>�r���>��ڊL��/��s�8sn�Ct��!���#Ŵ&E1 _PE�y[D�3㍝<)P�~@�Xx=��������)�͂d�4j^�ꭷQk�e�><5��޹$�������n�\��_HA��F�B[����j������γtu�������q<q|�������%|���C�U��A�n�Pk�d���ő,f&��-lP^�^��j��(�>����T�E�f�c趻�w�>|R�٩�Hg�d��|B���p�:�*��K�O$�[&�Ãa<��A�����M����B,��g>�L�n\���K0͸L3=�tz=��l�@ؔ|8F#I4Zge�0���d��f��se�mD:j�To/<{�D�A�Z
�}�#�����`�A��3h�<p�,�3R��� ьl��0;����'���򥳨������pE�(��>M45� 1�|�~^�N�&����S��:~�ӫ��`�_ǩ����]ʋ�J>�fC�I?���zvQٳЕ"EA$�A�Q�N<��O,�c{k���/�a�h�% D3���m��%�ņϵ���E(��'1?C@U�_����	,��چ���^@�� J���V�	ʞ�*���X詸�`Z8��Ą��Fd�E'7���p��K�V�q8��#���20��0�Ļ�ܖ!���<�����o��0D>F�����#Xƍ���]�ƃ+����"�t���Dʽ��
�F���f�%�N
���Hib�&t�FK�B�X�|ru	�j[�;����?6��c��G�u�d3fo��
��#��j�!��t�������n�0��H�e3��CG�Fa���2��^�II�� �\8Uv�}�[ǒ�Mn���8Z������(BA]6X�dDȐC���V��!>��[g[8{��%k���W�@] ���r�����S�����;1�N��kϣcY�w�=R��%k`d=%
�E�e���	�3ḑP1;9�^��_{n��L���F,�W~��x��X��%�鱃p�42�seQbΝ׋p, �ziɸ���}�Z]�$;$CƵ�_NU`j��R*J?3�E�����?R�3��dAʶ�F!���+=4-b����)&�I�H�C�my���)�Ib�v�ߣ���_A���f��p��~�4�ɹ6�RJ�1�b8��z��C���rz0�>�_�����Q��}~�e
��_5���s�Ƒ���|S��FiϝXġ�(n�������ws9�K%tz>N����l)ns�������5ˑfpr �Z8��?����@8����?�]�lҳ�!�@v���!��Z�O��,���mtj[�Uv�/?�o{�<v�x��â�L]��p$���e�nJS�H0̰p�ݑl���m��d"hY��vaSɡ�IW�5��QBJ@��A0p��qe���V��An�]�H�׆�ᖇ��JM \��vw���U2�$���p�	����� �2�������`53��5�v9$;��q`���v
C6�*�5UU�*�Qn�>�m��G�j�	�0��쏤��W�l�h4��ݏ�!@�9ǹI����o�]6�.��6<�\=���	���&��,L?��L?!lmв����;$���޸(���xE�̳�Ѱ� 憌�~z��-�'��[�G@W��ׂ�K? 78�xΎm��-y�唍4�G�!�X�5�?KP�a���6Dê�K���ǎ�V�E2nbd (��T8.�� i�o��?[�@@v{�&z|�=�o������G����n�Þ'2v�	M�N@�Q�!0���.
�"��&t3�Hj�Iw�a�0F�~���!�=��(Wqhn~x�{�7αl��%h-.͠&��#���7��j2�KV@Y�.��u�Zu����2�`0-M!�9t���~�D|��=�MT�6Mp�����o��Ư��J�F�r��uW����ȳ�z�� ��5>�#q�.��:Hƃ����v$fY�R���f� M5e�ɁG �G ��+�Ҟ��l����b�r�η���~C(͠z�Be�������:�"�!��&�Z,�O�^
�J�.n�[FOK���f���j����Ѵ��g���i�R��~��#���ëש#��ajz.�q{[�R�f�� ��Xy���^[|x�̨�0<څ��a+�.:^�<<#_�F��XP��P�f�B�JU~PNY�KgK�},�W�눏��op*!AB.�84��q�Լ����2i������^?s-KA�jK1�G$d���ģ���jȕmTy�	��an! �V6�����C��moϝ(��NEp�D��Jb�� v6��|�
fƑJ�ʝ�<�4�ҿ��JP��r-)�)E5����7�{x��@eh�s%[�LB�g0��b#�g��"R]%������b"3zllhh�-��q)�*�:|��.��5xl~�B��%�8{�>z�x�3�Th���e��)64i�mģ!T����h���0�H9�{}M ;��jn�Z��2�Meq���A��z��(&&�q}�;{p��@�@��#����$30<A.���w��
5��k>2����$�����r;B�d�P�U��`��.�&�ɤ�`y����Q����//H���/�%ů����f�g3ت�ʹ7�����f��͠O�g��8����1���op|��<��L4�T8���M�m��&z�T��;��"�Z�]��ۓ	s�ـ_ե��ߣ!M�\P">�
Q�rџ�h�2	G����z]@-�ni>C����Y���D��v(�7�03=��?����arj�dkkkXY^�ߤ�J�q,�G2A2����B���_�{u/�6�4�
�:�F3>8Wx:鹭T]���ߠ�E�V���S�"��������!O ���c(x��9>Tx��"��`]{]�Y�C�����d3�{�*.N!�����`�10D�N35�PfJTB�UU4E&�y5�{�����y,�����*�
�Lë�+J�CW6��p�:}u,9�.�a����p�GM���<Ύ�U���\;�*��bxrFЏk�ʶ<��o:�B�RF~oG��>!S��}9�"Rk�S�3�So"����QO?��pȃx��T^�?T*���~�^||M���j��������4�B;�p�)��ގ%�}nJ[���{���Q�M�J�R�JWo�D8�A86��*V?#�n\�Cu�ʁ�gH���� Ь�������|
?��B2�׾�U��.-m"4x ����i$�D�q�Ŷa��ML�D������x��w��)���j��x<)��U�Z<O;�p�hy4{i��l؍�la��	I��cY0%��[�.,����4S���%�	�H@����PH1�w��3�q���.�m6�eQ#���ۢxh�Z�O��̐>��VG��"�@T{���@��.^}�#��4=�l3�Iv`�^G6���r��Q���h���c����c(������V���@j�?y��|=ŀ�j2L�i49}�����d6����ۯ~�ν�DR���q\�p�rA�L�3����4���!����b���5x{���^�/b�����e��&��z�IV����3d�2FǆEo�H*m�T[������Z��9����\X�q��bT��'�\b���iT[6,���Ϝ�V�0�&E�R.vhs�X�+����ֱ1��"lc)$xV�e��A�^G4No4�9�q{i��0<z�X�h��R��$�~zU�l���Ye�'���$��&�vwвj���C������zz�{5aN�9r3�Ϝ�ܟ [�A�����u3H@`��f�8�ǀpZ6��tf���    IDAT�	K�랇�bUx�-|���z�ӟ�G��h*k�^��>��b�p��W�Y�*lE��p�3��&�!�&��G� ��-	 _\���T.���W���`�c��4�;rcD���$��:�#�Xu����@"��>X-��N��HV�,M��*�,f���&c���G��ck����a�n�����fP5ؐ���Q�H�L��+��O���v֫�%�ؐ���<��H;�?~����P�[Svf�R��� ��|�;8����� ��(�����Z8���4<���O�XP�!�/��v�js3�G4��l���uHi��'�<��j(hw,t���^�V�J���H�����!t��_�>�X�X��y�l�����IE%O�#���a�&�2aZ )@ֿ�����I��E�O,�.�f'P�ͣ�o"��UAV�~��UX&H�������h4�)I0���LGV7�ō�O���N��Ѥ��Vޓ�@�v`��Y��E@g���^�G4�~3(p��f^�w��"�n�g�!fX�<hԋ�ܪ��Fa3@������6TO�^��l���פk�ux�N��Q�Cj��H�+Q�A��K�FD�
��E�vdE�e˶d�N���*���E0@�/�%Ew ����%��	LͦDʷ����?��Օ44D4|H"V�Y�^���F�_��t�+�7�}�}�)�Q>ʑ,��.�p%�޺`l-,�ĩT�`f~�_��DG�a����˥����Ӧv�&���1T�rX�~[�o��r�n�#.,̘�Mf����Az�(�� x]�(q�?��s�H��3��n�XiC��T�;��(\��@�*��F�"��b����E��z����D�[>�+T��-�I3��*�Xu��5�a1T���*�ѱ۲�:�M��.L�A�����t}���vP��a��3y�v0��btt\�L�h)g3����'����-�ӓ`�@�`;"_�G>�>2�M7,d��F�C6���ŷ��q[�@��D�K�v ��(���{��:U�t2}aA�m����yil\z��D��q)�!,m�(&=���zJ�?��l��&4��Fq�H �hX D��#xx�0�(�DS�68��Ql��J��v:r���Ii��{MB�]��Z�����q\tX�AN!��;�y$��m��NҔT�
/�2ڍ�=]��\�#�a��x$�t*.����3ɫ�4��f����_­�&\%&R6��d�)����Q�lȖ������fE(|�N��O����B�*b�^C�j!�ɛ� JL����U��sd�d@S�09�Vq+�/�օ�(,]��C������A����LM"<0%2�J�B<C˪�0h�ϣZ\×���||���J�
»\��4h2�ڋR���Mhz?H�>�a!(�! �pu?���A����@���!/��F��x��۸��E� ���� Z�
ŜL?e
�A��*}Z��-�hEX�iP�{;�ï~�*��D[�H*h���mt}&Դ�������{h���²�aT���y�)"�F�J�\�%�dB�3OD4�E�Q��� ���4W����$����P(�Œ����L�A�b�
&F�i�q����s�*Ņ��������?��y�V�CI� �ݏ��!��0"1���-m����C��������y�n���?��Ąxbr��4�lq}��74����,6؞~3�j=��y)�cьL��&L_?�[w��p��)�8=�����yw	5 D[����s��Re���fɅ�h����G镏��]��:uOOB�泲��n �E��خ7�W�"=:��B?~�=X?zz��O��"��F��(eg���S^تU2=���ppf �G�py���d"�h,)TЅQ��߽)~����]��*�6�]�PzULeS����w���#�82�K�GngG6s3�Q���'08u���F��~���Σ����O?����{?�"�3��#:t�1~���6eg!9��*_��u,9�����eנ���H&��5!�j
��*�~�4[_��z��Xf�Fm����+hYu�����g�b�m�4� �g�K��q:)�_|����YH�&��%p����MD)t\^?s7�MO��"(7Z��]�tڮ%�H��_㖋��LME���Y�����;ShVy&�Q�Z�+�(W{H�p�^S�R=ܖ)�|�M�y��l�<N�P���*>z���AP�IeF��Df���l�P#q�2~�j�0�K�7�d���{p�͛�+��U�2��p�Pue��:4+�=�E��r�)Bc�\��c<�&U�����������ه�Lm��۷���,@5��z��V[�C��	�Թ$Z�ea���&0��-��v������H�|kY�)��t�����,���������U�!���Nb�ȿ��@j�]��ؖ��~#�f�85�<:��A�;�B"1̳�pD�T�������/�f�!�~ʟ%��uѬ�qtq~��+��>x�{p9x<M�q���	�\\8���4�L������Z��s9���S�g_|��o�q�"��8�D��ݗ�0����y"}��$JIy���l�z�7`�L1�T�9!�2?֋R�!�v�`�r��{a�gG���+J ʃ5͋Z���cC�Y�����������1�]��$�R��.t?��
V֛��%���!/��@��d<�p�M̚�%��^����,�Rړ�i��B�PG�Ґ)hF%F��0�R�fP���AЛ�������k!�Lv>=�` 	�����i�O����	t� ��H�F���ύ�� )t�()�S����Kf�:�<��*���d��_��'~���/8Qo6d�m�2順ݥ���M�\��Hs''m����dR�QmX�ῳ�e�6�b4�B4D<b
������I�{��~q�īQt�*T�ҟTӌ����%%���a��6��[��H�*.�{:�W�Na����G��x#p}A	b���qBkx���HȆ�����W/c��'(���؂���GC�-�����؇��g��p
��@�ן����]����3��?�k�M���"�h�mX�H��NNb[����2�K���\��H`U%���)�`>e���M���������v���R+o��M���95%�P��9V`�� i\�J �-LF0��"�z����%%��Yo��h"�I���ޥ��e\���@bXТ���B��䶗�tN�ۭ��{<��"���Ock��vs5�-��
J�f珉��G��%�[�G�^����6~fj�N�>d���hm �	���rؚ�'1q�Y�3s������y���.N�Aת�ԑ:4���z���019�&	h�������
��r��0T����&�]"7�|7)�����)�C�4��fP,�$҇ ��4�=�
���\Ms:�.��.5N,i(Y	�p)�*��k88?����:>���wjŚ(�
-����n�7�	�9�<脜���E�B��E�V5t�U�S&���O�ﳼDzN2O��
r�=$�Y��i\����L��qtG7�,�����Cy{뷯�ڇo��~K<������\5�����`f'�=�Fa�	��b����X��z�';��L�:9�Чs�H�� ��L�ʲ���FO�������L�'�gֶl�-�b��	� ��FF��F�prλ�s �S;6�\R�TE���|��<�}_7��Gl���6���3K:�∨�UK�YQ��]A�*Y�X]^��p�u���-��l���]�%8�w�N����a�N�����\�.p���ɒn���у[Y��2'6�f���6�,�<R���h�*`���SGwqpO;�|�F�J{�O!˫i��*��4ѾA������Am۱Z
��Lq���x���`Υ�]�j5� �W_:���C�}��� lS
m�o�=�z�W��//���#��G.���|��m���siμ���9���y�������:_�����%�����j���� keɑ��5҉y����^{�	�I|�-��e::%�ў*���%�x�A,f#�JV�ʥHYH�B��ߑR�,V��V�%����jq�P8���\���H;>/L߯���nR7�Y"�.Ɗy�ܵᶛ��,0�P�,�Hp�����Z�ө4���	���\k⠂�j!�P�ؔg���`5���x��s�kl�6�ڊ5�v�V�y+ ,�;1��fl����8���0����,��w���N[{��}\����y\ސڢea�z6����a�\�1��g�r����y�C#G����-<T��kp�� �Qz�B	r��^�T�a(��)��ؽs��<��o?~���W	�۰�:_�#B�v깭5TJll!��
(�LJ��V����J!�S:�jE\��F^�U�T&e�>>�[%�\���Z�J�����t��?$�M��'�2�\C�J�m��N��U��3�RTB��'���颖+�5q*Rޠ.��P~�����׷�]*c��Q7y)I�`�L]\3�mnԱ�Zo4S��ձ ʘ��%�;:�Ŏm\���"�>�կ��v~�ŭ{�ؤ_Z+�j��S��b;���R���G���-�+3Ј�VH�✉��c�F7�@H�%쒇�%Uy���^�z3����eJ��*��3:l����a)W��r�3I ��B������5���Y�h�%J����@O��N�aK����.wB�vW����*\�v�bI��.�XK�[��&�~G�bN����<uVV%c\gkmS���� 0P*V�:d��ֺޙd�i����7��X��P7�A^��H�v+F!��!`#�h�����Q�S.�ػk����+�TQ
E�8=B1�f�e�.��h�<����(�YPJ�=�y�co�����������]DeA�]����L��>�����x���J_aV��F%������{�^c3^�b�(P��ǡ3M�&g��MK����M]��-^�A"&�`,�T9���u�K���;q�����p9Y���_ޠR�h���m������g�f�h���fuЈ;Q�|"F��zܺ�	�����]�Ѯk6T@Z�k����t��U���yr%���,k�.p����1����~�k��E�L��%���gw?�BF�#Q�f��Y:-e�˳H�Į/�`R����D}�0�m�0vvo�X���c_�v?�t*�
�Z��s���ț�}E������Rm)�t�=����`��j��HA��f�&��t�<G2{&�8�J'$;	�J!p��#��,�i����@��t�F���Z�Q�Y�U����B/�L�� �B������;�y=X�v�ƚ���	Ṳ	�Y�ï?=�|�F��S�3v�$�{�ai�$K��)G+V�U�5vOt��3ì/-�f;�+���&��Q�A���r��ɥ�LQud��� L�eJ�,�(]]��WX�s��{S����X����kE��U�Sp�Ή�F�/B�l���`�͢xpcu����%&vY�˿���yF�v�؈��]h1J�E^b���AnҎ$����"^s!���ZЌ�����A�@�V�`nR��*af8<�_�!�kbu�L��B6�p��[�Z�L%�]��	z,�w�z�JU�����u5y��NvI>1��`���R�w9�%�+�D5��������:�@�B�%�&j��j��^@@�"�
�F�����\͎m}<��8�rB?	���$�ΐ����۸zcU��2�6w}��FnA����`��0�)�.~Li�5�ڣʠم}p?}{N��m�f�͢M���[���Xp+�G����g:y�w+|~�<}=cj����Td�m<���ä�T^��~��|���\�t(n�(�jw�<��`��OH�5^x�yj�4swY^���*U�T5�q��+ْ�(�b��z�bw3O1��C�
�fJ������`�ǥ/Kh��n,�&�DZ�"M�S��_�v��Y��N��U�M&dl-l�'S��Ud�z�f#G[ȩ�{Q���~�v�ʠ%v��^����/�`v�a�z5? ���؋-��F����v��u�gop훏Hݿ���ܿAnuU�iA�to��ޏ�}�+�9h�Fm���l����l��1��F
�ݡ٨�X}>�+6��,���rV�zN��d^/T.�]�G�|N�Frhx��ܑ	&:�Z��ZX�l�����1،\�Nrq�>��w����E�Ē)���f�f�����g/�"�7*_�$s����cC�l���R�5(��]�Q��/�V7���Խo}r��b;�:�=�,���>m�E��C��+�L��VK���]�CF~�_~����=��\�����:�swN��x���B��*�և������
�:�ޛd�f�;�ƻ��x��~���=���G�bcD������C��I�ʟ�d��ET����&���4�V�U�tM��*�,.��#D�b���ko���&�X��[l�BIr�uN�<�J�H5U�c{x���(��o�:�\�b�D�a���.k���Rk��3��&s���E��%�����#��l�z�GsE�r>�u�#���&�t��Lj+����:���u�����7���gI,-2���(��u9���g�?���daӨU9�m-3���?x}��7��tiJ�yJ���ghb���+�%<2VZ����+��`�X,��%hm���o3}�w�<p��n��~ˣ�yUK���i�)�"��<�/2�+ �N�V���#��VL�]_&�k�6��Y݊+O�����d��_jDq)�6U�e�X�l�GU
��[�ŖVe���a��#ݲ�%Srɳ�In.M%���%�*p�I*8\>2�.�U��\
����]}H���`K��|&N{��Gv��S	�b�F�F>[Pʦ�a�!%� _]��͇�� M���JEA��-��A9�+:�4k�ܒ0�T)����Fy�� |����*s"��3�9xh��Syf痕�.`�b��M��强 �b�a����Oޡ�|	h0X�4->"��3x���?�?��W~��σ�*d˔.�]��WKh�R1�j�A��j�,*�I�zv���e�ڽ(h
�����D뺸���ܭ<����c�3�iSEV�M�|o��ؗ�n�nf�a�5H�d"������Z������[E�˧�M��n��jR͕IldI&2�lF:{"��vU�r�++Ir��� ��A����s��V��'M���3q���Z~3Z�%�XT��*��-�ٷ{;�.nLϳ����������[Yl.�˓S!_��O�qs���|W��{{�Z��w~��~CS�L ���VZ��g}pE�1{��"a�~����	���i�l���t�;�t�!k�r�	�H�����Z�7pȝ�i�����m�K}���:\Jm�x�>�Q�U�(�˚��x��w���c�Q���䊢�z)�[}�vQ�r.��"�+��])���J6���t�(�����]x�ƚ�����ͺ�����z�:}*�L�
���A`\v�o�K�-r��.9U���(Ca��!�29�Ǖ�wI�S���ڣ����D�NΜ�g3^F�V�F��V6Q&jY�FC��z�D�bui�Y����i7��_��3�s�L����A\)�tK�VE�Iru��,v�7��a�<�E%��fY�t;��`���l�d�j���h/7�}oAQ�bb�/SiPZ>//fq�T�j��b`!+E�B��)�U�Y=N�r���B�R���&�{���R��#1u�����2�W�{�	����2M��k�fTv[Kr��NUlF�ގ�9v����*�a?6���M<[��j�-�ϰ����[D ��-HdQ:��F��u������u��]&5r+D$��a�f�c��2�>��7B�b�*��t�)g�1����)v���ֻ���L��'q�����ˢG;�l�*n����.��Uj*�yW�d�/�*+�.)�-:�Ϫ�!����O12�g��7o�XY�R�X5#π����"? ���    IDAT�i硖���G����O#!F����:�����H�H�c�p8D6[���*:Y.���׹1����C\�AU��tv˓-/���mU�6�]�g�up�����+���^�ca�i�ǂ��^�~�Sӳ����QϾv�I޴ZUk�����/|�̷QZ����à��N����s�@�uk@�Ia�.�=s�j!ɾÜ:��g�8��%:���9l���A.:�*�j	��L�XP+�:�%Fi�U�\!�ЖzSp�F\�3�2��+������s��Z��W7XXρE|�B�l�-�&�)D��(j��X�����E���g�PO=������֖�RQa��%],8-'7������\}����W��/�./���r�l��7$ ��RZ�=^���i�}����%�ٍ/��zpq�j�O?;� 6����g�d���$jR��e��6ʩ-ݙ��W������~6W�I,.��G`|w��X�� d$"TQO��ױ[��ڂa�]P���� n�"�խy��:�G�%Sk��B&���ˀC?Q��-ʞ,r���\$d��7d�f�t�nSZ�`����[��ht��$(e�R�#O�d.E	� ����^=�PL�R��ѓ�"��u�n�=�l�8w�w�,�h����ZJ�����ϾgH��f��d[d����-eP���=Ӝ�X~���E2�e^�Γ�<"�4p����s/	0���C���R�W��Rl�%!1��G�"6ۇ�(g��~�Mr�s��������^������oxx�!�� ���X��Dv�v�AΞb1E������J��R�Y�1�Lp���J����a��U4�M�4��^����Hg��j�!CC���n��dk~SE2}��6����,�,PmX��$_2bt�����aSۢl�m�:~�����v�����ؤ�(���ĦJ+*1���R�s��u�\��l�k/?E[���J��z�,i�z�YN�:F9#�T��� 8�ܐy�D��E>��Ü�����į��B�d���:(�G�
dDrP���Z�P���x4�*��"�lMU��|����#����-���B�9��l�I�e`�|�܁��d�jl��� �6��R�nu�E� A?[B���l�����ZuĢw�EZ�R:�'�NS,K�C �q-U�8>�%�H	��E�*�R5�k/�m�h#K�,? �§�BOm6pJ��T����s�s'&���ެ�˔)����j[��pԇC��*���h���q:iڌ��f.�\e��5��t��l�(i?�@�d��yO9��҇&��&]����
�⋣�y�`��)�E�7k������D�T����f4�H���ʂ�Xb|p�2�!�?�-�廭a�Q�(�^"��;��ۍ����b%���Z�ڬ�y�m�7�g��i��l�i6��̲��R3���(��x\.r�VcH�@�٬Ћ=�G������!��|�Y:y�5��ԗ�����nq�q����KX,.IzS��шC�jr7��y��N���\�F\�Z��������p��27n�#�K�m�8c�#�АG�Kx���fp)@F "�2M�*���q&J���LJ�m��*�$c�읔JX\\a��#-j�aS�$�L�L~JהeL]j�%�T�1�ۇ�V㣷��?��bv���^*�����D��=
��[*J7���@x��=�4��SBj�\��u<k�@�Z�8@�NTO��AU܉��3P�;��d��-L��M�6��$�ky�E�(5Z��'����k0Q�����ņ-h%O4�dd������b!K1W �L���62D���(\R��)��qz��\����mU�p����VԌN�sʩ��tY �"(K'��H[6��*��F����޽%�7�&.+���������ge9�w����0(��QU��2��f	��qJ5+����my�J1��<'N%��w�\dm-��!��vhb�{ts,�*�y6�%��%$��X�4�"vR��*}�BO{��6;��ȹR�`�����x�b��W��xm�����$v����/&��
FQ�jyF�bJ�E&S�P���&�6�����3$�z"�7p{m�3�6�j���3X��l�6�=��+ô*�\ٮȠk�n�=�j�4��_������Ln�b�������J[{ΐ�R���X�@��?�Ã�k�nU �=��ĖZ��p�H�]�����X��Lz�:�V164(=^RZ��08q����}!��a�QQ{)�F5���� �Qn�$�3�J },{�(˖G{����HX�@�R�ꔗ]+��BE���)�rx=V����]�2kS��N{�J� �^J255C�f�#ho�!J�_��~k9�*�4A7�?��(�$ɭ������.�>���n�xKnC�B����JUk*$�o�����7�6���D5D���aP�+-��|�� �l�-r��V�������KϏ��[��{W��^�K���!�ƭ�I�ݘ�d���Xhx����l&E��[�&jVe�f.~BY�����uSctb�À��4�~UOE��?��*��2�����<8�Ե,��v�Ȥ�˓�t�lS{a�)�6&�j�n���@%_ցUI�F�P��J���8xp��.y����i���"NGQU��[�^���o ��z��%(]��Z�\�X����'�n7����\���h���GD�N잠�;��)����bRj�+���1�����׸��2���9j�S
5��H@����{F�����;|�����x|ڧ%/�}������Y��^>��'f/Y�HV� @����K���%��=��û,��Ӊox;��q��:�����9B~;��"�f�=;ٻk��ė���ʷ9t� ;&���YK65Kp��,�`X�v�����n���V˺<�d�\�/��E�A?�f�v�	[y���oR3�����{H$���6�bhr����u�58�9�h�x��m�F�
��Z��U��<39�]r[���νU~�����_b��=<��a��y<n�m���K�|1JM!7;��[�Ou����x�cJ@;-˪��T5�=�Q��䅥0�ʕ�}m^��2Z�R��y�
%����/��~�mB�������9������8������Յs<�7�>��Ć������0YeC]!��HW��c}?%�_��[��9t� {�P)÷Wg�9�E�,Y|�ֶ����쬮,1;�����.��B�]ߛ�K���o�E�=�ayi���yU��b;2�������*k�"�H'�l�B�N,֮yO9Zj�~�n-px� O��Y��(	�j)�+l%z�v�H��������a���x�`��Uh�o��͌���
r��#D5j�����_�;���R�-1�J�)�`�dbI��[b�{��t����`Ӱ�)����j�J���0�7��Jl�g���5��{�>�-�jg���ek�����]��,�%�e2EJ���:G�����[�\��V%fl|��G&Wfn~�T�����pk���e#�N�ͧ��}�Je�ʲ�I%_P�O��VB���#���ᖒr�ޟ,f�.!�5p��h�\��5�� �BE3c�Er���s[�����x�F��ǈ�a�?�F<C�&$m;.�+Y.\�fkq��&��=�Y��	�n�pc&A���e�~��[�QEEiU�)\�����L��
�����v�A�����7X^^��h�Rz�$�c��C`@6�l�3�aP>%A�Lb�TZ���KmYJ��`�-W��������8Bmc�4Ө��%W��o� #�f����"���G��\d�R�2׸7��-��=���u��X�����*K���d�t��V�x�6��hYZXcu=��V���.���^ZI��40[|3UB�VS)�B6w:5{.Q��8qxa��(�RafP��6B��.FYP]�v���oP,f9pp?�wn�\k���ܕV�e����ԡI�vaY��.���n�}Rēj1�UI�\���6:�|�w^][cs+�j�A�'�#�}��*UF"��2���F��P@F��0���B\���8�+6���Z��0h6��l�K,�w	e���b�{��R�LB������j+�Ԋ�I�$P���w6�b�
������%������*Q��{a5�CŢ�\)OVd���٫�RYnu\*���cN�Rf����Z4=�VO�����O�h�k8,VB^/V��13;�P���!�� v���D��Wn�*@� �_�JMTk�#wQŒ,V{qQi���N��!��{W/^������&�%��F�ڕ�R.�����~U[�`82D���aP
���n �&*��z>NWW�p����f�nվ���J Ś`���C(�M�����b^��V����x�`�t�52���=��X��5Uؚ��j��_�@��Q۩�u�-Hh�W���cm�ҩ=t���e֖3������
�8|`'����l�Jd
yV׳�~�>�J�EL����^�b��ߥo]kV[�Nu�{��;�L���:O��1��s����/���.T�����{�W�VBrs
6(W�"+6:q#��8;�#igk}���;,�\!�0��A
���͐ɐSoU�?E��L� 5���X/%�B2���8఑�HQ�K�dE��K�|����^�r9,f�ĺlh`u�/^*z�D��d��[]�F=���,��*����jѠ�?�K���o�L5�^��SE���*т*�go���|��
���l_J�3�!�	�����|��z�[3�Hœ��u��ц�!�����ͭ��~d��̠(���T�e$\/���3L����K�d�U�N�rF� Bk�����3H\��F�����ů/�.y�Jq�\v���c��~�3f.}AE����àتX&�{�P�v���4�0/J��y+���g7i�;�Ţ�/���J��Ϣ/!���zdJ���>6���{������U�;�m�,}����}��x\������Rl����2N��#�JB2}\�6*�2�F	�Š�=QX��M��~��a�SP��|����e������	�6S��oα�����NQ7�iz����7�q�z�L�1��Bu9�c���ۻfS u~��hosp�N�KW�YڌS��C�Ngw���}n����VaQi�p#3�\��;va*癹v��gޣ�X`��Af�N���X��Fv��چ�c�@�(Nw�\<���Fe���6�yr�l�3	����
���N{������b�����Ʀx}�1�𵃔�<w�+�7��ߵc;��P,[x�ïx�����|��#t�\���٩���e:{b�xjޠ�o.�p��-*Z#��o�,o��#�/g#ɟ�x/�Qy�PCM`,5��Ud	���v����cr�O>y�Çw����s��
o����%�àK����'K	]���5Q�%�.��?���¾]c8M�����o|KJ�,�%�{�t���I�I�P*��z%s.VQfk:XLP�nq��ߐY������?���?��N]���#\�^�j���A±!�V�_̓ϭ��=������3��wq��a^xa/���D2O0�����0����rd�8����7S����,-nj?��S�������ܘ����a��8?�Q?��\�v��髚O{�ŗ����������e�m��rzI糚Un�Y�TMr��v��!�LV��=���Uojf��j<�{�~���+�����gx��`$S5�ƻY�0
�]@p.y2$'Z����	��PmjC�����`���w�pnI�D�D*G!_Ft���+�F��s[N8�7R����Q��_��7�<�.��G��2�à�Ltd�L�E�dx�|�U���)���ns�g��d�xL�s�����S��7ɱ#c�+f='.����뤳e]:��}���|�k�n����.��;w�I$�LO�U����*�v���ܻ����k�۳�ѡ^��_��O<[��k��$9b��5��k��r
������R�iT�r+g�IK�+�
��W��W��8{n�f�������K�pu����4�^=��f(1
�C�O���4�&�I��U��G���;�2[��H�E"��$"AӠ6q�/B��X1�P{�IaQ=d�*0 -���� =�FQ%�e�a�Oph�����pE;�t�)U3�\�V�s��{Xy�믦I�R<��Ivnp��<��K�;���;$�u@;r��[5V�V�������]���=��R�KW�(���l���(����gf�L[G�]�wP(����5LFn��L����b�����*�z�$>W�'oW⩩��.�l��$�������j��kWXX�W�`r�$}�+M�M3��ﱸ��f�aP�I�;�J�i�l�ݪ"�y�J�W�ز0��vE����I�0�F.�SQ@k�=�R9��;t1 �/��s/�&��@��d��[���W5>�x�x<�2�a���>B�����a����>�*�7oH��
��tt��xI�
��.�LeZUip��{����Գ[T�H8�K�D6��y�t��.��2$�)XY�H.7_.����"� ȗ+M���b6���҅h6�Log��{G�� �nAid�*Z[>-1�_JԬɭ�w�.�k���;v��0�V������?[à]���H���c$��E��[�b��tٝϥ�,l��n)���X�� ��z5����#�eW�C>�?���a0y	����.�:�=T�f��sd����&�d�H�����F6�%+�e���ie u���m�߸<1��eT���U�
�M�^3����l���V���5U,*M;Cu�['~yE���t���e�8�����WO��P/V����Z�X)�%���;�؜n�n.r��"kI���ɑ��zY�8���Σ��ʽH�LyI� (�ʭz�*uY�h���H���������������Cn�yH��'S�jW�(����5
!�,��M��?,�k�)ݘ��:��*��K����aP�#�-�j�Qoʟ-�)4B��S������Q�����U �>�x_'c1-�|}��f�����Cs/����x���,&��É���鴒*H�xS�;<R��<�F��h���H�I*��V"E0�M��nӌ�dO�7o��ܑI2��"(�J��e�t����kG	{��qڃ͛���V(����-�f����g���œ�9�c�X�����7mQ�a����A��d�rO��Z��,+4�!�j�u-�>rh]�%6�ML_����>�� �������v�*VSɃ4q,$Z阱����U?�"����b�k�R��'��H�v���jUk�Ҡ���#�N+;���Y��]��ū���-�����z��wPnZ0Ì���f�FP���l�lX�bӵ�j(`�J]��N�M��l:E�����(D�*m?�d��T�D��=��uݠ6�9��J�X� �zw]����{���s�\��>e�&e��f�x�|v��ϝ����:������ST�.>:;�����r1)��(�!�)� 8b˓gS�R,[O���Ll�mA&Ɔ5�|g���[�<���vS LF���O>_UP�j��הWH't���ܙ���M51ώ�n�go�^YW���N��X"=�:�p�BX+���2��r�=;���~���3x\^���8q��O?��{����Gy�{O��g3���[���G?<���x����>{�D<�S'����9�����[�t��?������y������]<˶�觯��h��_�)�	���&�(y�IQ��u�`������m�Cb��
��Ǔ%R���J���;�|eZmv�vn��3�1���0Wn��Շ_Q��֬,�[o�V����Բm�?�06(fSZr���Nqd�������DB�xe��4��C1��8�6[�X�V��(�uy�
eN��j&��w�$�>��z���;~??��O�2}�[��{��D0zc�����S�K�ZA�i�}� ~������dcuM{������b���7�矑I�����r���71���^��	�>9���$���;���v���_}�H����\d���v����u�)�Í��{�=V�V8��s<��I>t$ĕ    IDAT��7��c��	�;u��Je	�B��'�wy����rpYqۚ\y�l��Ǥ�.�gk�Paf~I)t�h}!���D����YM	|����J� UM�ɂK����$�-���s��ꣻ���ߟ �h��9,�d�ؤ.���ć_���|�P���t\j(D�[àv��*�0�69��L�~����c�U��@]���d*� �;��t��E�Z]zGiW��������,�ͷ�ٌ'��ُ�#������w�36>�ԵM.\�R5W�1/�p������y�ܹ���^N�����h;/�9��%�?���n�IWW8}�4A��۶�wr'�\�:#�6�HՁܫ$(٧H�|=��V��'�3��Pr{Cr�U�0�J��T�x�.�097����:|�3I0 ?@��h�d����ܸ��b����Ü &�6*��5�)�ZHy�;�ur�%�+�{e���<�L�|>�����M
�2�N�5#�|�BYr�-ȅ�ԉc��+01$�`��ȅ�ަ�zS3ISH�f��X#��t�����i'�ُ�c'����\��������KLOߠ����_=I�c�/��ܙ���^���|��=f��x��QF=�ܙ������U���n_|�yBA}�5�l�'�=�@���G���s�����>�C���E2�*a_�T�ӫ�9I�W34*)�u��#��8����7�q"zԛ
8��x�B9����<�+j�e�ڍy�έ�M�nrR��!ɝ	QXM����2L�xR�e35��_�l2>�ǁ���-����g
e2ٲއ�&��$� �9�w'����b�� ʮɃ�wB�]Gl�7�/��s�,|��������%�6�\�>K�\���CTjf�R]f�H�{����+E�oy07C|C��&F��rg.��r\]��wm�����Z�����i�h�oh o�Ã�M,��^�4�)U�;�$�xL�
�Ԛ�{w��!9��'3
S"�����l�����YZ^!��ƶ��p�#�a!�m0u}�DV�2�۲oj��0�vQ)��dQ�R>�������V)��Y�$Z�R�gV���X�@柰���aЍ?�O��"��a4���ԟ� �q�h���>��,[뛜:���n}X.d�;��V��Y���&��9=`��0n��h�C<� Wjh_�l�ۣn����Vˊ��T���Ӫ�"K���գ��t21K�Y�U�B��k
G	9���g��LT2I\�m@�Y'Y�b��MX>��S�Ig�|��8ԧ9!ɬ���y�,��t2��æ����O�H�]�?��k�Vjh�._�j�3���rf'W��%_vb���A�uh��d3��u��$~`���ė�s���I.�`uv����>���A��kB$���Q��Q��N=�j�I���%l��ܱ݌�����������KO18ة+)H��[����Hg
��
��=9H2����%�67��,twF�������9݊x<V��\�s��2+KTvL�`x��d����[l%j��դ��r�V���e������B5��TH�R-���Jt�bv����]>>sAaF?T��!,5�G�O.qsq�����zW��4Qٛ��,VՆv�Ig�\䄖��l�q69rp�Gs��;1�*(��l�Rn�����y��.U����X(��jM�M������if.~AuE�A��)"��lX���0��y�_鼵F�Ju�&y�������q�<3���m��;�ѣ�XJ�Sfn�yč{ɔj,ҹS�玒�g�wg�եu�###�v(����)��K���qت�����ڬ�G�x�#���z�ͬ���M�,=dn����"Z�B9H�0��/�&&N�R�y�ND͒�G	��;��뛜�z]���N>����Wh�=|yy��i\�.UJ�&�6�dL�a�|1'���u�)�]s3�p�O/�Η�g+��)�k�������R�%��~A���`5k�+�L������͋_r���XJ������oȬ��;Ldd6�DDzT�\J%]Š!�M~�2������*��{����ٟ����˯��������e��|���8���#�u�������!�oع{�7fx��w�l��?�#fW�ݯ������^�Z�q��4'�?L�`��߽G:��g�׋�g�_$W6����H�ڲ7��A��j̕$��<Q��p$L0���x�i1I��]D#�k[�)|�.�$_\���r�v����*f/ٚ�է���[mTj��e[K�eP�uU؋�-%�vmܽr���.����Z(6�m�:��7�
(�rY��CB9\�ع}tPψ/�{���,�������>/?�鏹t�������@/��{p����P���Z�X���_�Kbu�_�����ѣ'��ONruz�����V�����'������Ӫp��-k^v��aΞ����FG���Ӌܸu��_}����y��+���,ǟ8��/�磏?W�����,-�p�2m]zb�߼s����q��qy�zQ;���ҡ�f�B>��X�-�����9���&�F}]형Y�KPAP�n7^����T(X1�!-��YLԱ:�If��kQC[��4
�R�z;�r	��Bj�!C��ꥳ
v8v�	�f��>+&�H�w>����U:{G5C��跆�Z��àT�0�8����z�]�~3���0x���z)��M���goh�A\�n�bZ�n�o
˜:4��#>��y�<?E,����>��G�}�g�}���n����YX����/�	=��h�I� 1��z����(���=�7�W�������.:��M|� ���'����y��1��|y�6K[y�f&���ѩdK)⮕�k+2��;楷=�t�[EI�K�fI��.�:�J<XX&���k���C��f�W��G_����&uQe�/��(J�s6��h���Z�rG.����0�\ ��H��n���˪d
E���'�np{n�jCrhBɶ�ﲐI+��4�0h�a�����0�MT`5�B�bC��ۃ1І-&�TL&�H$h���&u�z�wYXX�ر�<wj'ɕ����J�~�;/�=惏�XY����G��_~�V�}{vR�m��Q���^�������[�8q��6?�/_U�QO��f㤳i���7��v�|N��f�q���Qh�,F��$�����v;>�]��6����G(P��P�3�u0�4�+v�f�L��P����"��V��-�`UJ&3u��<��&F�� �
x��~/��\b��m��X_^��q��ߦ��%�e����7�A�*�{�jk��lj[�[���5q!=��AQv�m�X�A�����q4US�fl�έ���s�� ���e�d?�.�gq��۶���Ƶ�ܼqKc1cccl�akS@TE=X���9�nO=���3gn����S'�1����f���5�W�H$8<nvNN�4x�r�>�dQ������p��+Ze7M{��`_�����$1>��:(��b����ry.N]�\�����ٮ�p���F���k�)H���c"��܇�~�=��TJ��⎔�N��"p�w����������\^E����旳d
��������Y1�p{{t����WeP�\��]�w������͛�����'�����m�\���2F�_��b��?�gi6��������̩�4�N�����"�w�brg���%���e~~������M(f���묬��֨T��Rq�H���m^?x�$��o��(�|�L���̕�*@�r��������s'9��]�b����?��͇%<�^���y�}P���	U��\V#����bN���\ޠ^����i�Qi�[T'�^�<��n�a��W (�t����D��������`e�k�7�,\՞A�q%R	YL����}۟&�;�=�blPjȡ��ك�<��3ӳ\�v����ݵ��~|���_�����(�}�|y�>�.��j21���՗�u���:׮�ќKG[��O�S����?�0s�۷���釋����n�#�e��^&v����5>��2nO�;�H����mw9�&�MoXy�]t�Y�Z��(jO^2�Bg*U�-9WQ��}����O`�'�]�ں��?�̕�u�Hk��TUR�vE>���X.B���˿tm������!��º|���"��y��:���l�aAJe#'h��]�rI\>�����.,�27/�i)�Kwu�7�bA�{,���;�� 2
`�Yfm�O<���O�$�Ns��i>����W��
�B�˗o	�����;|;}�ã�j�⏟�?��"��n���"���12��g��se�2�P��_{��nX^�[7�r��-��<;vl��cܽ�ƻ�^��b�FH�����nR5Z!�e�����NWЈ�i�Q��e ��抬>��*��>z`7�=a6��TLN>�x��2�|1LF+e���\B�H��l)�R�*@�	ŽZ�������?~��A*%��V�-�h9O0ey���r�5�*��$E�0�,��J���DL��Z+q���\��x�9�O��翣$�1W���.�m#��������ލ<VvC���s��;���_����y�GF���?�ùo��ou=��w�}h��|x��ӷ�R�;�_��Nv�7�y�W^{�SOMR.��YR��'����W��?|���4���`t�O>�mmb;��_�_��Ż��K�n�k~Y�&�U#A}o�c�K�}U�t2Xy�����Q���������
R�H.�l���˷�����4l��E;15�4j�Vg��߱�[l=��ˢ�V��&?|�S��/�#/>}�W�s����_�RU�{d__���J�7��nY@�mR�,�نZ�[�`���Cnm�#��x����X~~��?���n��c�Űz�w�c�w�?�M����"�O��	�[)~��#n��W^~�]��y��o�_��3���LӻN��t���9�$$DR)*�F��NX���k].���.�S�[^�ښ��F�� �@��9w��'�c?����5�X�*���������9w�2�7�܋�P0��ϏS*YX\����WX?`����^���^�&}�=��0�uo��>���b�g�~�Ǐ��o�ן����G&��/�~{�O�8��u ��J<�����sz��q���
?��f��-J�l��d�̈́%�M�]�9��)��"��0�%�R�\g.^��n]�J�I`k"����n���|!n��k��<;��M�����ޢ5��7�}�L֨����Y�8��b�3�g��U2��7��W5�4�=-Ȝx�5�?��o�񃻵�Ol&��o#Y��%?�v�
���5(ĈbSj���}�]�,���y>��$�]���+���b����k�c�C8������h�[cc��}g/ׯ�q��9� �^�^�V?�����_��=|~+���I�f8{�3�24��������l3�P��37Y�JA��h��� 
��Z��}��r��D�m�fP�>����Es����W�������A���V�[�̻��ryd��ٯR��I�Ax�M�^'�-U�dK�zAj/y�Bj�F����m��ɳ�i�z���Rq҅�mFƓ?}�bŬ4u~Zm2k�f�X��L�Z�p���t3XY�T[Uڰ�Us�H�vڇw`�E0���B!��C��̡��lqq��e�عkýNz��wGٽ�az��^.���_�G�g��4�޻�﫫����6�V�t޻����fh�ڱ��� ���l�ƦF�7u��X^�1:>K<e��n"����I���nQ���?$�X���Dc9�A%;!���`���&"M!�v��ɳHS��'g�eMd�5%x��8��ɥzؼ�N��HN�0�JxM	�tR���|���qٷS����B[����Ըq�J���{��'�(H �xd%�K��k52���O4�g��D�&l�iC���U���NUr��a�^Nc�Zn���M��w�~��������k�=��.�޽˾��gw/�s��%#���һ.��;���h��}Q MN�c�~�����s�s<��ô�ۘ��b�Y��-�O�Q�I��V-^nݔ����Ef�{��J��~$�D!#�E�^#���"C�C�7���) I9�h��U�[s�i���2� ���J��B�H4�lEޫAVu���dI%L	��бM�Œ���X�<�E)�����vl�"(I�����{qF'�j�0=P2�i��	 ����S��V6��ک��:)��e#'�����w27~��ћ8F�x�Q���|��)������465�>']0��d9|h��5�0�T�s���������?�b���3�Ȭ�x��>v�hbyY�;w����?��W_����1]H�B-���2��j.g�+ܱ����j<��J$�[�+��桥S]��ޛ����=�7tV�얭�x�S\M�i�Q���r�6�2/�9��b���@_�T�u{!��֍�<��r�5R�8��
�����4.������X��X��E�P��JA$-i%�DzϺu,��2{�6˓�X��k�P���L���_*0��Y��0��n|-͔Lb0�P�$��s�gK����[\�p���6���mk��7?��c��у��ַ���S+=z\���A��ʣL�,k��⋸u�
��l�?:��ϧ9�Λtw�����r4���ϕ�\�vw��7��M�j���q�րzL���.�(�e� �u�����H�H{���צ�k)p��Hv���,ǹ~g�t�D���ގ�R��nL�����9�9�LI7�v����S>y1W���i�Wp;L$���4�x�k{ɯ�P�hoS(�T�.h�7�4��˷1�%��K�b�`��U��t&����v��"��}Ν��P���U�b���k�&:�s��U�jX�5���͗�aߞ ����ώi���G�f�Cü������G�-�Oy�O�Z��O��0�2"���ݑܸ>����?�.K+I^�\.7��΋��eV��a����T2��W��J����{(�;�wZ�C&F�\��[jYz�n��]-|n�f��S�J暀�X�.��F5n 
�sX��ײP%��/�M���QΠG%x^Eyw4r�(�h�E7 ��2�jQ�$\�ZI��_��ʜfi���`�XXI�q�+8=>>1��?����Aͣ�!���e-��<%��L1�dۆMXJ9��8ϗ����%�`��%=��Zi޲g� ��>��*�tj�6C�JVd9ͼ����=�`_?}�^����L��ԑ'���ͱ'��fj1F�b��!����,���䙓��n�����h��rp��nN�(�\4���io�!!�7.�\���t*50;��T7n�\McA4N�f�i�3��Eu�-Edcȍ�a��)�0�H�W�;��åф���'!�5f��\��ͩ�zPy٬���K^�T���u�|�u������Ϭ��g�?Dk����cx��f�5�y��Ӝ�|�o|���r�k��D���dU�r�K>[.��������ɭN���u���5k��_��3$Uf�ܭx�6��cۮ���b,/�ⴖؿ���������?4���d�߼�6�zzx��G4��s+��0B�j�\�1������+X���V6���ص{��s�,�b��0W\J����rif���$3����H����R� vw��A&�V|���I%��Hd��"y���4x��9��`h]��L~-GaM�N�%ߐ��h�3ݼ.Gӌ�-11S$�5ꆷ,u�En�朊��bv�9P��:�8%�0W*�-�0���＼U��>�F�#��-�������L���)��6�*Q,(B ���!��f0�2q�㣜{��=?��ŅI�^����i�������x#
��M"
qvw�o�:�WV9~�$�]>�������5�Dƹw.���g9w�eE��G�}���S���4��<����F�T�=��ƽ�x�v�I*���U���m	�x秙�Ze)+���ƅH\��O��<��%��I&�L��F%��[BC!��d������FZ�~C^rل���2g���%�:��X����\��Dxr�    IDAT�Z� �[p��"Dl�/�V�����DީuJJq\���G9��-2�5�<���ν�.߸L��H��g��c�M�E�"���0/PL��Y��\�7��Mu�+��l��`
��L���8����nk�h���<�R��� �݄W���f9g��|��)�|h5s�KW'�+2pi�k�Ct�F�It��u|n���������$�Z���Q�g����X�1<<D6�Ry�r,I����oWր���!��u��)+$�f�Kx�F|.��8��Nd�$&�j�d��H`�r���+�6��[ȕ�,,%H�
LϥH$�wd��#n�� %b�� S�:6�*5$L,��IŗY���ޝL�-k�{c��B�gg5���cG4��򻔂2�Qߧ��#�&B6��[N�z��������͠����x�{0{����Jg�Ă�6��m��'g�7v���A}�!f&�<sVL�ރ�����q���h<ώ��	��9y���@;�0�+�J������œ�ܵ���1�����b���B���5���K��j��I���oh�*q�"�����&��%����RTE�㡣�Q�s?��S��4^LjK�|��bCWo�WϠ��%�L5y'e9!JQʈ�P,fR�H���i!����a`צ.&n�"���s�V%O�F�_M賛]N1:�a�0�u���@�i��E3�p5c��0�츼>%��i�z��t�01���[���K�ɧ��ǟ����E���+l���Oq��DN�/�)z:|���86R1�9�*�D��_|���/y���I��G?Ќ��>���{������+$�kz��?�����`}�Z���"i��A2�J)z�|D�6�f�h́бL454���n*R�TIe�[��t�9ɮ-7�3;���Os�vw����tk5�4��K���`f��ȇ >��Ii���*=�~6�o$��@��OKs�T�LN$^$���gn)��$�/a�;��?Z��bjT_O/+�3L߹���u�W!��7��V7eB���tn8���s3e��|Y��i^:���;y�?�ŧ�~��C����A4��՟����	����9��6>�d�c�Nⴚ�2��}�!��{���c~� �`#7�\���ݲ����C_o�/^�W�t�/�|�)L*���NOWn-s��0z��5K���U�F�C1	��$�1a(D��\���r�*LW>��d2��Z
O�]i�n�Iɨ��T~���ݜ���S�[E6��ʆ�����)��V�6B��Q-�)dctwyt�F>z�-|6>�d�������l�����8{��6�����D�hVo�V!���q��k����Ϲs��S�.�B
qy�-���r��n���DnT��L���}���§���������7��-B>��ǿdbb��v���o=���<�w�B	<.#��/�p��U._�£�bx�U7|�D���!m�9�.N���W�0>��~�sڳ�=�z����R�+צ8{mRM�F{�JY�?�g԰z|���G)��/�Ԃ�3Y-5͑ C]�*�	Hм�JF|���dim�P�FG?yu�/���O�l��AE�!Ԓ�d��Z=�Z�:��\�AKe�����������A�Y�!�uæm̯�y�ؗ��MI6�N�bQ7a"��fP<��b�{���űױVhٙ�'@�*����߆��oG�n�nk�U�����
���d�ƀn���*�.������{��B~���/���H,�"_�'lg��q��4�.H�d+��ɹnϧ���L�,����sO`��8{�8�r�5�?C*[�P�3���l	�W�A�����d�WI'�&��;�w��:ikr�-���A����w���U �uJ*0;ei9��{�&��R�*FA�W$��LU~��(g���Q���,�O���f}�����+�\8u�����G�����7o]atj�+�Q/��Ye�_5�"g޾a��Z������d����cr8y��g�75A2Wbz>���F��^��ؼm�J�ePb��Y�"���:bq
y�o��˓g�����{ɖ��|I4US5���'���F?���@�c��biy���>J&�o�V�A�ߩ���~�<s����e��
�Y\^%](3�Sɶ�$�R>�N�%�BB�WV��#��w�sCA�X�+����U
�����0�d^)a%�e~9��j���Ybk9Jr߸�(�J�:%�L���֛A��ĳ,��B)MM��������=Ⱥ� �\�_���`����l��D�h���\��l�!��	aQ��G"2�t�u͍�������|�g�]5m����t��F�xZ��<���9�oK.@��vcs6N����-=��+�ڊ!o�¹K�NMq���	�x�1��Ў�D�xܤ3)�^��:�!�����4�Blٰ��ƙ��64�LJ���C]�����TX$��j0����v��ɇ-�L<WU
�z�ś% CM�S��.��2�4x	��]�YDnO���%C�.�Mc��6?łI���1�eF�d�>*f�f��i��}(w�����]���e�T�()S5����/~�8�����f2��V	4��_�'��F���/.Q�9�
k��P��&y��3���g>���Դ��t�6����t?���K ��k�d+�uK*����u47:p�%���A��G'���4�-��I	�$�ie��>}�R�d,���)�wfW���Y]��i��CC�k���@�NWG��J����ڝ%��ISeH�U�l�f�兔�%�h��ͭ�m�4	]Z
�lFbI���� ��J�&���J�D����*�=�N
Ei�5��OZ�E���ANғ��-!�Y��0*�M�<ux3��A�KK�hmo#���e���&W1��QHlV���G��c*������^狷�A�E�*a�0{�4�(�0�9�������6�d�����P_�tr�lf���&�%\:?���<��3���[7W5O�V1���hkm��u]^ _�����!��,�K�'�I.d�4Ghm%�(�tvu�sE�:O��L����fs%���lZ���4�$�J��͆"^�]�����p؋�)�l�8�� tg��T�Ē9&�ט[�Q�ٵU�4�_e
�Hn����"��uz�vR��n3�����[ZѨ	����J��{�l�@,���S3:�Y�bk����X����A�_e�O#�؝n�R
���w���E.����<�������E~�m:�[x����P��_|H�TOJ8��~�#.^��Ou��̳/���(�X�-�OM��ǧ)f�|�;���q�ӟ��Ġ��i쳽���5����K3�9�K���4��*k�Z.���"��)YS8�����ǎ�a�v#n�w%��Q"�!���aXbeo|r�s�k8��d�e_���:��f�AP���1�$�hTB��"twz�t��f\����3ܸy��N����\!��a��U�-~	9�5ZB>�J��B� х9&�\fi�щ�u�hY([i=TCc��㌬���BQ�U��J�C{9�o�;W�p������������]��8����ܹ���;����;3��nz�<z�������ٸy+뇇����JE��"���"�i��z��p���;�hon��[�DL��}��5i�5���tkV��#�|;���K��"�k��My�"��L�C�km��5�C�(�2Fa?����"�|��_.��I���t�C�V��j'���6�"��Ͱ�o�4�&�����6N}|����РfV^8;�ɓgy��S�]!^{�C���5+�M�[�6B躲(1���`3(��O)̌@nI7F2�Y�X�7б� ����͠HNeÛ�c����{����iΝ<C_o��x�ə$����:�ܻk.�����ܥ}�%���'��K����*�qx---��'��p��ư�\�m[O�d�Ϗ�c��m>,6#��0=�b	S6�1X}��P	���í����JI,e��EE�I��5Dg[��!�QER��$�D�2V�n�<63�|��h�//���JJ��[u��M�e�f�*!��A�&U�[��X�I��O�&67���C�x�f�f3�;���>L� |t
������咵Z�Hf�x��E�ܹy��D��Z���޿{]��B�o�����C�c��M6���vb��X��Ҩ�t��&2��nN)HD �C$��T��O0�2�j!�3�70��AV�p\v�'�tJ�=>�<��E�B��;6rpgs��|��Q^x�Y��j���8m�bI���9DU(����d�e�h֫�d(e.�xz�n��z0I�_�O�l�dS ���D��r��J�����gy!�f�T&���W��O2'ߪDU�HQ���*��A��
��</`#3��y��<��tw���r��m=�y�}�"Ň?��J\d�r����6��K>��\c��A������	m����1�=��g��Tl��|MD�w�o���tV�&Lb�Ũ�c���C*Wmb-�J,���V)�R|�C�N"=r9m���x��!�	g&ikngx(��t�d^�N/�8K*V���o�%��q��O�[|��a~!��mA~�׸36���]((�B�6R.�(��E�����XO��kE�٘n��c����P�}:gd9�`fu��S����Ier���	R�������g9�b�{�i�fP�R�
tL�<񭉼ѧ��<��"ƚ���h�Y�eI��D����h�qwJ��y
%n����O�H��^$�n:���=^��=���S���=����).K3���j�"g�kc�9�_���$�Pvg�L5��kd��n"�a%�N�[a�ޤF�D��XJ$�Z\�f�`�z�x�]��9�S��$�PJɬ�a(�h
�Y��p;J<[b5�D(���g6P.8��y:;��2dyN��k.�[ kt�(��Y
N�S ٘D5$g[1Ʀ�ڛ�����`�oH"��Uv��P(Y^�R�Ԉ�$�Y\bfy���M4��A��V�PJQ3�t�!Q�ȀN�_rW�L\R�&me�-D�VlF�n����m��Gk�w�����O?�J�l���d�ƪ��̔2��7�u��[Ԗ�4�G�A�,U^<mi؃�y k0�#h��(ᰉʤ@6QW�T�)��h�dJ;������o����L21�,�=]���ɩ瘝��S��|�2�P��M����Ss<�w�7���+\�t�}�v��fn�L���d7�މ�$2�
�;/�q��4%�I��4;�v3��Dr�k�t��3�����&���"�T���+�,��P1�ȗ�8�!�6�B��杖�
�f[�=$�2��а$ݮ+��*E�:������)d���Mc2Y��K�)����ɗN$|��dQ�@�Q�c���f𣣯�4���?���:�� OO @8��i�QJ-��5����=H$��M���*�N_�!���1Y�\�2NL�.��$�s]W;�]�֪FX%�*���=��-��"�ʪ�g�p�6��-t{\�X
�Z6��b4����>!�&��A��ɻZ)�pXj�j
�{͚�춂WV��4)�9E!#�BՊ4y5
���y�+	W�$���b�x�>�HL�,�U�+�!ynF�SH_&w�ԓ$��ab����6��4�2�K,���CKW����\�T��E ��z3(kL��	���fo�G�Z��0���N�a����=��E���	�<G��MkG��WV���y->�n
9�8����k,�Ma��Y�q����-rcd��*U�#�������6��XV��&W(��n}�롌���͠H�*X%װ�]Ka('h�:X�Պ����p0;��H�D�b�xp�}*��IvNU��4s�2gnO2�bt�U.�u�j}(YH�fPf-�d�,�U���I'gټ��'����q��,��XNN�>E�j`ö��.�r��F�6U	��1J�Y�6���`�zbKsL�\dq��� =��fć%��C���-O����kn#/�|�r)�a����Pw3�rZ���B������
���+8�F��9��%
U����e��C���$�j"Gt5�yh�t�ٹ�Ss45����H8�b��A�k	�����Ѯ҄r9O����v�$�U���0j �,�j)�!���-�˔�n���ވ�-�'/�GM�%���.���h�Ky����.%��Oq�L��CXt����?H}E��UC!������\"2U]Y���#�+/��\�L,ɭw�Jvd�QC����Y�y����>��œ%hu�����2�f�m���p��g�^x�f��Z���n������M�R�z��B�x��}�����Ko��\����������o�;��}�V.^N��H��Rh-���d��^2��W��2����\�Y�P��R�@2�R ���Ϟ=I_'�jL##�$���L�CI�^A�T��N�L�M��!.A�;���*�w4��&�^�f��m/�t2k�)��*I�"�R(2>9�B����
U�K� ��~�M�Ƽ�L�r��ƷZG��].K�����FX�r�
�K�&�����%}�M�&-�TJa�j7��dǦ-��]?��As~Y���{7�K��M���J輳���A1�UB��iS�w2��� ���BY�{�N̦���h���o&�+P��h���|���K�O��᱇�����nr������?!V2�7?��f����5������_(�R|��/�y�f~�ڛ<����|�����W<�R��8����$\s)�ӻ��g}+�TN4]��&|�n�䜹7[cjy���)��I'V�#r���ަ�.�*��W�8���Ɓ���Ai�!��V`?k�dD�f�h�n��H$ִ���v�j�藚���t�@#I�
a��B�A�Q=r����ߐ]�������V/����ZL/�XC��7�nh�����A�:WK9���X��Jee�%^H�+�Q'�JZ�PCN1N�\$V�طs�}�����c���?�����ɏ���%���_���ᵷop��-yxG����?}��?<ƞݻ��w��ѱ	�߸�/=��[+|~�
6ODQ2e��T�<G�lt����;�K�@nm�ӌ�)�?�B��
���3�,����e�<���������7Y�p��*��f����@S�A�C}E�Ng�X,F�U3���z�:����b\�@=�6��X��R�K6U^��z���DK�3Y����4t�'�������͟i3( ��^�������J����j�sx7��v\� �:�[M��p��t�X)'�8M*��$Di���!�ͱ�Hb�	46R����G�؊�b��_���H���/2re�[�n�c�!�+o�w�J���O?D�:'o��!׮^揿�]�;�6���!r���ĊV
f/5����Q 22���y��V���(��T���V��Y�&�ʝ��*�wzb��RJ	�[L��:I�$�Я�uhU�3%���0�em��J�<	�G6��]��X+�O�i�S(&��2;?C�P/��]GŢ��'1���d�-��L�c1SHeX����f���w�.�a&��`�"4N/�M�����l��`u	�-��n�*Y���'�/WE[�-ԦY��Ŗ���p���Hē�lزq���[9��9��'y�٧��=u�/D�@;_���<�[��}}�S�]f��u�z�q�mi������EWo#Ǿ�`v9�И�HV��O����nZS��P���Z
��e�x�d -��RU�TK	r��tV3L�llm���`���'�Lͭbw�VE�WτTp�ԭfYa!Hw/O�"�p�(�d4��b�,q�݂�l�f�\�j��M�ҸK$��Xe�%SI��L��|����A�=X�{h܆�}�W6���qa7�0��X*I\�2>�	��I.�cq)J:Q���� ��d-�����(��-��a4���V	[T�%C��:�ܺ5Ob%F[S���[^��ūtww�cg�YFJ�}��b���z2�b1�5�HjrS���\�%6������$�Oʸ����|���)����HWW�D�9��*'%j+/�^D9�����N�.�Jie?X�J#n������PLL�A�%�./��Ҽxcn�����1>���$��z���fPknC	����24��    IDATfЇ���0��CX���~�	H�BK����7h���������ttt�g�V2�,�����J�ӯ!�K���A�Ϥa�.�W�j�����e�ܻ���'�NR,y�ǱX\�z�p8@c��h<���h���T�AvB)�['
�\,�(AW���tD�4�\�.J��2�I������.�Hd�$�y�f�^X&^4����̲ͩ�%�ՆI�U9�n�=�(�h���P�Ba3�m;^���#��ܼJK�Ek[m�~��f���e�W�
9��\�ɒT&�2��T3�7�����+̏]ee�"df��3V�P�kS��A<�����ԇ�����L�X�-���$"�ύ�4�-,�s,E�T�$�����шM�F:5����a���m���3���bueYM�����8}z�DBBtWؿw�����1.]�ȋ_Ne^�x}AF�׸t *@տ}LB��+�;'�y����u�p�8��&:#VL��$�)q�N,���D�D�B"���|�x>���"s3sd)�E3ec�p'�LNu���A���!�ue�z�D?.�M��M2���Vf����^&�|����̲g�������9�8{Q!&�[�J�\�W�i�z�f_g3�R���3v�c����i�p�d�jrbj�D疃4�۪���$�A�+"C	��4�{��5N�;G�����vkd��%�b�`q�XY�a�p{wⰯ*�L���zJ��/�`vaU'�6�o� 7oNp��<��S��42r�.-�,E����Em���K��U*��N���Z����u�@y��H�h!'�|�ՄOHu���ŵ<K��d����c��!m��_�uD�Ro��l���(�OC�E,�LI7I�Z�F�������&F���ֽ�o���=�47���t�+7��Щ���귐	���~��*g������BS����1Q�,1�a;��>���1Y�xD&�]�f,���@{���D�${ʢq��i��;,6/�<ܙ������k5�����ܦ*gN}IW['�����Jhl��J�w>>A�d�/~��+�w�JDyh�>������;�<�"m]���W���1`v5hCPUٽ:
���pk!�s�6ph{;y��f��l��I�ݺ�l4���k�2Q~�J�UZ�^�Z{hm颱��ݹ�}q�՜A��f��J��yL6��?��?���D��������b��?Z�ʦ��R('bQ=3�_U��D6TE�<(a��e3x�_�]��=����FÖX0�<����\V	���Am]4�v)<�,Y]�$�aZ��j)���W��bwy��J��Y��o���'.i��M�8���g��g��}}�ڶ��B<WhK�f���}��BA=��>�������M��V~��X�e���̩s��W%�1-e"'���,���Y�����V�9�"H��5|���1Ʀ����G8����8ini 
��ނ�렻�C�l�����~w�p{�ߧ�ڄ�T�m����"F�A)*��>��r�D!���4c0	,�#r:�Kbg
:�1��,ż�($��:�R�	K3�ɿB��mO��s��J3(2Qim� �C5�1z��؎���?�g��f�R��6��\ȭR���3,c�ن�T�h�F�����lnq^�$2���7�Q>�;�����v����1yo�뗮�7�����;�U��s��e��o�A:���矡%��c�ؿw?O��qr� eGX���qT�V-RN.c)�y��V��<L�N�5 [6S�yb���tv!��R�BN�f�e%(Q!� M]!�F.\���H�e	`2IĀ~��$��-����65���+*�m�JM�����Ȧ%��A��b�,N�*� �b��yqHa[��4�e��?~��`M�A����L����� ��C Tq�v}��A5��Y$�Fhp92&wO�h ��+�g��U���wl����l�F&��"���uN�.�Mihd��><NaA�������,'>=Ok�:͗<{c��h��'������5�@�D)#���1�R���*�I[XH�ݷ�Hk6w2���p�	aԏ��565_Q��w�4�^@5U�C�H��ԗ��3�$�^,S2<��Р\���Y�UP���`�����k��т�h�q�_'��/2Q�J6�W2�z3(p"/��u���'�A�lC�n�<f��H��V,:R�~�d����R�J2�Ռg�x��Y��\u�g�7�q��U�\�g�g]3���-��<��߽F2g������|�:�Νe����ܵ��Fq�Z8qzT�s�۫�m�٫ߏxK%�f*b3�عa�|CY��N�y��,��X�&H��c2��)K����,p��R�5��JT��:L����aQ7�� �d��\��R����y ��:|z�ș!Tiy'�N�=��֤��W͠��W͠��YͶv��p�z���^,gu�2�ي�ZS����&\n�b��^�EI�-���������*R����R�Dj-��ߠ������N$ؼi������\a��-l��ǝ�1"-��0��q�F��P���s��y1���^����S���n�X�=�Fd�5i<Lf\J2��L3�czY��)�qr�&����F���f�P�I.���L�eԦM��u�A�3��Q)�Պt��tu�i�T�=2r�Rj���v1���D��g'�T�-M����$_�(��Er9�ƚ\Ojy��[���w��K���PMb�%�⬚�:y"�C�Fi{񷭣j��e,�5��.������eш��k��|���e����ϧ	�K��ۏ0=6ͥs��\����w16z���i�y��7��oߤ����|�y0e��[��G���#�.+��\f��]��'y���T�~L�3K3P(�t9V!��45z����:�V���+���Uo�rer�,�+I��V�K�V�[[�\�����v���*��zt�4��JԌ���%kN�;��b>��O�A��9�s�[Ȓ�lF�HK�p���S�K��c��`	}Jb�@�(��z jog3�b��?���O�����H�l��!��Mtm=HK��6=��*;��"kk1�n�n�mV�<�p"��%�ժ��ɯ���b��ґ]TsQ�}�m�a?�ᷘ[�r���y�֒^��������\���gmm�?���m������T�̏�;���l��iDA�r���`�������NtfZ#2������sU�%&Ƨ��f�Z�ɨшGQih�&_��KP����+DVǮnT%������X�h��4�eR�U�t�	_>	��aX�:�S`C3�lA5W�WM�I2M��R)� 2�?yg5� ����e����;�G� ��A��v7V��D���ݛ8t�UG��\����l��]������V��-8z�$�Z���P��cmc����L��{D�~U/�*F>�p���$f��P���][�3���"�Ϟ��Ͽ��o�B���?����'S��HZ�<5`V�Y�R��5���G����b����v�����|��i�b9�E�@���m�^Z�V"Nag �Å-h��x�7�}�Zł��Z�P��]�h�*�aY��_&��fPTi}^"%5��{�����ph�v�,H�Lq��[�e�l��[6ۂU��ඍC�c+{�W���9�g���������aziAñ'g�
�i�A�e�P���*�,C���d�� V��E�V�t"dv��t�5n��Ƙ�Z�s�m�*D���j�q���LMMj��������kX��=O�����C��n�Ƹx�,g�]��o��3/r��<��c`��)�v��8�|�Ì͒'�g���KO��#��ȝ<���~����)��444���Dw{3-��~+.�Ie�6�Q��o�(�e���d�B5M+�O��JIr#]J�.i<��d6����)d	�]h�E�B�5Z��Czo�J�j��DM6�q�Wԋ#��|�"���㫜��H�&����ϙ������ d�z)X�|tl�l��fРt�Ja�����7��@w@<��>��I"�������%�]��$�Lj����Po�!��d�X���U)�����j�~C7�۰Y�
F�Z|ܻ6�1#�X#Q^;v������dl" K|���a)��4�3"2_Ȥ�x�F���+����$SB�6	E�hn'�w��[��-�#f���G/`u�����4�r��,6����1xP�h;Q��x%sWďVR�K���-U:�������Ă8\z��d@��`(�4��|�>�>=Jm�>&*/�'���-��2&O �߅�!�6m"vmd��0+�iR�����6�F��S9r��紓.��}o��h
��K��V�rSĂ�e����#���t���Z+s�ڨ�;�Vm�#v���y&��)f+��l����K�XM�1�L��N2y)�Eh+gk��A�qvoZ�`��ܚ��B�5p��Wn�%U,��N�/���DBn|'B��������x=���wq�"��.�r
	V���%�C�������P�U%�BT|"��S<�"�1��}D� �rQB%����CXɉ�P��-����6�f/�|؛��>��2Qw��Z�y���A�4��+�!�O��?�R�|.[��� qb"��Ĕn�;�ٲ����i��o�8L0�cqv�å��s���=�{[�e�X^XPօ䳞9w(Hw� �n̲M� �*�eu���k
�lF��ٳ����rz�Ʉ��aaa���%�_��O��˯�Z�����B>�2#���~�\Ti��N�-Q�Jp�Y��u0�4�r~�3(��fќl�>K��L��lW��j�
ޓ��?n-�2GC�鿬UL>L��z��fme�c��dKd�%<jϳ���!����*e	����H>��ɤ�<vp;�x�'�@bu����?�p�����={��/�O~r���*���wtR��W_gz�>O=������c�X�q�zf~���c����V�kq��`1�L����6���&��+��b�Pǖѭ3����|�Ʌ�B}��A/���F�!�d�Jf�ō�h�l3ɖIa=�Nh��[�a�Z��P��d21��MUpX|��|��XU8����ï�L�~�.	U EE��<�ܚR�֓\Ybu��w�՛��,&��I*�T�����7�L�_k%�U/5*9��"�jK-O�/�ٲn�d�.�g��.V�AL��YZ�j3���?8ȝ����N����ޔ�>���^}����瞤P����>Ҽ�_x�t��[o��K��>�$����Jr�8"!M��!��L2+^~�a:�V⋳�|� �T�J4�&��`na���(��9��C$Z%���w�f��2WG氺�����DT|�����ʇ��%���W"�}(�u�"�1;]v�N�	��l�(�1�:E2lUͿ��DrS,Qy�S���C>͝K�3~��?4�&�,2r`h�@׶����f���N��f�T�i�.;Ns���q�A��æ[M-����K���c����ӛIE����Q������_d\ho�nr��3��'x���F�|�1��W/�P���-[�y���ӟ��s/aqE���R60;D�_�`��P��B���k(���[X��S)��h��f3%n�N���QZK1?;O����`�p���������\���SרY\X�}��t��ř�,�L�J3d�+�M=	9Q��Q��26�5�invF���H#�b����dKČ����P}[Z+�!k�[t�'�`1�d농X�9&o]�\S�5��q���\.��\7�5І��*�����
Aٽ-�훫�^���:�<_�����_��l�y�	>}���>9���E3A1�")J�-y�a�[;��5���e���e{g�c�z�Y[�LI�f	$�����ܓs����}!Q3�Q�b�����}��O@@���h�]t��d��f^e���B>��ζ�L*���b��Ӹ����������t6��y�i��z�œ��V�>�*�W6�����ƽ��nf�?=���O��W�B<���C��4t��q�,�H'����<3�6*�L�;}����G�!�,a�j�$�ry��ɞ�PFy�>��`(���J�N[ �-��f�-��Q�C&�_v�M.��
�`p =��������X��w�;���ٿ����7^�������ц�D0u�dG#�,ʞ���)���ˏ�ܼ�˿��n�#�, X�s�O�,j��};��4Q�'F1lo����X�/���~]
�3�N��|J\������f�`��%4��c�@A���16u�s#���*�w�b8�b�K��FjMR2�0�]L�u�᫏!�6B]��/?�Ds�	L��b2C>�2��kJS�k�P� ����qca��:��ް���_��������#�S�������@,�i��ɉئ�~ؑ�IPc�b�żHNΙ3H�z}Ld�K���/�ћ#�������h4�C �ǐ��QL9�Tj�DN�y:��[͇�����dF�.�*4D�n�rF��������Ciz�0=�Ѽ.m`��������8=���6�i��09��C��B�R�v����/��dn�>��Ƞ�D��v�N����-$H=l7%n���xcEݮ%M�p4�����'W	���幞<>�l"�l��*��m�n�t����נEG��65�RWB��r�hy����^�l�U&�[<<A��˱��A*Es�
�#'5�F�#J0��y�74�������&�]j~$]M	��`��c0
SƳ���0"*�nc�<���R���=a�*Q7�p\�({�p<.fS}˟��"at[U�Z��ӈ�C⇑�%���1�"���[�s2T엗�m$RA� ;v�R�R�z_ܩ��!	kPJ�ؠ�=(l��+�ȧNO�f�Seᮉo���V���Z/ ё�b�E�fgȦ���z W�m�ڭ��,Ȗ#0��0��Ո&S�V�'����mt�J@���w֪�Ep��+���W�.�OE}(�WEr���/�AYwf�&.�b��cHO�h�n��8�Q}L�&p�h	��5@y'�tG�����e����=,>XS��N�q�M��]����DadD�DV7+�3�=�`j��ÇҒ'<�zX٨au}��Q�M½��3h��Q���0���74-���,<��q$�7�3b�{g	w��Cj�h3��rO��g�4���Z� _��@�>�X2,N��߃��S҇��cQ�=ʆ8�{�m���kdN�[�`W�]�d1�A���kI������B�~��z�������s4�`����F*�#��`4ED�ʆ�
@�#_'�7�,D�p�k;��y����c%,޻/�EO>~��<X���m�͟��n��'Ο��ϟ���=��N�KX�O�6f�N��������k�D�J��$ص��l �w�;��b\�AY8���۸�ZF�;�1q��g�h<�l>�T*�b��b)�`4���n����,]�d~t ��)�����sah8A0(]��uh�FD7�xC}<EĒ7/ ��N�a
x �pL��"1�����*(߻���_��|�� @͠�k.	%�@񸸉&Ǝ"������u��M��cb��đL�����/�����o����h6�HET���<f�~�΍�ݪ�ei�ā�߿�����A<v�$ΟG�^��*�խ��r�S��?������7�!/@U^0*4M��k��X�".��w��L^G��@��Y���q�����3ٽ�Q(�"�N#�K �ӑ�l4-�ؗ?��w>��P�h�|����羨�kK��}���p0�űD����Yvk�E���\~�1V8�U�JL��q�9B��675*`�޵����e6�
M����S����c��(͝��h����졐���'N���cЩbl�����=FX�[֣w*���C�:�LΟ8;��'A00�������Q1x�t�:�.,#�I��̩�)�>��߭���[���+x�� ��ĥo��8�5Zts�(�?��P����x�	���� 0�>�� ����X�fs�҅��,&�G��.a�-�Q ��e\�l02bB�	�����x    IDAT�����v�����'+YK@~ ` ���j4�L���h�:}vWy��J�X��x���,V"� �N'�E�����/���7�����pKL`$�c�Dq���G��	��:V[܆_{�<�x�^^Ļ�xZ���Q��l�=6$H^�X	݀��� �ڃ�,#1p��i<v�(2i��F��aa�Ƶ;����t�פ ���ٓ�PÈ�be}w����,�����L���%d0R�L��:���4�:7��rYe���6����	��)�����S�h5��`ċ�������Pi;%rr�1���C�'� E�t 	�(iҥ�,��"b�A!�f�p�I#�BP�����T�� �)���%?4H�iQ!�揣�(�?�k�?x��˟�_B�{��^�����Vm;
-ss�Oal|N.�^��^g/?w��������{ТI�Ri1���j��=��FE�Tю��o!s�Z5qh}��0|T2Z}[��+�I����@O��1|ǎ�$mO��v�n-�e�*a�蜪��t�I�|XŰ[�l2�?~�id�z��%��.3�"�!����6[0T�/E�=݀V�s���">���XanP�'��g9�7C����X�T��!�)A�K��bD��c��V"�u4�P=�R���h��j~�	�ҳsl�ygt�(��82���������� �z�vvVp�Ɨ�$r�|j�R'��F2UD"��{/���*f'�������F�����ijy*',��f�B<�E*��s��+J ���8P{ǔq��Q�T�t��.~��gТQ�C��m�0����v|ɰ�CS)T.zM[G��0��"�e��&�t?o@�{���_�H^A�ن�zhn޾��K+��;��CS���$��>l��k*����c�H�qo��7yz�$Y�����*����`�wVg��F�Kd���Y�j���|��V�/������5�h:F�]����A�����w~
ow�ӀG�6#)�ⓧ0r���$�d�la:w�t ]��<���:~���B�����W�ڤ\*:#�4�!�s��z�+���lBLhRq��Ǥ~l����
�ךh�S�9M��*��Q�T�d�z;��:v��/�2>I�dIɇ�"���`���1�1ЫU���D�o
;��C���m��0͎4�ɢ�f٦]PH�g����Wa$K�.q'<�8UrX�Ѕ���鈱T�`�ȊS>�z�.��l�W	��,��þ��f�2q:H�-t�#�d��,~�[2ei0jB����HO0#M4�@<������#�8}<�F����5q�&x␉���=�	QB�h��� M��	&�p�4
s���P�� :n���y2MƱ]aqEyϳ���(����1z�l�B1I{��pQ���� ��p���x��Qܿ�$��t��f�$i�i2�txRI�D6U����y�!C�ƙ��d��T�S[��x�X��V��3Ǖd���y�u�R�B�=ےK��8�K��?�h� � %*6��%�������h&=��8�8zt�O`4e��e�:nI���{s����KXY���h)�s�&1=�D:a���/��)��r'Ӹ����w��$,�����q>4�p$���M��zw�<��SObn�8.��;9�wU}�j4���U��x]���1��l�ET�.�G_\�/>���E2E6�@>�D1�F&�D<A,��f������ǵ����0�!���PB����I��\0ME�B'/M(Lt�!đ-?�t<N7XD���\�2�%﷏d:�b!�~��݅���p�՛@g�������62��c�Bfz�dУ�+�.�������bg����]����x�*�Fm�jR,����Z�9Bs�����an:�Z���;�P,&1>3�`{q�;=4�mDt��L	����[�-�nl _��O`u����2�9%��� ���?woЄ�vP�y���}�Q��R"�=E?�~�B�b	qfM���� ����fƄ�~~�._�c�4,�/*dE��w1}w4_?�?�Y�t>��n��!�P�N���F%����Pxp�YA:�B�n��3�+`P5Mܻ����Il�X#A��(L��ԙo!?=/TeZ�C����sc���=& �R.���l�@��C�C�9D}��5,=�e���!`j*��S9�sr���3a��x������*}�6����麅�����q=rD.�O�\�Cb-.Ih��u��"���ū��c�joV�݊ �Ͽ�_�F؈���4��J����P5^Ҟd��b11q���e���"�#,�*
�y>q���&��tf�����Z��ٰ�z;�%	�Baq94emU+;C(�.��&�̖��
��qq��!���姸s��
��������'�?znl���M��{�5Qݼ�o?w���zm�և��pO�t�e��E�]��Hŋ�T*��di=u��w	d��>��6vwv����Z����	����b.��)4%LNe����o�ރX��D�3���$����Q"@'>'K�	�ꠂ�]��S��0�����7�XP��i-U��|T,�Ր'3�(в]l�=\����w�e�_$	�Zư8�r�T��+����B��ƣ1�S}���ވ4���Z�z�!��HL2���"�8Z�:��-]�v�-������y�'����O������6^z�U�1$�E�\XA�F~�U�NJFc(���"ڲ7^�?�_��et��
O���եY��<Qبa�jӂ�n ���WÑ�a�4g0x����7�0jƃ�L	goo����eD��n9�\�@�^�h��Z����C��%o��/G�[�<�L�^c�E�޷/ g �jY2���Mv�cqa�p�:xH2�^��c�LjnX�i���L"�>�AA�4L�դ"��r��딈����$W���C3'�U�0�|��I���O](Rȳx��.�V�iGT����hS��ݟ��_�Ԡ��^}��6�\��p��l-�H�0Js'�.�I���u8�³jH%��?~Z�'��?��hڍH�z`$�����o�0��4jJ!O�17=&1.#�tv���Ɗ�h6+�:��2�,c$�x>������"���X_[E��ai��o�c銬��5��x�4������S���鶡3) 1��,�d�����0�Մ�`D'T������~�.��r�q�ԂY��EN�8���~M�z����EZBN�y��q+��]�R�"���	�Vl? ��)�m̎O��������o��, ���{���Slb�G�85�G���d�!�7��>�S�5�wi�+���0`(P4J�Bzԟ�i� ϶Щ7172��?��,0�h��X�X�Ça�@1axpZOӬdG&bht<�<|���-ԪMѾ����$=*z=��lؖ���{�uDs���i��6�uZ ��>�v�뮮�^���c�h�i|������;<Xمj��;�M5 Mz0�y�z�\G�.��O�n�>/Cǒ��ʅC�	�$E��֖|(ו�]:�r����p!��h"�w��o������aͯ��-�Š��1v�<�l�&
�����3�.j{����x��<V����O�Ca�' 3)~����t���ҁg��`azj�c)�2�+���p��f��S��:�}LONbt<����,fjv���X^mJôk2���E����Ҽ�+~/<{
��*�b�t��Q��EsɻBh��U��>w�{l���Uٸ��N�,?�5���]Ȩ%ߨ����:�+�bj�9�Tp貞�?p�)Vf<������>��쥜- �#=F�u�E0��yzr��L!C�>�6Ο?�g&q��{h�Z�\W����plMn�ۊcusO4|i�a��F�01^Jcgw�lǎ�F��������k"
�V�@&F,N�ޑgP,����hb��,�`� ��XG(8���9�v��ʳ8:��M�e��6�}}�� ��cjr���a��E��@�P���l�^���7���B���x���g���r��H��B�L�x,��I	� ��e�Q���S�&C�iIK]��>�ɨ��~c�K��Wn�]�W����j����1z�9d�N"�L��I�H����Q������U\�zED���ܢ7t�g�ލ���CQ�H�h����Ve	G�&��QW���"�<�`�M\�t��Џ�py1�0R�brt
�DӇ�`�p��C�]ܖH:'y3C�e��h��P�]dc.��/`<����t:���]���`bjJL8)J�5�89V�;��I(G(�ۗn�ݫw�����}0��_�}>�\'�\;�g���!H0�_�\���C���4-,B��(� 179��9���>���a���ɢ�����^8E���F
q���������[�`QK	�'}�|q�;�ؐ
�+˾��icvf�D�R	�3��5�X�j�������(���͡X��̅'�`��vms�+ח�6U�h�����:�Κ�������"{ ���0P���l2j"�T:)SjB���3#��i�X��F����p��L�y��y��#��f��iyԦ���hDI	�b�&-�B�)�\ܷ�[`ө��>���C麉��&���X���ǸK0hV�[�R�_�,J'��q$'� =yD��l]Vu/<so�6�/o��.*�KK�ɞ��M�AK�`��H�c�����gq�xL.��-N��`iq	fς9����p<�� x㕋x�IUL_�^��k׿���EqH�0���g�1�9�+8�{D�ۘ��<w��a���'�r�T�4v���#J&	��ge��f����[��VC}�F�#Lm:m�m9kXDL<����7A!�\?*B�S
J5�t:�.M���XB:z�%zj&h����3c�Ç`6��ѥ�PY��'ON������=/��
ʕ��Q�^XB���x�u�'��d��k�]xn���4N� ��/>A���&ON�Z��h��s��BJj0<����u�s�F�ޝ,l��͇��iDR	�{�����������p��/�l�%�)�ͣ���p��<S���6Qmu��P�X�d.���$�r���0q��A#,S��f����lV�����w�G��`���mͣ<3�t�W&.�N��n�����:(�����H2'�P�;�d��%��2��:� U�=9	�K�d>�c�y|��?��_�9���7^}��>��C E8>�a0�p�(
3'���Ӵ)�(m�;����t������`P�1
�3h
/EW%p5�;�F�=�.�\���g���>p��gXY��.�*z^lN8�P<�ɑ^y<�d(���}ܾ}�N�Dy��plJh��E�t?o�	]h�C���k���p�F����J��tG�^�|�ɱ��p��iA��zW�F����v}l�[~3(dȝF��q>U' VE�s�A�A�=6_HQc ����qk:.,�����ɒM&�P�,F�}�&����U_�>|����B�,�E��Sb����)�AM�a�dQ���S�19�������E4��<N>>��а�z�u�9���X�q|�����2�������Z���3�w�Hg#82��D>
xq��U�m�K��1�48zF\"�l��,5�Aτ��X�f�c�����#F����u$5^��b�)���ȹ�6�	X����B��f&��f4��@�_�R�Գ| Oʨ��8���� �ɓ���S6u���X1�?�C�����$��� J��(������?ze�b]kA�$}�G���#gP�;�P� #���GDsQ�^�S���g��~u�C�ß^1f��w:��ť�A���RCSX��OL���`��4���=TvvQ�w�sRpɴ��G�qj.�b�q-���㨉�v��A>� LR׃)�'	�ګ14��b�(�����G1^4��&3�D/MHR9IA������	A��@��i�ض��ߓ�����c�xX
�S)U�f]��4H�.R���t�s�i<9���e��9Δňx��6��G\(�����'K��ǠhId3���P�8{�Ξ�������2�t��F���Q��!IK�'��鈣�;���pxn�B
�X�܈{�����p�&m�=teD#
f�F13���hz�Ӷ�������!M�iq��ۈ9J|�-���a���EM�j�Š�]���XM.�d2� �#W�S đ"�E���������%(�C���t�eS=��(���������"@з���F��I����C�� E9A]Zes�@Ҽ��x"�\>�~����3���SP)8��l�A����ǿ�׿������{2��1;P|	Ic�A�J�X$�Cc�+�X�D1#,Z���6vCl�{د��V�K�0Qa4�a$�E� ���F��j���:t$T}
�*�NL���=�o�E&B0xI�au�N����lH�f*�B*��n�mIQCZ3)M,��b�������۫f0� �G����]���AR<̓��C�#�q�'���Iq�N��~U�a��d���M��,i��>�^}�_�G�����!�@Z���d���d����zu��$��߽����O?�K =��t���@a�}����@�E�ZD��|2��3	�B�'���X]T�C���`m�!�QE#l�8u8�\*$S{r۷�C������Fk�JW��3��H4)�*����so�
'�=���1<=���o�U� ��Ħ�F/,�i����n�t�N<���!��l���Ԉh�5�)֜n���C����o�A�}4����°tN��P�S_kA2���t�a�:6������w�S���W���uT���hc����Ƒ�8���!�r@�0x��k��(���V�W����p1t�1dG��9�VF��6f4~O|�I�B.�a�P��9$�!d�*66m�lU��XF�>���ɑ�-!�px:�Ѱ_�H3e���N��~Óib(^�v<ʓ�$�<���=w��a�ZP�P��.`�-��ҵ�;����&v�{ةT�^��g�d��2���r<+I�;@�e8�Y�:)�������} $\�p$"tLk�BGD�@�H8����2*AR ����(��
�}x	[���ԩ)��?0��W_��tiw,c�2���o�0y�lV���6�ĩ3�P�'���Q����SNe22Y�[}9���80T�u�����%�aK����0$����������X�.K�$fx845���N) ���x�}����[ب���\##�-�NW\D���G6������^9��0h��][&<lV�bQ،P4�
v�v+el��-������H-D(�fPǧ�0N<��Vţ���h8*�F���=�eԦ;)���{6��/�֏�w�E3O�G3I���͏��;��/�x}���3h����O�����
�ad�"?s��Q�(U��`�^��h���<������\ǀ�PWHs/���N$/MܠYGT5Q؄� �+`r"�BR�X.
��FO�������sL�g���d��`mm��	��X߃��C >FoEt-ѠFT��o�g�L�p�(�RA$u�م����Q(� #���f��*����[i�#4]ÛOB��c#�SҰY��i-d5�tI�)�_/Y���������oq���5���P�Ć��k{Y��bLnv�6;�|�b���
��c`w�փ)`�f?Q�Ǐb� fN�zۓ��x8�h(���.����ڭ����)��
�k���QvB�X3��#�Db���Ϧ�e�=ɬ��KK��XPj�\<�|:����!:V�������JGb���&��}UWL��'l<yr�g�L��X�eٜ�3���Q�JYA�9�~�+��>�i��ݯyֱ��W�S}�����/,�Ȅd�v�L�,(���#�&�?�	���$�е�C��B���"    IDATf�I�; ��R&�\$��~���o�n�b:��i�/@0U���y��N�fЈeP�g	z0;�?1���g�����Ui�G�)�;������Bgt�<A�NN���=Alo�����VeWˍ�.��J$�D$�����L.�Z����w��[G�����t�V�����!"Zq��\.줸;\|�0�ƣ ���`S���]����LtQ���`��G�i�VgFw�� ���cn���>���E�M0�g*�ZqM)
=E4�4J��y�q1-t�]8CƷ�A8�쀃�GȈ� Ƴh�UG!��y����T�'�q�S%�.P&�/w��!�Ϗ��W��+WP������șQ
�:A!1s�v(f�8n
�yqD��4������}��ŵ�'M!MC��gg��P���֒@ku�a���Z�F<�����H�0H@JN��t$|�"f�1ȩ�]#W�/Z(I�p]�� ;@Ŀ�Ţ����*T ��}\�N��24�P�2`���}���_?�>��pF���+Q� 9a�;����ub�\P���F���X	V��b[&���1���OuC9h٣9�,�3g�ҶVӥk`��84���OO��C��tI����Eg�7iU�2��`G��u�V����>�o?�B���.cii�[[x��!&'N���i�<��)\|,�����>��>�~����-xFL6X(Z��=�m'���ё.K���=����O�蠉N�-��ꇝr�M�B�|�z0,�`�4Qk����E�����6*mz��P~���}�� ��}s2������\C^f�fSGA�LJ��� �Ő��kv�=�][菳S�?����l��hH�`�p>�/����5N��+84[���o������'#Q��R��B�{VA\�P�Ej8��;x��1��섈��v��"n޹�z��:�O�������q���ID5�_�ڗױ�V�CmS�	b%�o�4i�D"�B��!<���;-�Ϟ)��7�mT�h���D�χ�Z�h��T#>=bco��r���Y݁�e0�H	�'Tq�c<$��ɠ&4q��'K�b���1
r]�`Á�\���z�uJ�L͟=���Cҝ��S��첀AmPCyu��`p��9 >�k0��p<�h�Z��G��#��dn�W&����z�@�HDt1�0�}��R\��t��-��4�����'���#c��
�������BĦ��V�T/��&fG���������+�g&1<0��;Mm��xf�>O�͋��h(ӡ̹�uQk���L�lT��Y�n��J�.E�����#i���`��7/LvJqc���,Wj��C�-���P�+���yqP5�y�#BӉ�R�17n0�
�d�@�4�����7?�ų�x����;�}�V��I�~����6JG�Fiz�|	6��tL���h�햼_�l[�{RX'��:21����V�]�[�p�}��ׄi��@�8���)��Ev$���,���5̔5��s}��'���g��'�*8x���++X�m#�˳��ĢC2iԮ%Ӥ�R
o�p��j:�I�w\d�!4{
v�6kM��5��[E��i=�0�#2u%���&�W&{4���ہYϣ��G���7��#��������!g:�u���-������05�Đ��0S7TC:��^����_B��x��O�k�p����z����>���	���NDE�Mz��<�F'��z`2Y�H�vTh�N�����&4����5����Q[����\	#�$�'�Hǣ�Z�v�������U�mc2B\uqd�F�&��d�:�F;�+_l��D��F�)w��!4�X\��/<vG&h�c"`��}��.&5t��8������j���r��)�k6��`.�G��|�_3F`���'���N�w��� �#��YV�v;�e����>��n��(��xM��3a�6�V�*FKED]7>�����/@ya���0t>A|�8&���` �G�Y��8�aaCE��/ξ��ͤ07;���+�ȠӦ���*c��,�do��!��M$��L|�6�h"1�T�D�D\b�6��bH2=���7�گ�2Ŧi�@*����c�����:������M� z؈����3x|>�@ߑ��IO%�f(�����g�*mX��A&��wlV��c}*�Ir�ר�>(F�V'KK���f�?a����(ce\���[3K0�M�f�n�a�-��F�A�a�ϥt
�h�Û��Ϳ:���	�TO@�g����L�^�g㘞H��sp��ZT�}�2��FP�&Q�!���#���Ƃ(f�H%��:"Aj���r����A�&�(&T���h����f"�[�P���!t���K�Ҙ�H/ű�Zu{x��4�K1ݮxLh���a��t�7`�n��Jv�ށ��̠yg���������7y�ϧ����]�)�B���&���-y��d�l�d��q��kɔRv�	��ȼ��Y�8J�x^|��? ����c�?����[���B���r&��m!N%���K�z�^#	<�4&
,�Ee����-,.�
��Eĕ-���K��߿ fbn�V���B��GwB$Q@8��l�nw��i!I���T\�ݫA���W�}��2�:�P[-v5�i(R�B��۹�W��VY����>8�T4�nej#�����R�t��U��xH�Ս�&��T^�t#e� nNB����l���):�(r�z�}T����h��:��&J0h����9zŹ��5x`a~�����U|��G>�	F R��IxJX��sPDj��-�92��@T�	G ��j��խ:,%�Zk�j�ֶ:��M��Qj3��w6�����f�,�S�˚��A�V�v�{Aڛ�ŀ��D����"&�
�^U
.7p�I���ZD&�>�P-����V[��k�	$`Z!��$S}�����ߜ��ۡ�jp��A�vS&�+и��;;�j���'(/���@�H�'�&z��%gp(`p�7�� 5�g1u�`�v���&�S�ޫǰ�6�����0���!�,�*�uao��:�FH�"�<��\����8�uҁ,�,�t�c�X���@	�1Z����F���E����~�B��bw�	�1����d0�S��wyhI')��ׅj���S�q���kJ4'�t�@C2��^l�u���7��v�Xۮ`�����@$;��#�`R{ �B�>���_����I�������0ր`]�餂��/Y�r��`��������ͫ�w��_����{��a��Y��&��8��&�Y���'���q��tO]|K+-|x��8{i���dRҹ��o!r���HG�ق5l�Z��t|4_���ql��S�R�����c�o������4����H"�'�y	=���na�nC5�B5��*�.��1gpЗ<��O����H� w�Sw0�X�����6�����o�p��
�3���^R����P
D��&%�`���o����]�6����0fR6��zH��(��0;5���I8�'Yw��2anb��饟a��e<u�0����C�5��w_�g�4��Kk��jad�[�9�����A'�b��[���" ���'Ν����`}��Tiŧ�	������rA������o�����n�������N�c3x��'	yX^,ci��e��ǧɌ��f�a��f,�S��^GtÃn�L�<w����>��ڭ�mby����a��1�d�s1�1M<�#ͩ�^��d�R/Mţ@r%y��Dz���h0�\.i#�&3+�hw:��e�tr��Q3�"a�g��奡B4�{"e�d騎C��������2���<�����[��t�@ �"��(̜Fn���t'З�`��>�vS&<��9}
���{�d�@7"���q��]Nx��nYc<��H�눇u����.� ����2��u�F���`��}��M�VJ�(�ObnnVLV.������P��F��g3���H�sЕB��gO�[����5O@ Z��Ke,o�Pm��ܩ��k�Z#�K��+ P���ZQq�<8IK��#�'-��Ɂ[(�z�v:h޸CG�����֪�0���k����¹���t������/Wd�����`0��G��"1q�O�I �E8�A$I�{���j7d�mV1l/�p7o���+7I���s�*#�THUir������3�PJ���"�!��P�y:�D��`i}W^㓓8}r��g�@��Ayg��5� ��k�:!�v:1)Qf����81���lZ��ח0�z��Z����#`��mf3��Pj�ϊ�i�F������A���N�R蟮>���)+�8�szX�j*���
�&:�6�ݞDKăDs9d#(�°#Cj0��y�B(����&�	Щ@6�)Q�ĠfJ9|
�C��s��Z����.���֑�*N�i�XC��ÀM :�+>��������Y��eؽ*���43Sq��I$�a$r�Z�I�뷙b!F]�4�#���男7P%�ays}D�i�k3�V'jЌ�
���'g03��>?�Z�t�9Ҭ��`f�F��'bF��Ve��\I����.	&?kЏYrM��+QZ�K���7E�P���l6�#��v�NO�x4��8V��C(���}2�t��4	����\�XNr҈p�����aw����U���C�f��Ц�B1$�'䤦�D�C:D&�`zb����7J�v�
ܺ��V��B6���� ���l$b����V�0�����i���%�e���A��H��?��˘1�����=�d�C�`��-ˑ���^�j�z��,L,�"5�y-4>��'A��ص�����!G��|n�h&�E�151lְ����
�>�gW���z7�N���D*�|���*���'� 5��A-%5��#ϡt��ɬ�A��S7TLO�`{{{��H����f���#�Ѽhh���׭"@�#S1:�G��D��D ��I��v�>�
�V�/9��Lc�Y���H����Pkqo���n��o�Z7/��R�Ah�3�V2l!����yf5OFe��Ԕ��sPo����b����N���V�O��3����pH�vDBW%�����韦���F0Ƞ�N��N��^���$?�Ji��l�@�mѕ0cKށ ��}���@�M,\��]��y�mHgFDä�N���)��3�l�	�m�+���dA֧�]���QE�& -��]h*�f�>����N����v#�9:|��j�MĠ�B���ƽ���٧+��l�C`����Jyf�e�J��1m\����m����0q�2%3,��h��n��g���r�[&��\{H� f�y�ٳ��S�g,o`��G���$�B�3�9x�ϡw}c
6|M��P
�	�LN�%���~O�M��L�|����g�Hgr�hcOݳh�|���ٖ������P��_��A�,J���d09qX��������a@����@�����%�����V<���ad��ҥ�t��k���Wt�x���96.Z�H�����h�C��\���o���a��a\81�bV��E�a�Z���:�VvQk:�%�1�Qs�h�üM�z7�hGg8j��Eew+�!��mT[D�#��'��L��b����!\4�}�!J�ɤ�,_wNk99���(��7`Ч����#��q����E%�MI�-:��<gy	n�o���#@:?>��NC/$�uicO������ ���������{x��sx���&�����{��W6������P�<����\8}-1�0;5��
��p?��,~��}���u�3%�逭G`�q�ہNF��D>���מ�d��Wu
�q``��A���~�\��B~��&ǋ��)��q�m��t��=�7���vc�D�(\-�F����qC&͒:BQ=2S�hA�\m��r���*�]�f �A<7�@$��p�S��4�h�����X��>f��&eځDB��*�3��Rx��3R���m�����O,ذᄑ��^�VC�W�X��C���A<G�� �� ��,
a�>����ϡt������Q�����l7���s�O�@jl�8s��l⨈و4�h�q�(S��k��t��_��-W��m�`B-�Ҝ�!h5Ӏt4&�N���ˉ~�� {�t;�>�~}��:�}�^z��VNw�r��ō5��z�.L[�^59�F͞�t"�q�h�e�Z�_���G�ę����B����>׳!��c��R��0T�N&��5��-uB4�h� �q��K��5mH�N ��y޲I@0H0_٫��o�V���F'�0���+��l!��RǎA��vT��CԈb�TD�#M�>z���ʋb�e9=L�B��������%M�1r�G=%\��5<~v?��#�u�ě?�,g��dq�J�N��c���R���iX�VV�06���Y����+L���M1�3ꈇU>4�\*��������6��9D���%D�סF( %仸�I�l���:M��دVѠ��Td=5�Z45�Bl�Hz�%���~�S�	�h(����`B�� �G��d��b�Z�Ny�n�g�p5�`L��
j�� �K%����HQ袍F�H�Tڟ��&>z��
�&0 ��̰Ύc����D�n��$��<�K��v�>@�T*�S��p���e�d"mȄӧ�r6F��.F�1�B&�J�Npp\��G&�ps��t���3����+��o�#R�L�������j�B1���i�-��Y�9�l<vj�ftp�NYU���g��@�هi6B���x1W";Q�~dH�۱��VjTik?� `���}����e?I���@������n���^y�X"���;���I�`�.i�3�y�O==Y �`D"V�N@F�j66Ē!�aX��]��4�+RD,e�!��'��`����K���_�Y"� �-f065�������akmG�x!���{�b���+&�ΎAg`$��۷n�\e�g�dJ�;U��i�a��HG�?����85Sv�Y'2��SN�*-lW�(7;hu豫�j���u�'�d!�Ki)t��'��#x(3��SAN*x!���v6h3��	H����|-^��|�+R��(��(
�<�f�����^�dp�?2�!T��@r���a��h�ljy�!��*҉�L�q�t��.�6��ۋ�Zj���``k�F�n! �)�c��T�R��h5L���GȦ38~h鴉��}�o�J����F'\D�y�5���%����%�T�.���Ԉ�&b��?�ы82��#�I��j=l�5�����N{�.��*�j���V1�S�����=��;,��z�s2<x�4ku4�u��	P��i�G�� �T
��r%��e:�=����@w�xp�#,]{�����:�"�2���9_3�q���ov1������3��O~������{����-�� A $ER$E�H��}��|�d2��_��$��/�%�O>ٖmْ,ɔDR�$H H D/l������,$٣�e5$p� �Sޯ�|>�mð=�kL	��s+Xm:m�p�A�Ȅ�+�A��ٚU��ʙm�J��m[:Gq�]X\>�>\�T�cG�w<��X���Y���	���O�P�=�qwqS��.�Ss���69u�[oV�~y��}�yLmFT�P�ө�xN�0�62l&�$�5
��Als�{��PD�BSnxn��d�E���CR� �b�\:M&� �JS+0�T
�j�V��Y��~��
�ŧY��b�ϭމ��f�Sf?yk9���4d�R8���3( ����]�L�q�nZi��W�n)�M/06��������)6��E��4���r��K���Y��;_y�=c&>�d�L*�>���K%Ξ}��>+���Y�G�F�����^���_"��������1��_]���k��'=E�&���6*.K���5��L�".�I#N�F    IDAT.��@W�?�Z�L�� [H�JB1�����MDK�;��)��s"��{�����ey�{�a����I2���[��Fl�ש�"�Tɗ�ec1�V�4�&�e��1�n��93=E���܏���{��ڳ'��?~�rr�/����W܁�+,m��>Idx���e�	����2���\�pd�_��$����qw�k[�Ԩ���xv�$_���~�V%�'�? ��ҹ}:����⫟���E�}p�'����8���A���Z�32<�ذ�u�~���U256_X��R�Ƚ�hH� i�
�-D��݋�j�J$ڏU�767��"�b���NA|��n����f�qJ�t8���d2�F�/�6o
2op]R�y�]�z&3�J]'���5��q��I�	j%���l�|"���Oe��4@[εZ��^����+��_���6g^<M�R��͏U�Aǋ�?���0��i|}���qV��*7�*^��V3tG���'�;|��k<\�b��дyh��8Ml��Eo��N�ȁ!��2�e
�Q�A��c���/�gq}���A��M_0���W��V��/dfs��d������\Ǥ�v�;���r�
|������L��Y�<�B�lNΊ�n���>��(fg�z�h���h�l��_"/����b�C������/����(�fP��R�,/,�A��,����.E��Ż���D|cMAb��{��!��P*j�P_�x�f�bs����J3h��:����q��c	�pu�q�4%Ւ�����qf&�y��1ffx����{ DRɩu���ey�J!�`o��?s@�/\x_�MRl�cI��{����2��lp���ք�luN�<��H/�+�:d�����ūBNޠٲ�rA.�l[��B�s�Z�v)EO��`O�f�BST.v��Iĭl�s4D"-[!�4����:��6�
��-��d�b��O��^�dɯ�l��[(u�	���f)/C�	�ǋC(�RgK���0?7Ov+��y��]�ۿ�hw�t:��̞�����G?��ne�,D��/�d��3y`���V�F�Q�/9�")�p�D0����=:�soQm,͎\aQ.���e�O?y��.+��|���|M������oϩ�|�D/s���>:��|�D�@�T�(�e���Ҷ��7e9&���
N)�
�=^"A�I�%K6�&��Q��T�����tE��5���K'绨��~A��;*
���mI�M��2m"#��u��V����� �[�f�:I�A���s󳬮��w�0��pZdH���ˍ�����$�=�2Q�=���aq��G��v���]c��c�]ܸ���fRZ%E�6�"�ѩ4MR̗��ʌ�qYT��T�y��`uH��.,i�@w$��"�����
�T��;L�����Q,�L&d�"�3��JW-a�HZ;e��ϟ>���.�-(�K�e&D����j��x���o[��;��,�eL�՘�cIm�D�'4-��
��_j���,&�@�LB��B�)�$�T&q�1^���4nC��٬Yc�V]�@�OWw�h��~���c�*)h籚Z�D�aCh�����M��а9U��A���%�������A����(>W��L.d^++��,�q�s|&H���n]rU��n�m^6�\�p�����G����Z�j���m2�[�5�^?���T����f�P�ְ�����r�t*��M�?���n�"�،�(Wz�mm����hJxg�;H��)�Xyh�@���iɃf3r����{e�+֣S�.DZ�ۈӬ4T�ⴘ�:\8䭮>�:��M�"�v�h_7c�w�ȗ��sy�썍��h���!��w)�^�fPB�[21���!�>M�葝f�bHv[U:�j���L^|�)�+o��"�l�l�-^���6��C�M��f�� 'Q�VT*)��J�� S̒*��|�.���ݻ'9�;�F��H�Ň[$�)�m͒�B�$�dk(z]�@�fM�ȵ� ����^��8�o@���f�\6I:�cc=��z��G���l+��h�]�����y�T���H���ؑ`��]�ilO.�{cRhl($¥m|�<�uAW', �R6�o�,8d�!�}���x9�Ӎ����8}
�2iț5vIx��Do_f������1�v 2�`�{���h3���22�u�߱f�Q��Uh�c��:#Wh����3�KK����%O��9_+P���ݯ�D��_�/YZZ k�E&����?d�1���Qm�|����'������-.r�L.��'N39���|����gi=�78�ޢ�L,e���}����kN3��V���	�>)�J&�2]���J��t�)�*$��l������d�'�*S�;Q�GC��ẹ1�!������irٴ>�"�:D�!���*�*'�o	pca{e��7n)�h����Q��4�{�&��{��$V������w��zl��x�t���T��Z�Dp�0�����G��&)-r%/�D=��`�˗^z�s�����O�o[�Y�{QHu��B6FO�¿�͓ėc���	�_��B���+��ѿcq-�G��V(�����"_���<��!�]Wi�d�	�����^�E�����p��r�D\ ,�uU��������cLO���©.�f��2˘x�5nͯ+P��mN���1�j�vb��'(��/;�%Ϣ�]0����ߡ�v���,K�ϖ������R����ϣ>��v���u��͜xLʂ�Og��0���������mO�x�����h��؅�� ��q��!\a.�MsJ-B)��$�
>���^y���?}���)ڎ0&�H�: �:�8:��m�;sB���>7���T���=v���!n?\�$��V���C�����slŶ���8u�ި�D���,ne��-���]i�v�]m�V,��z�C,�/.K�ݻ�x�|/�E��d3���f~#��R I[2��)	������(���5գ!�����s� ��u5K3"_Q5�{�.��GB�e�o�ex�r`٤����c}i�r2���3���%��deX 2�/������C��"�F�l7��>�O�AwD�A��H��Ig�-�L\�jGz��o�I��4��"�q.�ڮ��֫7���#4�YΝ�H2/�U�f2OO�r����­�U}77ky�|NΜ�!�s�MfqIx}���f��M����v�6��)��4dK&Ϣlݪ%"n3��
TK�	ML69CMK��U790K��Dz�\%o[��M9���L7�F�o Fv�j�����/ĵ�*�rim}�P�)�Co����F[�j�iڎQH&�=��C��>!�o��F].>x�M�����Z�Y��!g���A"��۵�?��參;��m9��wH�Z�`��3O�%�)���9-ɇ��U�I�B�f������N`����sTK⬴Ъ��ym=���x��?���.2[�}�$}Cae���tT�M�ϦX�NPE��G��Py���´��RL�v�f��Cb���2���C�d�Xk�� '�ᦘ6�N��@�WtLj�)�Nt�gU�F����s�q�Ʊ�I��K-mx:��6���"O�Y][��+W�X[chl�'�8CO$���@�S�K�i��t���2yp;���3	]I�g5��W�8��!^��.~��u�_�����m�i3(�@���J_�]��|���RxL����,[m�&d�%~v�:fs����D�p�MWW�F��l�זSd�mj&;��,M�1���j�w2RD6a�Tp��Fu{5�'�ʒ��)U*��d�d�� ]�FUX�*��R���q���%�RE�����	�"UZZ6�%�)�ǣ,X	d����C�T*h��4#��<��j�:�hP��r.�����(�܁js9E��V��3ۦDv1��}��3X
�� 4�k\�+�zA5ԟ�1�3?��UY��q��īѪ�I�7q���/�e����{+N�*����,�;<I�l�{�x�d�D���akrp��矙�V���v63In?̲�U�l�^�+Ȉ��T�)5P�2Q�9*풯$>њN<Bvu�;B��.���܆���E[.��ϦR�z�#��D���h�4Ӡ��ĹN$��<���ŀǏ��ֆXZ���H
ڒLdYVV�t+6:3���$�N�D6���axx[�����*��\W����T�;&��f�g�&g@7x��.�2*��MP�R���5ȿ�ﾈ���|��RW�������*2�<&�i*n��SGy�]\��fd�v,�l���{�x���߼�O��71�A���_aa����������+|z{�d��Yr�����
��,��Jj��6���yz���JA/�X|û�J��	�XJN�,I��ȫQ��I�&P��:�V+�!=�����M�}��l�����(RBD����6��8���Y<�~�Pm��u{�s��1R[��f���0:>J�ݠ�l�[L�sjm�p�*/��͠�'���P&Gt���}�-]�F����Ѵ���R��q����'�q;�z����Ziӱ�ɖj8<>�B����MO�V�YKs��O>���V���]&���L���gO��Q�o��6���F�]���ݼ�Դ���R-R���>��r�tь'<L�*�F���D6v��P�����;P���ڳJ&���+Z�0Ir��*�s�B}�F#d�rnTq{C��B��0]=T@�>rȘ���������Bje�Z#
�ZZX�P*i���ń]|;IS((0��lk �[��Zm6WVXX^�3���S�գѨU9v�������_�S����S:�/����;d�9���Z��gp7{���.^g�_c{Z�[�������J�U��|R�	EOl�T	E�:��8�Ts|��ϲg��g�a��<&����)v�ܶ����K�w���ؘ����{	�,l���e���=9��#tlBME��J�)E�H;ER٬�8}b//>�ś�p���*a_H�%��Y-�f�A���rki�2��B)�ƴ�\cbn/�U�~Ɵ�0��Ь���_��m�W����B"oj����Г�=lx�O�Y^X��(?�?q$���ScCG|<��1?���bmy�s�i�˜��}���q����=Jpx�@��u���R �~�ȫ��p;l��$�&'_ �͂�)�W1�4���88�ӧ�yxw��~�g�T&O0���/<�����ślgr��u��2�G�y��1l�*ٺ��Z(���՛qr5V�YJ`z�����b\�<�/�\R�xO t���#��j	�˫���{Y>��L�PZ�B���Qv~�� ���d��'H[!�
�e�A;�f������5"hqa�JE60���M�Ѱ�FY�zMf���Ae��Ilo����۲����RO���0n\��'|���h��p��ԛ©��0��H����8�F�G"���w��J��O���"����i��B���$��!��R���$1%�ɞP�S<}v����\Z��������I&J|ze���=�Q�f��N�j�V.������T�@�e�f	�{_�*��i��YT��O,q��!/>3E1Sesc�d.��7Q�5RC���N�nR/�(ش��h����i���6WW��r�D�+[59G�A�n�B��-�Lı���i�hJ�)5���f+��V��#qnݦe�p��Ǖ�.��l{<>��9'��|K+����J3 <�����0N��P8��N�>Z:m<6����9��G�W�/P�
�O�R�I�"7��銸]m�>sD#�>����)ľiiZ�D#���~�[3ܘ]�����-��O=���٥5���;Ig�ܾ�"�-j�\�l\��9�m����e���+hcd�KWH�uM������{�����1]�Xl�Y͛�9.�����V��Aw���p]w�;��G�
�3X%��ZFN�\[�6��������mvJ���|v�2�f�ǟ8�ީ=:��;����=Hw�$զ��o�;B�,7��`�R��s��n�q���Z��;|aL-+�jG_>b�T�\%ϡ��x�1ܙcsmQ!�����N0sl���'*鑕k1#��W>G��%��122��� ���TCJ#�Ů�֎�KXs.[�N5M�� �4��k�`�eR�F[�&/K	�喒B�y4�R��r�ɋ�`�?dr��*�_�yDe2�-�$T�L:C:�֯�uy9};�Qy�(���Ũ�M+&;��;8�7���Q�@$�r5y�o��e��
���fo��f�����4�v��ɑH��oW�zy��C�m���5�����Q��-%�[d �\�f%����M9~��oSʴp�\�	*�2_������W�V<�ir�U�:���?��s�%N>�U\��ᣏok���,� �ʍ+5�%0��,�W�4SL���#�w���O�`���M�6X]!*&�"ћ����H�"�!�i����_�������#vS3��K�t@|�ÑW�Uh�&�[dydœ���F<������h�BM�Ef����38�c�����5(�͠�ǽ�1x�)zw� s%�Z;��Ye5�P���+�?�����w�L��#ь#�Er�F-�/�>���>��E>��dqQ(uS��+�s쉽�񟼭͝`D����y��/��'Y�H0���}6�5>���ڽ�����T����ra���8;�*1��;�W��2�r{�8�&�ξ������� �ʂʖ��<OVm�fP�Z���fАe�����P�4�R�.�h�)zX��ܔ���`m�oUt�u��[$�q���gtj�L������.�&�w�p�һXJ��kib��h��gr?U�4�����Ӳ�����k�;��N
�%,�<n[MI��� }��*u��Ҭ,oPȔ��d�V��tz�ng�'O�a߁~5��+_�a���ek���X�eȕ�<��1�����u�,������9��䪄�ǰ{�(7]��N-ſl{5��2hZE�F<�����M._:����94-҅
&[����͎��P~��u	��
-'H�K�b�W�l"w��*��b��v�!MOO�j���e}N}b�3�XlmJ�%_W��͆RGj[�`qy��̱3��x�/y����m���7�o��ҙ�|��������+�D�gsqa��X���z����r�#�
�R��Il�SCLhн��.��I��?��a��@pP�p��&�vqb�0s����R����T������*R=�������F��.Ĺy�o��Y[M(�����m��/ױ�;�e�.�n	�.C$�=~l�_m���,�w��戄��:�@���WX��)�۸}jBcTs��W&�R�ꈭ�#�B� Q걹c��ϗ�V�"�0�R���%-�}��ad.��<�\N�]۲x�Y���V@I�Z������gckEe�c=A^�ě_�O:�8��c�l5�_����֭x|��z�݃g�[�C�f4���������)�b�{�tH�M���)���b�\�����-���Y+��9}r��=�E��L6�:m��|k������u����q#jE;�\�D����5�պ�>{iڼ-M��Vd{n�U�����J&�Ξ����nV�\�|I}�I��f3ݡP��v�i�7�,4�@��FΥ���x��f��Zj��J�� -Ke$�j��H$@"^�֭[x<����J�(_R��x�j)��i�P�eY_]"�b��}���V�396������p��ߡ�͔��*`��hY�x���;}G�(֐4�l�uQ�g���,���9�o���d�up��$�F��`���jSێ�T�F>���Td�����0�}�:8J'lnș�T�}~�fo��,,�ۢR(Q/W��Tm}�Z�nj&�ZE��!�I��3�p��t{-<{z/AO���-���E�-|f���U
M+��mX4B�A�M!�:�����\�G�߰̈OM(�R�J�7����խUq��.}O�����ZG��5�+WS��\������ϱ��A{��-�`���ş���o~�Nzs'���X�p�4���30�w��ǥ�#8�%���T|�VSM!;B�a��MT��;ͦ���].J��Ȟ<���>�-��3�jm<,���    IDAT.����=���̽�����"2�7�g~��TU^|�D6_&��`rȷ$_S�;�WY!26�j���'FH'�,�/*�f��dk�D�&>k�KG!M�!�fP`9fb�<��1|���]�6��ϧԶ�ZC���|D�!DGe�&��m�+%U���z��FF�9����=V�3(�`��oh7�����'B�$/}1�K3X��J�7��/ĝ�ˤY"�n������6%E������x��W.^��?#	P���ř�����|��W�%3��&֗02��o�拚&�I�@?�F�t��;o��i�v�bʴ�H�i�vv(e6	�;�c�PH�?�Ms��4�N���~x�ŵ�H/�j�JU"+Ļ&/�GA�jc�)�\���/���;(�n�e[rn$������am����r��d|!�өv*��wd�����Hx�LM����Rl��e��C&ZKb.�h���&c3h4�gi3(���\�t;� B@����j�����ܢ�f�l�:�D��T�
]1��9^�qN������rF7M�x"N^��ˬoW��7���Q�����c�8{j?�I�C6��<��(1M�x��;�eY%��q�X������g�ЬVI���Hp��d���\�ŵ���/��I���Wn~m�2�i)A�(@��6�n��%NRȈ$�H�L�U�'~R��lB&s:�kjS�ҧN�|9���*�T���~&�e;ء���l����g�ބҚnReR��`�>C�CJz�)�HC���/J|�a����_e1g���ҘH��2p���\J`mUx��^^|j�����{�o�*��hw��_}E})���)VE��&�s��'���j��ȵI�묯�Y\K��iQl�Lׇ��Q�����Q�Uȕ�8mz�M�x�	�6ۛ)��Dna�;~�`y���f���xĊ-����?�x	*`I��_�j�'p�="�*yn���D���U��y�^�BIT��"�l�\V�|�b������e��(O<u���9Lm�H���Do_�	����l��i3�fp� 5{�����dQ�;rK���cn�y��8G����Tl��*�:m�+kku~��9b�Y��AjV'>��Rl�Rn���^vM���3LwO7��f����145E�i���������$t1�[ [(������Đ�6T#C6�2�a'5I�fM	�(��?�ؠ�LT*fj�6W�����\�t�rMr�$��JCv�E!V����(Zv��&����W�~l6�8�3�'�ʳ������w��B�52�A,�:Dp�E����WV�%Z�4��:M8ԭ���3ۼ�ݿ�f��S��ǿ����^{�
�:V����VS�z��������vX)U�XIzV�Lq`�=����m�8I��Z��[�?e+]%�5�f�����m|�Gg�90��R�M�����C�6Wp���N���rd<���t!�T�����N�d��1�����6���F��ݼS�۝��8F�<��S#Q�c
\�R�ƙ���\c3U�!P1��JF`S g;�%f˰��,�5s��*A�ɴ�eW!rC�E��*!�
t�AW$B6�֍��z�%
E��\Ș�/[s��y�W��>�X_c׾v� ����aWO��W�����d?{���ū�-@݅�;������ÃXC��4D�ӪVi�t�mL���gw����n��&[�&�o̳��n���S��4�IL096����
$���훬d�<!ZV7ݑ g�S�l���!�B��I�JB	5�v�ퟡ��QH)�նҐ,�N�ǥgM.���P�_�8w�7Tj,�K�Цg���{&>�9�0�<�[�F]
Ry��r!��\O!.�t^��Jl���z4�_�~P����!��RCɶI,�G�2>O>4ORd�"��W�J|k��Y�v�+�B<�#�8�m>��m>~�;����
�1�|�q�oJ��1l�.i=���JY:�
ӣ�<q4B�PP�D��K"�z����_]ȱ��M�.һfK�D|��?���'���|���+�l������E��{v�դ�W!_�Km���ۘ\���z�N�c�&��N�j������,r`r��P�/��\�ڨh$�Аo��R����:V;�l����Ǖ��M�֬�4T�y�>��+��6��?�r�Ĵ����`�^K�/* ��0GbcD�&Н�D�I����&׮]��_a@�?����q�'oq�Ϳ���Ƥ�`��Ch�>�5����}8�=ؽn|!��Ē
@���x��<">>��?���F۬йD<����P��%�:v�	Kd�ū�t��oƒl�l��,�'5f�̑F{ͤ�b�i�3%2�"�B�@(��"�;�ي�e$��,�},f�,�����P�Ǐ��Wpia�Ƞ��<?�X�D�����/yn�NW�U6�R{���T����j�i2"�>�sQ�t�)h\+i�fp)#g�fP�g����rio�޹���~����F�;�����`��n�e3A� 6��vCtȢ	��ܬ������`jU	��%R�2.W �͇��Ә�j�@_������.��4O*�ԗ�������1�ɏ?&���+�gfj��������T�mW6�[ަ޴�MJ�f`X�	�fP�t�#�U���'9s|�|"΃�ի f��nZ�,-g�+��FHf������F�!Օ��*��Z�I����γgx�v>�r�d2�Z]1k���Vy�L��l�AO�G/ҝ�tz50<�96�ZY����,��;;���_jE&�h3�i��iCԅ6e�}��J�YU����v���7�*�e�'�Sm���	����yy������t�ۄ7�g�KW�~u�����8���v���\!�]c+���ւFT;�(���VÊ�$S���$E�Ҽ��}��?s�W>���+s\��M	6���n�^RY(T�X�ݴ�"��b֘.K"�x�Sֱ��P4����Ѩ�t��x���.�nuu�l&����\y�VIo#�D%6��H~��C&�d��=��ݻ���L�jahx@e��?a���(-��͠�����S�>�=M��!LΠ� �����6(����V���
�#*1�(��ȧ�.�^JPpC|�>S����	<2QN�4�M|��F�\����{(`�4�?9M_���J�ŕ�v�T�R�B�i���#���W(���ѫ��Q����a"������1>:A�@�q����![�Pl����I$j�L6��������A�ɽd6�8&�z8|ޠ����(;�!�{At�p��_�n��#E�l�+%�ܥS�r��)�~�n��Rc�������2QW�����qt�һ� Uk��|��J�m	aO&���R��3}�����Ufg��o��]d��G�8~$L!k�ß����Y��^~/^S����H����ᵢ���5�߻C�V�m�R.����\v{���&�d�̝�k��3L� 6g�fS[�ni� 9��]�Q٢V�15�O4b�vV��X�����T���6����ژ��g�?D]�z4��.�Q������T��]���!�ɩ)R�K��Z�<~c��l͠�c<%Z��Td7�B^}Q�z���eJ�O=N(�gt���l����bs�=:�����*Y^z٠��6b)��{�ޱ�x{G4`�֖s.A�������-2��F�X��V##�LD�>[����LT�9]z��9��y��!�n��6�e;�Os{�͆	���y�S;��\���8�ostx����OgY����,ŧ�e�m�~ױ:��*%<�6���F���3J>��h�\^$l^%�5�2%_��K"�7(�!��A��\/�l��wi��0���
�I�5����vu���f����XMچI�!I��&���Թ:lnX/�ܹMtt�CGQ��=��}l����_��nq��#H��O�ѪJ���Q3��� ����CN�6�����.O=q�=�����Q)�(lm3�7��H��x���9��#ܭ��!���'9�o�`X�J���O��p+����PH���������fG������1үY�q+�5	���vP�A��5��bW'��p������A��hTV<O�P?7�~o	����ϛA��E���t���p)R-�ǒ��>B�͙x��?�	El�D�[w���0뵖�W���{3�>�=��,1��L�[7����́�5�llx{������;ߦ��d*(�P%������O>��wvm��<"��А�쀋gO�7d�����/o�C�fb5� �ɱa����b��*v�����P��2�%�:�𻃘L5����-�,d�X[L�GٿgVaOd�p/����d��'�7��-A2�����P�ޖ����XZ*�u&BE�4����
S����"�Pi�0�#t�n���٠�_*�~$4����0��r!u�HD��h�t{�twQ*W�[^R����P9�ԋ���ͣl!��|4aiw��:,�ի|��
�:q�1�N�n{���f��@`umi�- I^���=����z��^�RGR#�P+�q�Z�b׈��6vfriyoZ��m䊒w�aq)F�(���Ɲ��kX:9�M�224FW ��m���E�-/Ӱ9��x\N�v<6
h��F*���Hvc<]P�M�*C��J3(����͒;�#�0����!��~��LG��B�̓�,��Ic�!�nmw��B��ttiЍ��A�M��T�4�F���E�g"ʴG�������/B�D�?���'?{_���{�����f���!��q�M'�� &��0�[
il��p�%ҡ�ԞQ66��g/d�$%�-W#�'�/i����b���̮.zz"�jU����b�7ﬓH���+����W�T�ŵ�����q3�pC����Q��k�_l%D\�����	G~��a�86��B���9,bf�պ�E�ig~iKe4�,&х�&I�,j��'mg�"�J��Ҡ"�G���owj�FyUV빬`��x�^��e�U��[H��/k��XE�!o����tu�0>=EM�探`��,��Y�wyg3����xM�a�``�Yz'�`��
��&��j�P���]]�w��y�ߥ$���l��H�S�ɥxv+E��,���/�E�W'�k����R^{"�
X��5���.�b��oQ*��Q6�����<�x��Ԫ�e)4I��&�F35aU��*o<�o���NP��ɥWiwjTjf\n�s��q;ƃ��� u	Do����
��OBy�E�ܶJx�}3(/H�Y?ȦA��ecҫ/
�a��V�yK�Pm��T�`�����w4�w�V�]$CCX�un\b���o@y�U���(��^=E��aLN	�׊��F���R��w�9<3L�g����H�[(��8ۉ��nfqJ����b�����H��ScCa��[�έ����mr��ؙ��इR&Kz{��d��L��f:u��9h�B�].7LJ���\z�d�U\5%�f;x��${f�'ϰ�BN|dV�O\�>ǥ�w���4-�걣�CY�Z�d����fP��l!�m$ #ͼ�fvvV�A���M�ɚ�C%�Q�2��hԵ!�I��,�= ����}�)=rjlK��ҽϸ�ޛԶ�t��pOC�m=��O��Md\6��z��DW"%*�O�/��>�w~r����*���PSm�c�|���qt�������G���̱qΞ��֪jN2]as3��#p8l,mn���ޥXk����/>�H��w6�v<����������nb���E��eͪ���F��LWa�j�+S�,1=���s��nߺ���8{!S�r��}�ΐ$w���eUˎ�)9o�Bfo��R����� JT�4vR@J�115���"+"���Ӑ̓�6��*�Hy�EݨS*��ymu�R>��ǎtiQ�wj�J>��o}���}N��Ϳ�:�J�^y�����J�{o��������)Ů��pxW�ϟ�C9[�w����6�@��ɡz	��s�\����o`w�������_|*J=g��]�P�R1�`��]���=._��@W!;o���׮��ɸ1\�ԓǘ_i�w>�e���5íٖ�+�>W�=�[;X�e\��c0�烟��F��˯�A�P�ڽ��e*M'f�l*�*�`<;��i(|Sm�*}V�����BF	�"��������&��f��p�r�����Җ����}#!�el-�lpR(�~���^�=~�F��t�ᰗ��w�ǯ�)��:ǟ8��k���h������%�w���><c#X"ZNc�.ȳJb��N����d�[]f~3C6��T�1��ˁ�	���ب�w>!^l��ۇ���}�L�h�\*3��'����U���u֓9�E=#N�bt �E�zl��K�@���2�>\#-�B�5KN���x�u`��㲫⣞YSƞ���ߺ}������:`#U��	�l{Tn (��l/�&)�S�����(�bH�����q�ny��y�f���K���?�!�?��֨,�eb$�i�ڤ]R���V
9��]�0��i�0:8��U����p�o�ޚsZeȟ5�s��'puO`K��G2�6��
������,�ns�'ai�T�\j��`��dl����Y��j����
�q8;<��)��6�o?`;QQ���� �s�������q{�|��T�y��iT�0�e�7��g�ᕄ�����T�auK�r	��`E
_�`��F�=\�tQaf3�����If�ll��l��I����h�'͠�#;�A��Y��ԚV�7r6	PO�X����fP��t3(QimV#�LzQ���W��
�@*!�#c��~��ҧ�>��f1<�>?��->x��!��͠OnmM�^UX��4���� &K�]��)�G�8yh{�Ir;N>[&�Ȟ�`���ްJ���#8]^*�,~������pwSӂ��ҼĕX��T��\Y��������r,v�|U�E�n��J|v�!�J�7�0�f[n�a�j��L>�E���7�e��0�\��H�D�ds�/�Ied�V����D}�jFi�m&���X����Q�#5�MZ��,�Q��t� =�4�J�ݩ�����J'�WĦa%�Ji�&���������/8�:ۘ�^�;-{�@d�FG�Sz��vڅ�X�R�0.��$++�� S{�lmUq8:�ԤSE><�vۮ���P�\f�F5�H��)i��R.VY�Jron���8���J4�g�߫��tf[�!o���UiJo��y�ne� 9kM���-Z�<�j���=�7L���u��P���[/�'��aqu�G0ò͐I6�;�Im�E�b<�tF�f������ng���D��" �b��%���Z��2!�@g��Щe���֥�U<� S33ZH����;�9V��۬�����N*@�he3h��`�]�U�{��;�͠מ�Y�k�E��~L�˫1�|��V��MBBU�W�R]��S�����a��و%x�+dsu��A���V������(��n�`�DQ{���4�	��:Ȇ�*r/Y��ߚIV)`w�W����cf4®�~B	\5��֨f�jc�A�[8�]�q���lc�.�j���af��N���A��+�DP�m�zJ3��D�����0pۢ�Wo�6�R�ʗ��֠|J1;?��j���{qz%����H��u���g�(�f����&`����c��Yz��S�I��bq:YY��H���gf�3>A�]�\mh�ܫ]�>h�X]Mq�ӛ�ꋎꔨ����ʳo����1�,)jlnl�pn��x�K�ZF���X���e����hs�����;lī�Z6�j��Pߏ0��^��vj��ܖ"C�^�����m�q98�a�>Xa=���АbPiR�HK(�M�gj�7����L�QSa�Y�F�Q���o�1�ÚEh޹��='������]цp}m����S��ܨ29:�����[|���Q]��@������<��0ݓ�U&ۃ�o�{��� �cfW��+�|ti�?��o'�=E,�ctd@)ewn\�7�5>��4_�ˏY��O�s�ff���~�>�\���?�b���������_���[<��YN��w��=n�^�.���}3=q�/��h[    IDAT�W�����g��Q�o�v��r��A#�Z��������	�m����3�ڗ_#S�R�7�JT���>�n��l�S3.�We�"ŗ,�G��/�׿�m���ʷ~$����642������y�����8�%��h���|C<P�}%�ߕ�d�2s`��0�3�K�����l<���N����5�F�W^{�d*�'�M<����Yz{tWdW0$1�XZyN����?��ﳲ���{Dd�r餒&�����{$�m�����R9����j�񟿁�ꡧ���T:�����︷���-����ի��o��HD7ޒ붺�������.���>�.
��JQ��^�S�%��jjR�l�o���x��˛ܼz�3���=%���������������	�]�N�
�����Jq!�@)<�[f�"��e��_I�����^
ق!5ٰ;�K<L�ݺɔ
�e�4�2�1A�R�������9r��v����d���7�Ο�1��*GO��7����i��P�����G����;:�5��r(~�\m��T��׏��?�ڏY،����vc��qѤ��q򱃜��~�y�~v��h7��M���l�ǹx�2�̘-�;v� =�!>��ͅ���/a~v���/*D�����S����Iν����eZR��L-.-��f�â���T���!L����u67�8��Y}��M6��_��d|p�N�jж�뛥��XM���gl|ٚ�,d�"�JG�jn��h��R���܂�Of	����"P�A��rÈZ� P�����jV���^�H3h�4�q�].��w���V	�N�p��o�$��)�n\76�lL��
�<��>N�õKs\��3�nA�p��4LRc��<�?��_ck��?|��X,.�!'/|�۱4?}���
eKDC.~�7�O�����+)�/����?��w��ꦿ��Xl���e콟�J�s���9�sF7r$I0Ð��p8Q��(Y��x}]7�Vm�z�zk�`C���[^�lK��F�HNb�`&@�  rht�>�����挮��� ����}��>�4|�;�ǅ��3z_���d�v�!�ͬ�v�t��A���=Ȯ$p|�wn��YF�ɋ��'q���-�$�@h��.������\4�S5d]\י=n)�����f��\dqmE��6�ڶ�f��*�D�̫�*#C`Ej3-}��3gNɿy��Ӳ6I�Q3x�=�f���PM�䪦kR��|1Dۇd:��0B1�Բ@5���glGGDǭK�1;�@�c4y,�TVt<�SwH#u��$��W����[�jX[[��"��K��~�\tt7���:>�tSΙ�=�Ѡ�S��He`��D�z�[05��əE�-n�kR����y�ح�T�M�©���hB{Kׯ^E�lE,�UבΕ��\@���°�!K6�N������'�
HQ�<Ys�l���_te&UT�J�Cqo��D���d�dQV��@�)�N�¥��t�qBu�X��e��#�AY��Bb��4l�6�ie���atuz��7/��CWA�<�"a���0�`g�]��o�׃�����c�@-/���4�_��2�� ���b�ZDow3z���]�vA>*%,Vqq�>f��2�PI;�j&�phz�٬&,��b]�M��17���9	\Yͨ�����3Ȓ�L�YP>J�$���#��7���Zo&qr;j5iy�l&6�bl�_"ݒ�rD��êL8�&թ�M�
LM߇�t���_6R.N�����M�22u͠%��Z%!*9N>k2܂���h޲Vo%n̤/VL�լ�:�[��B���&�@V�ڸ=l��cW/�\�É3#b����Ck���6��	�si1�p�n���*N��*�+N��g�څ�ΨX�r� 7:���č�9|p�
9+"�X����)hf��pV�݄S�|����N�<\��p;e��J���7<>"�6��qDo��u.u_���R�hc�����6Ѽ���~�FǤ�a�Z#j�4	R�h�Kz��
���"<���iq�b���D�̢���r	S�.�d0-4�E5�l��Ҷ;�{�ք&J{jb�xn/^{��ϯ���}�瀵T^�4z:�������^�c����������f<�]��Nz2��B^\�>�k7Ƒ���3����a ��"ӈ5��XK3:[�XX���gF�H��u*�A���T�Z�MV���ICo���'�I���=(���6n�B�dEٮK3��+1�b$!@!�&���fP�v�.X�d�4�x<�P(�[7�ZV����#�?*�U�Ir�U4�KS�p�g[[]mc&���!�Ϣ�������]\<����@{K s���l�a �wD��'ލ�M�h�?7��@g���{ľ�?�5l�0tO��
~7��䳏����
���������-H���Z�t��W����:�w�i0u�.܅o}w/~��[���|������6������y��l�˫a|�.z���_y�/-�셫�[D�%]���e��
����Y�/�"&��8y�=��h`��8��}�K�_-�~�>�� ���<�Ej���9�S�º6�>%l4���D׹����ѩ��,�)ք�x�&�d?���V�`�B0�_�SQ2@M�3Ud6�XߠF܍��68�N��[����Oࣷ~��ыx��8�揥�����j�h��������/��Hs��`2C7���{���/��{�{�k��a8�1�`13	xly��V�O���16V����������'_?�Ĭ���?"����3K�XI��������3����_���"��o��(��p�=������x������?} ��Y�������@�\GoN�j��o��_ކӨ�KxbO?~���mc���?��&&�$�ᔭ���w'�j6�*�\D{�Ua�oCM�OR>%�\UT#���9gԩhl��*Í�Y�3��s����A�8�RM�&V�i���?B�%��[�)�$Wn{w��\�/��{���a�����5\�q^m͌3�w!Լў��:�T������g��o<�������7x����I/�m�R�����x������)�jD ��_z{�b8y�Ο��p�hNf������Ӹ0��S�.�[^u+�}{}p�èv����׾�9\Y����-v-:�6/���0�Z�-��:�/���E����;�ѐ��-x��������I t1��ԡrm���*Ү+�9���Ѭ���@kI�X�x	���ͭ0�U��>B2����!��.\�ʪf��J� uO��[+�X��Eoo7zzzP2k�jm�a�����8{�W(��j�t�%zIoމ6�Q6�Q8�^hnF����x��܊�wa��&n�L ��$���B������m]x�@?n][�G^�l^�G7f������XX� �/�{�Ж9Å�S���Ux�Q<�³�۳�uc��r�����>�H�v�8;���e�v���@X+'ۥ<��k�{k5�ޘ�=�W%�\��Q���/AG_?��ܹ�=ԏ��-�����
S� �-׋:#�TPj�}��c��@�&����[��X�"�8F�uX����i0�{*����Y�7i��n]����#.͠���f���z3�,��?�H� �:�C���4���YM�;~kT�+G�a+V��[ �̊�8�T��� ̙�^z�^���>�ߟEs,���l��q���R��=(�m�h�x�	�V���%��e|��O��˻o���Ձξ�x��!�~7^{�Y�%J�~�.reJ�<r6;tMjv��hN�Tg������azr
ͱ��.qn��ܸ��c�a�c�*7Q�@���M�8��Õ��z�xl!�{���s����^*sa��G�2�`�){3kJU��ea)ҩ��Ç�qkNÍ{�#���f3�����lAx�m�k>��>x�n	r�qd�ߎ�^�'��+�Ǳe��O�h�T6��v���=�x�ݫ�{�B�
�M�����E�XY|���U�8�ڻ�`�,x���X_K���G���f"���%$7�(�) ��o�._ o��,uwv�,�T%b��D�M�	XK)�wưu�##��5�عG2�V2�;>�?��WH��ο]��#�(�h���ƣ���$��!��4N��:��)��Iw�H]���Q��9�<"�g�[E!�ǣy���bC�>r�ӉU�����ݫ����+*k�L>����KS?b�O!ַz�U��2Y�%>[	{w@sXq��Y��,�A�f8����l���Ͽ��Ҁ����b3�GSs;^{�(��,�}{��ޖIc�j���g�����|�gp��x��.�t7��Xx8����͜޾���h�l�?��Y�?D"�0��s����b���o�RMc�@;vE�;�x��c���Fw_�8E&�	\�:��DA�j�fBA^ P1R�$�m�*^�Q�B.Ş��F�Pu�Ѹ�\ݿ?#�5�ҧ���f��S��S�V�w��#��R�K������\)���6�KeL^���'�|x�>��Z��Z&�����q�z3�M�t�L&y��o�Z�6������,	u�4=j���9|�K�Þ}��ٛ�qsz6���V7����X[^�;oUn�D��؏��f��O�cn��{��?}������I�F������αIܼ;w .zZZăM��'6�`� ��o~��͜(���/����d�$���w09����Ʀ]�I,�-
IIi�ԇ�y��vcR��s�� ����D���0�'��g��_$'���8���B�,�&�Ƽ:j��b>���*��]�=Hf��pk(a��8.}�6�#�.>�'��kG�o2� B�C�5��f3$G��I�V�«��ͯFg��K��qs�&$�>��&������������������{��:ǃ�\�:�յ�v�u����풻���Ӹz�&�ع��;/bi��n`~y�r�xϾp�h���XZII�t��ZH��
źF�RqG�ށ��0$���AO� v�m���?�����tF�%%W�`x��勨�7LTC�;�mu@TDh�A�8]i+B{-����h��{3H�2p�41�"��g���*�������5 �N	E�S���8B���@�������)���؎c��������n kC*_ƕs�Ѵ��̓ul�3�fr	���׍�~c7<,���q�����j��!޳۷X��?��s�������1���ݛ˸q�&r�4\A'v؅��4��E{���0�l���a5Q��޾��Gs��<x����k��?^�{�E$�8<��eE�#����,P�)��h��׎���t�*~��B���p�Q�>
7lt85�>r,]fH2u�tS͙rp�<OR��fOr6�)Ϲ2�j���f�6�3sȤ�p�z�a���ZC6���Y��&�pX���$��z"�X[��t#�لߣcgOf�\ů��oPK,b��!��%\�zFes��f�e����vvC�D�F��)�����+Obǐg�<���G��(HD��fG1����_���hnv�?>���EC!l����p��C\�x��`g������]���å+�8�*Z���������|޵dV�]&�{��~��{x�hU��ig~���VD�T5{��2ڣ^��s��,��0���o0���=O���9\�~Ob��X��h��t�T��\��V�&�4�R�P-�S���2٬h�[Zڄ�0����51�b�� n�
�C��tN��M��1Vkea^��w���U"��[[��WN���_#7{(oH�@�>�-����$\�>�!?4Onw�c��a��A�ǚP5Ӹs����GH`Z��^�`_ +ˌ ��BA���ż��?���B��N`��"��3���=����,��b�`�n�\õ���u{�l��/m���F�=B&U��↡{��S��PD�ۅTj�B����a�3 �wn����:Z��`�t�:?��͍�ɳ�% �u�F"�E���$�����1��l5jm�D�V���p�wy�cƮ��Be�ĺ�. 7�G�x�𬤛ybcs�"o�adR���h�zq��;*t���JR�19�6|��[mD�s;�p\�8��QqQ-�$4�����*.���͕My��4![!�n!��W�{.�����Br##�דv#4q~� �+�d���χ���W���5qP��C�'��xD�U�H�7��	����,n�MJ� ��q�V6�W�V,�TLb�/�������Id~_Tdn��B�5�K�g1:5�7�u��}���5�1����i`��x<$��^��
}����C�F�~����: �p f�
�Ӆ\>��{XX\E4҄��^�\V�\X�_���i��l���|.�#�g��ā�8zt+�z�:���a����ZW(fQ,f��X��7��
Ο{�S'.C�b7��/���;�8u�4���I�+�20�/~�>�`��^��'��s/������h���V�ayy	O܍�_݇����G�4~��?:xҊ�L���@_w�eR�yܛǖ�N��t/E����9$3U8=M(V�'�)�7�F`��7����1CP�zn���C::e]m���U�2סX����e��$i#�eV��sK�W}V���Db3!� ��F��nSK��5,ύcn��� �E�(�*iٓY�A4�@�{'<�v�i��n�{.��;�ҭ�p����Y�\p,/>����_���������o����[�%�2���1L�Ϣ��gI
���7p�@7��{�a~q������Ʌ���A!g"�H��{w������v�G?���ŤhA�u�jQp��a�Sz��E��O�#������7�ㅗ�bu#%([�@��Ņ+w�5#��#���I�j���5".U�O���_�x��ɣ>s�Q/�0o�KGr3-Y�td��l-u]�6��lH��Uh&�A*����A(�������vh�*&�]���SH��@-� �f j&yc;ѹ�Dz�Q�6�R��?�Y�n����?Fb�����;8<Mh�ى�Lv[�r��1���!����^ƭ�$4����-x�>���'11>����ol�;��}{���<����N�<�#GK��?��[�����-C��d4Bgg��wG��?�������M��D�i��Jm.�5�¿����uu�"^~�s�w�R�"^|�Ｗ�c��/Т�bM�
�n�Rv�8��͠Ҽ�~3�)gI�S:�x�\.�Lx�B33Ӳ�LWf��͆�W����Bs��#on�ɔ7	"��$n�=]49(`��(�];��gX�� �h3�};�Y���<��Ν�:\RL�Fj����
�j���3���i��F��H$�p��x�#8������}�2FoO��k+q$$֗q��n|��v\�[�~�sAn��?|nOǎ���{���!�}� ���DSĊ����bz�^}�5�q��"&&��d?-U,���k$n��(xK��b~�[���������ױ�Jcߓ$G���+p�]`p�
E���>�I�PR���gN��;�/�魚�ә��;'JM�����@fy�y��ᫀk����%C���nf�t�:����)�¾ �0��<N��,>���ڎ�I��������	1�!����{���5|��>�,vh.r��$�>�/>�%��;�-c|b�++�����E[�##y��4rf	.��KKhn��՗������߾�K�.`����/���\��8�\�->�SE<��w�p�F��::��ܑ��;y�P���&�R�)��,�J1'�X؃p�#����e�fK��2��+��Y��{��R�s�T7Q��c���e��:��{t�ֈ������z�H&�X��L��Vr���*6*��S�PB2����6;"�(�>�LXB^'z�<�{����(/L�ɧw�b��¥3phn�i;`��1��m��i���GMg��w�Pή�+����C��b3_�gVp��4����8^���������Y��|:8���]xb� v:1����q���g�=�=;xt?�+W��I(��`v�l���߽}��x�����Z���    IDATW.�E&[��QM���/�+���P~�|
�����0��ׇJ����uL��cǎ�Ҩ�>S�K��6iΥ���~Ƞ����e�+f	�ZG�,��d�T3~����Ű���g��ê��ƞ?�'���kgs:��l*�׋��N	�紱�)
�j�޵���[H�g3�)�';eV7<�^D;��n�3��٢�ހ�� �������\wF�0?��xK���*)LM�`yiժ!�o�d�N��I�;=����9t�u��/��s��}��b�"�G;c��A/R�2ܟD$�G{���Y��%1<�1���D�Z�I'O'Fv�� �аT�^����P���.:�ۑ�桹HdLX���M<(-����Y��������5`սôZf�(��儦HfR�^	��$�����QTd��y�,/���';-�-�g2h����qჷq��4��W� � �9�>���"�6W�Y�%!?,ּh�K��m�pT4���I\���eaV����DoG���8��N�}�j�_�y�N&�p @�v	���v#q���"����}p�n��X�`��:�&g��щ�-1�CN�]���y�Jk�.�S�%���YH��ُ�q��-V������%�wt�pYp��$�����z	����A5祦V`��Z~�Em<%k�;��W�J7H7�z3HJ���,�ͺ���E�(�Y�ss�3�,B����ai~�j%��(-��B���=�T馔��}�p�٭8�n^EW�6�X�XU�5��Ãx�a|p|�n�C&]���A|�K;p��m��8��h��k����x|'?9�]O������+�8u���lp"�K�a�8�����d��tۥ�)��U��5���@_�������~�;�O���Çax���MLM/��
���D4�E"��z� ��$�U�����B	a�4:x��j:��22�LR���1�HEWEM���͠ZԩD�\^���V;;+�-q��Xz0�G�ב}0
��d2h�ea�W�!�X����ُP�0��6� u����E��я�m�}�S�KXZO��y�;9Ia��>��� V���寏#�3Qsy��K�bK�׮���Ĳl�T5�x��~x�N���G&��3���}�������b$�v�d�|�Ž�����o�5��/�VK�T�)d��ؿk+^xv;jU�̊8f^Ŏ��Qs�p��&��(�M%s�HS(]���E�iu-�����9u�4,j�KN�����+eF�5��$��cR�Bb(CG6���2m�}�"�����_ˡ���^���S؜��Zj��f��5�]۞A�g ��t%��g�J
��/��u��#�|��D���/�X�j
O����}phv����t��}��N|�!ܼ~�F�I3�ͥ�4��;v��w/����_���H�M��N���k����O���� ������73RhX,n�ZH6C[����P_i	���������j��J�/�A_�Vtu��������sp:��N�q�-�ՄPfHDS�z��4^�yU�Aڋd�0ό&43�pD4h�3�J/�
�<���1$�V9h����l6%��hk�.�4�����s�\81r���`~�m�0��w!g� �2�X�0̚�JI��:'���dL	���˅,�NL Sȋ�wk;�F�XY[�W.������l*�@���ېNn����а:;;e��̠XR�l!�J�&V���'�����R�Ѐ�P4�`A&lU���6/�"���ઐ_�ݡ��Z2����׏��x��=Xa�?�5�j�3�FL�l�>� ,�fQ�[�����
A�i�h�J!W��{���,�ceE�qKyS ���>�}�؈�*�BK4
G���o�sS��ґ]8���1������B(F�����w��oG��AD[Qbl�SC��	3�����?��09����{��L��-�}���H&0~	�K�x����Mivc�<��>|�P$�x�H&7%2� ��܊�---�<7��(��@ (feB夆�����Dꈙ�˺k]ńYd��r@.����EV�LVeT+�i
8�1חrN�g����s�}&J��k�l�F��v��75��͌<�̙�6� �ￔ9t?,������;��y����R1�!�&F��O��q�?��j.����F��h���>tl�Ok7��8��s�6�(d7��jغ��C�/xkl��ǀB	��B�M�3���%���!��*�B�{�W���-��?:+v�w>�P@�����È�s�38��Ǐ��&��̽�x<N��n"�ɋ��5�,N#�\�,��|�y��2���p���f��rB̲b��f��I8�~���₭hj���WǽCA6��ɓ8���㔏�� 0��GC.��+T���L�� %5*_����<4���Ke$*�� ���>�p���
B/eq��9\?�.23wľ_���J��w!�1OS\Mm�9�2J�Y�<2*T�<<N'>'ʦ�ia��]��u"�I��V�ژsL��JY��J��/�D2��fӡ�v�Y�(�����<'�t���L�zBV���*��y�V��6�8���AY}�J�9�t�7�a,.5J�zN�죌ekLqiB ��~}��4�������_�z�B��o���������l<٬ҹ���wUtkY�lA��A�����
������4U�&">ڂ\��m��Ϳ �@9Ez	�ɔ�͠�u|-}��[����r���&K��hn�a��^t���3k�pi3����04�.1��2���5x<~y�~��Cm��5ܝH����#Mx�� 6���=�@ W>�n�C�F\x4_��@K܍��2���Y���84�2/�C�Md�Q~�q*MI�O����Y��2��{��I����I��$dz+D���Z4�t�-S�Rw	�7�揅��>Hp�*�������1�fP��j�/�A��5`ai�K2��'�#��9D}6���V�����4�c ��@^p���8xh'�"���"�4e�67�Ѧ ��ۆ��BH���#�*M,���W��0q��4�M��|x�G��Y�w�=���!}ᅽh��b��._�)�ʾ}���@��S���;��p8�>;P6�,�_�$��rA���`p�	U��G�b��C���W�����3cb�]f.�Ր�u�6�66�%��h:����*�D�Y���w��c��r.hF6dstīB'��f��PR�*�-�D1��B����߫�����bsmk��Lό�f0�rb*��ڴ����ًP�vh�VT���
�n�`�����B�n�m࣓w��A�p��6<u�����g�p��=8<~	����Ã�4\����><	�iǫ�=��� .]�Ĺ��%��pI�8<��������@×��t����Č�l1 �QnOf�,�.x��� �����lE<��b-��)��-x��^�M`trV腅;�&�A�5.�����tbb����É���Œ4���Ba�H*����pIA�����RhWu�!�B��QU���lFBR��Ʃ �E����,�{��(�&z3�N#=��4Pb�N�shM�h�v��a�4�j/�jɢ�[�S�vc��v��N����wA�$��o�|��2�=u�!�]��Ӊ�RÀ�ه�.fe��ǑLm�+_�
��p��2�߼.Smn{���{;Q�[��o>��R
��9�g�����5\�6"4�r��q<���}�Xё�n!�"�r)#9zÃ]h�Zq��f�bǮ��L��N�HL�q&� r:��\i���r��IK5�\;�Ϫ�}�
�J��^��-�b���ܬ��l�`��V2�x��V���hR��fDw�F����KH���`?�Jsw�b|�4��F�����ܤ����S�#Ժ���(T5�X`9�p9�1�<���I��r����W��lFr%��FMU�n/���h�X���y�P��P,��v��R���s��L&�q��2)���i��w��t�6L�X�<u���ƲZ+�eT`�r��HgO����G�T��fníhg4��Z�aD��F���ˊyQ����?K�Xפ5>`&__G�H$�p�M��L��&��\+��/׀RAMaC(��Q�����k0lt��°�p�w?ţ�[x���x�?�-��/~�OD�GEW{��M�{��oB�B��gkEds�[J(��l�@դ��)&l��;6�ITIѳrJ��=�#�l��UE���^�y���U��iYE�"Pq�t8��t�����g��9]#�!p��,R�L�K��i8qe��x��ć��(�EM���YH6�L��5��V1�n�~`�g��Z�#O�kBY2\\�Ԡ$Ew8%\Z$0l8dJX�,����A�P�IKe����)��hsW��O�sqOً�����)���(�PGb[����=#�I�
�|�r^���4aɗ�M�a+W%�զY�/d0�1!����<�^�X�XO�Z�n�(30k�(�:ͥ�?g�f����F�R!��r���Y�,��|��1�@Q�Ea[g��.1���MA�H{;4�Sܞ�:����O��R8��c�(S��t�>�W�w���o���s�ש4�����dŴ����X������`@j�*cIt]JZ�A���]>�+���9`�K��FŢ��D�c������f��(C7H�d6�)ε�	b ��Q+��T�
�KM�-�A6^��YQ 0��h��g���Ny4q�%h�ڂ�TN�	*������S���x�q�QC�"Y�3%���w��%a0QG�k��.�ס4��l��#�Mk5qҤ>>��v[�#� dE���1'M(�[��8���J�#&n|]i���H#�ڐ}4���C�E���RQ�!.�x'�c �k�� eԄ����
_k��}p�[���&=�w��!���^A0������"�%�=Ls:��fX_O�5���2ű�σ�c ��bmmC�.��n$�P0���"p2�讃~��L�qm�"-�����5��/�)�E:�{,w�|��a�C�;ŋ���t
�

�24�#5�by��QM���C�3��O��.��]�S�J&�����'�M�_���p&��u
j�*���8��x]�B2�mVɻyd2�?J3H7Q���` VK�l��G���O����14�[0;�����z�x�޿��#�ph��v�[�;�o�iz���'2��sG�{w>�d\�,p�:���wo/�iΜ�HF�<��`7o�!�4�d�ʫNě�/^�T �&j��A�PF�okF�P���IY@[z�h~Ch�NO��"���+��Ylx�eñ�3v�DZ��2:@��Mn�\�D��J4�I
�I�Z�eD8}:bU�rE�����Im�u1������N��O��ǣ��H�ܭ7�˰#�Q�%�Z��=J3؂��>8i����+���+��pskr�9�=]&�q��8��]��i��Q�֎V<�D+��q�����r�r�.�ٓ�@�{��j���f���� 9t��3\6��t[\d��9��4;ں0���R��I�R6�g(���u���6�mo:�n�a	��VIF��V9Q��l��Z��h�+���^V�Nu�e�KB��p��"��qK���;��9D�(��8��*R\���a.,�g�p�l�cE�X	(����^��
&F�a��idF��C�L�YO�ꇳimC��F�D�ZA�Z�C/��[C��aKw��i�fڊw>���fJhX餶'�ɻ�8�y���/�D!1���z{��t���3Be~��ӈD]8s��Д���I"����v��ޅ��I1o�c|r� �/���n'�&\bb�V)�f-��S�E�V���B����)����D�T̼����z1*�A��s�MB�YP��_�hJ�AN=�U�nG$��Y��$c]�aI4 Ղ�rC%�CQ�,�8]p{�b䔩`���>��j��^>��ۗ�uai�>��ߺ�	���:�¤#Uyd8��l3b����g��y��֪���M��4j$S����P� �F����~��P�eizy9��␎�6k�� �k�{���%��HΠ���%V�%T+i��5�]����z�J�f݄��G=8W��z���d����^�����T�$����żXP���s{�zd�yd3y�sY��߶ȁ��5�*L+n��v
6kU��n�@og��>x�X����ލ�~�CW��o|gfG����K=�V��`uzQ$=��(�AS@�X���y������s)X�ynC�8�S���������W��T�������PZ �,¤�0��`�r�����G'��1�dP��Z�:���5i�f���o��ko��6}�N����J<�j ?���w�����9��rj���W*��?R�7�r����0�0�H��C�ID'8n�Ch�|-5���t��D1?y���PYy�g�=���Ņ�g(�Z}�zB��"�9 WS�PL��%S
b����1/���4G,ƭVt9�)���4D/��<��k�iC��O͡I�M�	u�n����'���e��YwOv�)�a�^��Բ���P���|�*�N�6�cN	<�����漮ͭX�v���������+�<?�*E/��\��w�IqS 8�4��[���g�^	[�4R�D.�������/&��&W�io*Rt�YtƢث�rN4����0ɐ4K=���ԉ��!�"���&X�:��jQ��t��A�EX sM�
LZ7AJ�$����96;��&Z��bQ�q6�lY����2���S[��h�D��!��Ä�lP6UN�z��zT}I�Z�~�f�}K�a��H]s��"�TY�2Ard�*���9��iD��d4���d����Q�&] P5�����M!'�&�Gּ*��*�4�L�y�C�m6�U��&�� .�8��o�H��QS�xUh�.X�-2�n�3�*�A2|C$B�̺J���u��*W�{�O��R���av6C��߼N��,�5�J6[4Ϫ�X*�fqX���祖g���wE�:�s��2�*lD��3���<���23�π�%�5<���
��XI�0V�L,��H�m���� ���N��ɓL����>c�~��*�?�l8�z\i��%�r%����Zd�,�kݛ	J�fJ�c;��Z��j������v����n&�):�h,��m[dA��B�@��f����ݻ�`3����*l�l)�e�������wwA��h�a���y�H|^?r�,�6U\��n$r[�J!T(f��Ȏ�-�i2��KӤ�qv
)hD�t�,A#-����85�t�v���G"�����8o*�T�Ϋ_5�{��r=8U�AEA��GD��PHn�V� e|�9��Bɓ�O�m��@�T*G�<�� ӂZc%o�F��)t���^��?@bzwo`��,�e��ڪY)�M��#-����vl�mF����%��p�a�����F7Bx8��R�&NZGN��%
,0"�BY�pc�A+��P.�:@d���L�X�1d7��I�kY��,�C�&�`�ͼ�d*�@$�L�(&� .M,(�0�6�Da��R)T*8=Vd
i�&�73�*�]�
����	����$(�fcCH��ž�Ǧh(j2�@�������2�=e�`!�ã,�5�˪�y3��,T�v�txr�i��Ã�t0t�ʸ;rn�F~i��,j�M�$,> w�64<�`�0��h���������K��]���g�.,�agh@�k��<)5�e�_�R-��g,�J�`�SLq����:lrx���J�tB���x�+T;�Y���H鴣P,�p�����8}"�X�f���EP\m��$MO�أR��M3�u�F���']ձ�s�^3(){$Z_�@���ވ��4��P ��&��fR�w91��~D�� �'���#�ƃ�u�������[�ൔ�|�.�]9���3B�M�<�����u�	d�'ڋx�6Tu?�5 _*�V����$��R**9�����LC9��N �"^+{�sDj
J�:    IDAT��I 7F�p�������,�ą�4��{�#�F�"��j]i]尩7|�U3ǚ�C�^$'�u*������g>+�H)��j ޢ&*�Z�S�}���A1��*0_?p��!�v�;���r9��s}�![%�n��/�L�E�)�W<D�Z�lm����Go�k����ˇ�_����귾���3�l�=��4�z�h[��#��U�Z��]��[��p����.j�T�y)�d-��,i��b��I,�}�j=�Z�"E�H�)��,n,�~�5�@�Y������bBTY} zܳUSY����礘����곟UO�h�?��|�<6�S�����g������������\A&a���:45E�5�d��40���F��`�Z)eQ"�_��T�<�^'���X��;?�T���̑�(2�|���P�.�~D:�aD;�
�a�A�%���Z�Y�Y`׹��V�Y&D�uN�U��i��r
Zh�|`P��G.�m	Ҋ>���R��0�4�SR'����>�K%�[��q�X�f��B����ıv+4�S��y����Hu����	_ݐ�?߫hΔ���Z�	l��!���Vj4��C8���B�g.���.]��:T��s��2~`��BaW,E����7!��p��e�~�W�̌*�b�E�gsb�C0B�p��p��p������f�,�M2؄��5�$E\�p�L�(Ey�v���O5��,�/�jy+��T�;6�P���ܑ�ǳ�����Zj��茯EXej�Gz�f�u^&��U�����xģ������z:8 ��*�C4���uƖH�3�D���$(�Lxuh�U��R��|T���@�h��YNisP��TIu&U
&�^/Z�~\��N�����0��r�ϬA�D��h�3�
�?�b�Nf4WrR7�%�P,P�f����D�'�N�Zl�>��"݇�М�D�pݑq��:A2W�z,
X!P̩#�k���Tl?�t���U��<��R��1'��xDf_�@N�)� ����Tg2�U��P9��M2������r�ֽ�s�?S�V~u���2�����3�g8)�eyf�&�C�A��1���%��f�TӚ��_�d�/�ty[a���v�D��4\R��HIri�}2J
Lww���pw�."Q���B�p����F�ARrp��ջ�ƍ?�T*QG�5�K6)�j�f�N5.gN$�������CV\X6�
����tRȉĪ��h}��)��d6�L�3���H���P�KP5���Q2�׫�����!�[q�̇�ҫ�o2�hn�|�x sBYa��b��E[B�h��Ux�
1�b���j	�S��� Vg��<1���[ؘ��%��V`-g�� N�zZ�����f��FI
�2R�5$SKBg	��0M�BN�J&�"��D��nE�q�P+aTkH'Ұ�tE+W�qt0�Ԋ�Y��Q,������/�n8\��j$�i8}^i�v	מ��m~���Ic:#Υ��^�TN��\AF��`���<�� �5�PF�&�\��=ڪ	�D�֋(6�lx���z2��n�Ad�u�$:B�5�n*d�P�7�N~�����[a���{�fn�Fae��,��Mbo�B|�>�&�"o����j��R^�
�t݅�?��E/�`�3p�D�"݃l���\V�c��brCԍ���)[r02�*�U&��eH���C��?��.�}����~�6:��Y�`������K�Zsm��sa�J++t�C(ڋ��L�)�Bo��~ﳼ4�K���y&��i
���^G �y朥�,,%e]53B���k�T�:�@��l���V���]�_>��WN��!��,����ch�U�Z�Qռȓ���Pf��!ج���x�ZOʔ�p2�K5S�?].�����b���oI��ɡ����&��jE*����'B
�^/9���<)���H 7�(cA��~�Wa8��^���"���"g7������n�Ãz���g?{��%�7@�Э����X�4�P"*{�E��I&�T��ppJm�e��AW4�'��f�^���;��*Ks�����M��r�fŵS�}���8�f٢	�Űi��������9���R�KӮ;=����z{�1%^{6���Ypo4�, ��������+���x�)w��և�ᦒ*�0�9reɭ����*��VZ=Jc�<
��l��>�7�+��c��qb>�{5�䴚�?\�B?�;��g���E�Bד�s9�M��X���'Y��H�,
�ȭ�ض�A݆��1��G���#<��\׮�(�8>�0|l;������AsќEqӕ�kE�2�!˃���|^�s�u#u�L�L����f��"?܆K���Nz�,��_>���9c|�|^tv�.�}r��W
���oI̙����2r�p���w��Pd��g��i5i�"o��!�\�F�D(������p5&��0po%M��^��)@IUH|y}TsX7�� V��?�(VL��<�Ŝ8��a&����<N���G��9�S�%�fp���[���h���+�F��R��	���'5Jk'�%���6}�'�Z|�VpbƆ��:�F$d�I�T��"k�p����#׮Ҵ�L�ul����)3'�r�U3(u,�.V4/�F���͠���*���P@��9�[	��V_�j�|��Ⱥ洑�O���D`3�kC ��<SR�y^<��)R+@�!a�Z,farZ+��,/+��z����G��7�Zz]�*�A�1:�����x� �t�G�t�?Ʈ��aQ)!_$��Mf`�'j���rxMx���b���\���{�^��d[��EY3܇��U@N���r�*`\]���\�Ru�`��=�[~�l�����o�����bv�v2�SK���YP<�������u N���r8d%�>��h��gy�����vX��fG�r ^�}8�$��3�;�`Yg�B�|����M��A6����.�fv�,�Io.�@541�F��L&1;�P�cҳ�u�J��)�6��ˁB1%�].�{,���faAz�,���yn�<���_�q�(�c�k����Y�\J�$7!N3�í�d���G�z���h�E.��0�u�ݍ�P��h�?�_+t[5�2���h�	��1��be���3��@6y���S.����;��[Q��d��縼nl۾���0z��F�� K>Kn�RZv�pE�G��چ@[?�p53D�)f��݁\.%X0Ѳ�7���PY>��׬.��քBA+��'?+���P�����
Qx>l�` �k�l
�A
�Т����N�ld
Yr`���>�1�[pr��CR�=쨘܌�~ N�Y��͢��DV�ɑ>�Q������B�`�º�$χ��R���ca���=�N��P�`�vp3����^x"��662X\Z�f�77�,dx ��a������WKb�=}�����$�P�&dr�������{;!o��C8thv���4)K���SM�(2��Y�;�F*�I�b!7j��.�o&dzA!?6h�x�>p�&����-�%8�&��z��3��ύ+�'�S�s������&8Rٸ	����U&��ps%x"Yeu���M��~`�&�_Y�
�U�lݙ��dfQtW|��?�s� �4�T-����%끍��~kr�K(y�z�-�yE	n4Wl�vn��V���(�.}���g��%�afR����ڍ\��;&.�p�n��9��%���9)���&5>bf�(@R��ȧ��S?��껬��|�5��WT��A��y/MyO�3M���	U�&O�X�dR��� ���&���q"NG;��L��S�7�HH��QgҶ�h�!��q!��51�5r
W�t�U���l��p���@TBcUq���Pd�a��I- _����ː�x��|�[�N�ŃO��o~{r��O�w'&a�е:p��U��#�=o�vo��"��,�b��2,�X�K��Uї	�������!o|( I9���_�<6�G�R� ͍��\�0P�D$���A�e�έL�#�Li�q�t�2ɑ)͆��>�Q�\����j�P��aQM�h����K�i�$�;w6��֩lt�c��;`�!��D�C��e���Nl��Z���I��G�7*����]�e7q���:o��ok�:���8Bwz�k��\;Ԇ	8��*N�0���ե)�}P���`I1��(d<�uj�����Z���+a"���Z�L�Wj�CM��O��h��v���R"�Vi�(��v�u(��i~J3-�Ou6��?<����_��4��Υ�kLe��FC�1|X8�:i]�(�/���~^��J��I�wq�T)h|&�UM�e+5+(P�*�l+��0v,����>|�HO�V�LN�x=-��.ĺ�a�FPs���a�I����dK(�|��P&��Ҕ��jRː{�Q�+�YF�P�Y�A:-=
%yf���d0s*%���>
,#=�+� !&�%�^?(�G�W2$b�S���hvU��:C�n�M �}�!Y�V�_�����<�}v���>��U$*�q�c��k���I�8��
7vl���7��'�Nb����4!!ԥ#I����}f��g������Xґ�f���_y��}���b�,�� ��{L�8K���7���~��Te� �����3$���Mf&�Κ���*���5�&�k�4���a=������z�-%	�`�k'�r�B~�9���J��J�rf���Ƞq��>�F� ��9H��=?��R���*�Q��:1:
��<���A_�x��A SE���\���GS�@��t��<ܓ��ɟ�����<{�xl��g@��OC���%|��я5��x$�0�~���}M�����G"����xn�=̈́]h�_7�x 0��r�0H�:8�>趈�J��O)i)2�����OV��O*��(���G6��`�	�97e���w1`�S�Q@$��\sJǗT2
W��x��j͛
�=�	����,Cw�2�C�M�V������m�7-� �8C�L.̶�4v�>=�nJ�20	pC����N��=Jx���}� L�� ~~v���j��N��`�C�y��F�Z�nw�JC:s��Vo]׭W^���WT#���'B�խyl�	CfX���fO�0��Dy8��A[еcg*�8�"�nՔ�2.&㈂<��=��uW�"��T��bP��.�&(�Hzg!g�J �Q�Q$��1�iy�a���=Ǝ0UТx�	�N��r4�-\���8"���@g�l�C�E�)���_���<@���d��lJƠ��;𹿵�:�2��S*�w��0�e��:Cc�4��C��ep�Bӱ��b:y�b���=�5�~�q��_wLH���>�e����Q��K�#w(R�����A�L*�۪c,"� ψ��.��4�&Խ@9h7}����,�߷�эQg+��A�?hvMO�wo��V�BuP���oµ)�y~��] g9�y�F�Fy����3�L���.���2n\@O�9a.qˡ�$�"�˸Ѭ{�H��D�+���s�E���bj��0y�U�.���:�Bk�vw ���{'�,=ݺ|Ng���V�=���������a9��왻Տ�Ȏ)�*k��S�Qvh�9[�.�zhP��5��bB��+���"���27@�N��ϓ����4�jy"L���(l�� �8�6�N�w�4�+hLׂ���M�!BП�z5������|a���a������@-�H)�9D��{�`���������:�[ߴOq"�sS�R���������7dRl������H9A�"���>��_}A�>�%}ǃ��˟����]����gz��y՚-��	=��*�ܮ��w*�/���)�)*��5�R����g���D��:�<�O ż�Pd�����!����ɟ����З{ث۰^8O9w�T��_�5�,�����z>��}���B00f���.o�W����;���?��R��׷ri��'��pn�i�f!��M=���_�@��� ����4f��г����\�RG�c��w����������z���X����z� �ōr|A��'K�uIې�5D��>��y/�gr�$①�i@9//�n�H(������z	����9���d��7}�4�Tf�K�� �i�X��p�G\
�l&��1~��"q�N0k:�72�B
���1Ⱦ�&.��AS��h��/����u&뷘�\�^s~r���Q3�8�8#���RC>+��C��4�통�4�խ�:}dN��e=�g����ה������c��=� ��Hg�pN��|����� ��i:M�둾���R�<0=��r�҄�l�',t�h�1{1S�&�=w��b�Ś����p�{��L]� G��H�'ge f��IX��]��]��	��N����ZR�kp�L����)�i�NeZʷ�rݨ�<��33@qcz8 S��f\�@P�Q��ؠ�7�[B#ծ�53:�S��z����/���ȶ"xyta2[)WRvxZ�ʔc�♂b鬁 ��ulL�=}��#��@�����L�y{e�Y�>���
����ĞZ�)��e����p2�l�U�_�UjjA�C�1��>&SO����rs>u��p"�	|�lMa��fj�6Ѝ���Ÿ����;02h�i�=�'
�@1e��%�10c�\7��� "PP��Lk����������(2�?яf��H�*/z2�L䔈q���v��HW$7C�epɳ�CSH�E��a׷��	d1�	C9�5ĞMM���D�o���m��< =��l	Ц�|f�\�t�L���% �� ��t$�C4��D�ÅhD)Ɂ�e�?L�<����þ����;������,���sـ�7}�F�a�Q�#�@)Η�x�������5�0���e-�M7/���ڊb����E�Š��ZR4���F��(7:����ٔ/ý��rK�msB4\ �S��iG�Q�~{G�Z̆��ID�<T����/��]�N]ʻ7*��y=�`�I��n�J�36�.S+׉;k�4���_�%�j��B�f=^+8�qY�3��5��sYL=t�X C@{xy�7�
�@�(T�g$jW���X�B�����\�A�3h6��6Q`�@D����2I��������rY���T�s#�TY�옆�ܡ��)[���)��-%zi�\|&�;��Q0F5T,�2������`&��t��Z=�iA�o��a�L��U�8=4^澳_m�5��D��0����E�.��p��[W&�K*��M+�)��Bx�l�hHmN@A�8����eG6h>������ v�X�i�C\�b�����aBX��vp�cJ�nL o��q��^��OXG�4\N����'��ym]{MSc���έ�J���؉�5<�����oTmV�+ku}���P������L�(��dm-`�q��j�D�@[� z�	Hpd�3	lv���a�\r�2kЎkj
ϝw�ˡm����0���7�+�h@�|}k[B�cq�t5L��n�}������d �g��-������	���d��
���І�lc�`��1�5IL���9m�N�$���ȴ���Q���	z�XԱ/��%�}�1-^|U���o��Ư���������͝-����H�K7�=�����i�s�|��'���t�Q\���ڽ�
%�q�db�U��y2d_ �:�G�Ш����ý�5@J4lP���d��1I]�,��F��y/jL�} 0=�!�H��a�鼧����k�M\x��=�JŽ��(Tޠ�t-_#~׍��C���=Ew�N���_G*�6����.�wI_*�]�՛M����|���$�	��.���Իz�2ю>�SwkI�>p������}--��\��W27�{��m*��hqyS��Õ��5�
��0'6 �"��@�    IDAT��kt�&����^I��B�b ��>(l�e��2e�}���0�Z�)�8�v�aP*�X��a�;5k�q�d2���g;�P�։��k*���ș$���t�ƙN?����r�c-4��;Ҕ�<-�y�"�%mO���d�P5Lt�dN��z�+(�|v�Y&�Q�3�$mK>*%�*f�j�����P^�7��c_�������=��%��t��7�42�f7��l^�8�f=!;���`r9���T\�9�"c�h �]��|��8'�Lp[Du�h�:�j��ӚN�!Y�i-,  g衟�a3͟g:ɹ8�7�sˊ���hb�D�¶�+ji�U5��w�8���B��T��d�9�|F@�PP��y�n.���m�烃`��h�nd���l�nA���78�D5M.#�@�f-¾�4�:25��RA^zN�yL�־��!�$S�f�JG��VrhX�xZ�H̍���@4ć?��m����E������}:�q��������O�����xjX���l� ���4rAv�~vַ*@�P� '@ؿ xب��>w�ݭ���]�I�~f0Q�Z%�
k��;p/4؇���a���H-���
������e�i�9`�a/1��A�J�;��?�Y�Ξ�)lմ0YVd���ǲ�*�̩��d�IC�X��X�'�`����F��	�a&4|}Ƥ4���$ݱR|2bE�P+�� �: E�Pi�ds�ƫ݊�B3�D�����8��`=O��k�����?mO�~L�x0à��y���Px���2����	?HW��)>l|���*�����/�d:��#��T��=t遲`�h�J0��Z9���f��ZE��򕋺��K�__U
D��#�knCєT�<����hh|F;�������t	��~7�Ib���B��hg?8/6���A�٥����n+c��Wϴx��|7;��ܘ�9��.��h�@��&�̸9p�M#�ei��}Ę�Ā8fF硛kཅ�R�¹����-��U*}�ab�K�qr��恵�Q""( �4�����]�C��߅�W*��e�Z�z�@���d�g�d+ ��I
�#.Y�_��ё�&'���uK�>���ׯ*��Sw{]=�XbYE2�*͝RvtV�����7=|ј�ź.�K��ݬܠ�X7���R.�����EEhw44�SӅhyޠ�|�L8���`�d}���4��my���T����Nғ.O�)��E�׍'���������O�3T�Â�	�7�>��o쭠
�ns���iko&�����??<��g��4R.jogS���*������^|^��U��v�%��}QCǏ��Gޡ���>G{�)��M*�����.�ȏ�9}��������r��d.�g(�3�+�E0�A�D�sn���!�<4M7͜5�9{sm��M��:���H� ����)O*mTp)Pd��8�Q�G�T1u����K�ANŹ�W�7�V�Iޡ$�L�S�����՗3��- ��hR)`h����<d}Fq���7%��)�����aLk�7���&���I�:SW�>�h���wH��~V��m}���\g_=���]�����=�w�M;-�CS��9�B Eۜ0p�����(�l"X��_D����A�gZ4����>͙���ýý�>.���45�QHд�2�=��g�B}���{q΢k�=0�9G5L�`���'��I�������v`u��ϼ@+��	���b��`�u�9:#L����8� 8��aS�Ex.���Z�`bB���p}e��L����HŬ��E��ɉQM�c�n����ϕ�T*嵽��vk{�N��\Y�Nܡ�ʄv�X���B�;���Ď)Q�OS�:MUwwU��[ʹ�.v�7�%s�5+b^w ��vS�[�j�Օ*��]���LN�ժ��&�&=ybo�r�S3ݺ����A&Z sL���C��X�~���j���6���=Z+g=p��%a�6D��
�?�&, ��c�`q��TJmt��G����0i�+�L٘��L]�n�Sk����/f�p�5G��u�=ڪmkem9P��M5��s�_�����5m\|E�r ����Q��7��̜f�پyy��s�*�W�5 ^nBS�з:����(�v�%+.�$܅�w�5���+��4i�9gyG0\�O�?��\��	�.^�46�n']7ev��!� Ga	�P����w�a���M�z4b�����,��,okk�	�|����*n��M�b83�jݡԪ7�BaM�nb� B 2R�`�cFQ,�F� D�Ȥ�.��/������_���u��I1����_ &��!M.�P�P�>�Ci�!���6�]b��0x�nbJ].��L��@�كY-���F�Aޡ����F�̲7`4��g@D�H�h��}���i��r�C@�n�4bAvDN�ᆜ�/�>ӑc1�5�@4�4޻�{~��!��*�w,�h��ym����H�xO��n�M4�^u�@���t�:��#1S6C�o"f�]X
�mS+���t��b:���������I��0:慤�&��s��j�B�� �QT�	�@o��@�	$�H�S�#jz�X����e'=�%ry��K�(֔��"��Eqi���h}�"jzB:��E��#@h�g�|@pp���8 .�Hr<�\�0����/��Ѩ�]�A����V���q�5��H�ODj��0������`]���d|bB��/^��������R����R�j�L\��e͟�S��YmU���A4��(��:ȶՈ*�][S1Q���"�e-�k�ư����b=��bh�*,2rɸ�JŒ���v�ִ��僨�#�3�M��V[�R)��p���ASA�6���r8L��V�e�LO7�@�q3��b(��8�^�&��g�H�Ns���*&���QzӇl�O���1yb�J�Mi�c�a(�Ac�(h�L6��.��A����4�B>��PJ�;˺u������#l�(��	Uf���,h�F�IB�t^͝�
�� �,h"@����V�7\X`�@f�H4�Yݐ�zMS��`o���=�rV"�v ~���.��7�S���zc'Џp�0�
��i��E���>�i>�&�I$ 
!��.����˅l��n �]�����*���B���r�YS�ⶉn4��M�a��s�Bl�h��%4M�B�߱54��4=KW�3dsiUFZ�kg����R�[�O=����&�.軿�{577�/���翨�����������|�b��{����'u��U]�|��
����T�{�p�CEKd�o�?�T��A�bt�������q�S�z¾�uph�b��@�VۯkiqQ��uEsyOd�[!w��D��C��ϭ��e>�Zm��#%��tI"+r�@�A���g�����N�,����L�^�1���l��hY�����أyOB�M��oa�0�h�B�1��ɘ�6-�זt��1}�GD��_���6W�o��G�G��Sm�W������N/]���tV;�55�me`�0�6m��l!�V����-���PQ�&�%�Ր�#��RT��p�e"c���I��I��m7@�L�9}������l:@8�j05�D��IAǙ��$�O �x���c�뮭m�A�%C�WhB;^� ~eP��s�����2����&��3㵸���Bu�2�&���%:r����͛��r���ꚋ�|P�_��k7t��q5�7�SS���۴����7_�C�Uo��>���������]_��g�ytfBo��v�=���x�	�OϘJ�g�������ܭ?��?���/��]orh��_{L�RIã� ЀU�p�nkw�yj�tJ��/*�/��=���Im1٬z+�$�0�_��1uM$����+����H�s�>[��g�9�Jem�8{d��0�[����3\^Y��W�iVT����G�.Z)���#/�;�[�n����V4]�m��!FJ�FK�S���&�:z�'� m��{�����Ą��W��2:�㷝ԥ��kucU'O����v��T��݄B9�����bkc����Ԥ��'5Z��#?�s����?���빗^�s�?��'O��[��ϟU֌�%�C�Q!����F�`�T;�LϪ�����)ڥ�VV�U,�T�L&C0x�13�=����;�������Z���:�@�C_���Y���.]R&��#�<���q�Yi��A0L��~��iu;���.n--juu�[\8c*�J5`q񦮽~��;����9l����&M�e_q�����*g��&�
��{���>�Fk�@q�U9��+�Ʒ"gF��ڢ�=�w�ŗJ����<�l���~y�����A���Ɠ>G���v��Z��������&@�F�%
j��i��e��ܑ9UJE�d6�~"�ŕu�zQM��k��ҕ�L��9�&k����g�qqN..�h}m]w�u���-n� �	�u{���С��ܱ�
�
ϊ{l�����u����W��0������-��Y3H��� ��0���P�C΄٩I�#� )�?i�1A.�Ӏ'�����ى�摷�I5�����)�/*��e��_ח=��7�'�Y�@��4��O���Ġ�p�m��a4i�Fh��|+���O�#�&gO�VG��8�6������c�0	 �d��t�A�t��{��Ԇ�2�����t6m�ba��+��X�J9rD`���ν#đ��C����!E�#�(��1�A{Glj��V�V��/Я����v�|FF���tB,��ִ��n3�@�y�As�:l��و�(�g����P�0Ha��(����3��T,���'#�c�����֊.�����6�f�Pm*�y��_��ixlF�ʄ`e�3͏�[;�^�4ZR9��TY�\��n��7=���Y�ln���9pߓ�8�]"����]�b�@�j6�s��wTH<y�����P���@����g2~[[�q�g��;��w�]ʖ�az��=��m�C�Z�8�[O�h��W���"Д�}L>�)]���Y3 ��`�q4}���o�)Bq��j�S Md�&����B��a��Q3�CKl�;O\�Fr'Ǧ|`Uk[�ڼ�Hw_�hS�=��F�X����Ff�hhtJ�.�x��ߩ)��9��Zw��8�߱�)m��9G���F�"�w7<4D���Ȑ���<$�h�y�O2i�0���׈U�4��҅������@�Mqy��yD¾�:~rr�T΀�"n����ycmĴC�E����?R��K�D�K�g��T�՘I�'Y�\J:�F&���"L���x>4T��}7��XA��P��y�3%c�,Q��HAc)iw{E׮���JN񃆵��sS��XSi����[��k��M}�Q����>�?�����XT�4l�,�R�s�@����J�]��� T�0^h6$�Z%�\ꕊJc����fr�V�哳�>L�z��66�u��M����eu�L����:�.s�ɣ���Z7�F�`Zu�gN$mNs�N*�?�x
4����C͢��H�+���1�`����	�� b����EL��<2Y�rY밬���lzշqU��A;�;c2@�f]o{���'��~�g>�+/�~�W�O��������O����7PK�M]���t/�{[]��	3E:=�l���lx�h���W/{12:�F�@�=\y��A|O�Qխ[���ٳ*���0��g�Pt�0yp���d\Z^ұ��t�}��,"��ŋ�����Ԕ5x�  �0�Y^]����͙\��Mi|�����nffz �h��+/멧�Rms��\��� �� �-|4h����^#w>𐎝8��_z�{����뱯>�ѱ1=��#z��U�={Vw�s��C���9ML��{��{��G��/���o�_;��z��KZ���;���^~�y=�ܓ�{������-�is������~����=�N�>������k�/���W4w�����6���?��N�ҟ}����/���N%cI=��ו�4;?�K�n���v�9��+�473��RYg�֎�o}�A���jmm� "��0_<�&�@�5�Hi}uY�.^�{������~��7b|�W״�����Z�X׭[��ĳ����i�i
��C�ߗs��g�ҥ�^2����s����d�<Z|$2-p�:~�]�g�gt��������ܬ1.]�d����]�.��k��u��);z�M��ڪ]���������ָ���]92\�o�_�����~�CZ�vE��;���~���ʟ|Jg�|�R����+�ʪ�hh��	�yϝ��]ȩ��Y$��_����c��s�|���fg������/٭P�������Vo\�Աc:v�zD& A�Y�${�e�g ����K/�6����n�O�x���jTj�z�^n�I��Duqq�a�������ƦL�@M���'G=�y����7����nC�I�[Lix�tD�L:`Ӝ��u����_#�vw����3?k�� ��7n�HG�L��ReDS��f�ݸz1���!OՉZ�dW[�>�����}Z?��~I/���~��EKK��?�3�����-ڂ:����Z�ٻ�������ϩQ�jf|\�x\��;���F]wn�ϡ`\c�5<>�k7�⹗Mi=s�L`�a^��l�s6��c"��.]���W���|�����|��xKS�vHg��邁H�_�i�,�����00L���6������f�a�/���׮oO���|tg[�Fo~�JE���:K�{��r��T�3{gg��ށ:�z���L
���d�"�A-�'��x2���wNh���'?��^x��RC�0��Wj���;�c������z�O����x4��I�b%����?��U�S,�v���QO���5?�RgЄEi�c�����@45àz\⫫K�a��\�4;p���5�٣}Bt����H���0:㬶�S�p����z;w��� �lv�A[؃�b��-��C�2c��|ܺ��������&�v*���b�شP�vPy���y�LHhH(@AǠ���Ώ�/��y"h�dȊ�����
q�L�@hw֗��t�}>�T��P��e&��UP(vL7�Fȁ������͆J�aeSE{m���{��w��>���������\o������<�Z�V��P6�V�P��֦5�š����NS�*t &�5�R���\�X+�z��kwW�>�5]�|Q=
�d\��&yKŁN��6p�nLu�jSSS���w�yki�!�
�-C��u�Z�+K�:M�M�1a��h y� d�ھ굦�_
����7�&2��r��u�5�><��L�L)V2��f����B�w�G��C�<nc�GK�X�{�)`S�bB���v6�u���onYX�w��t��{t��m�X_ץ�Wtߛޢ˗.����z��UA���g>�����MhsgW�S1�����n�yE�}mn��ʭ�)A@�iS&��^b`U���ٳF~��T_cS.�� ��e��a���g���u����D�f�ꕫFĠ�����]�ݕJ�M4M,`�u��PgVb>
=��:ἁ;�2�¹�� ⥁A���#>G:�ra�$�B�Z�iff�����v�,*�h��Q)W�VB�{;�'��?�\Щ��(�]oЎ�_��絵��_����?��?�+.�>�)}�ׯ��������*��.T�a"_#���aRI�K���	��4i������<����:~�	��Z���3׷����C�	���[KN����s$��~G��W��+�vs�@QM��c�6��6u���&6�q�K<���6		�{���F���`������ۂ2K�h�I9�}0`����p�ŕ(=a�D d{K��$����9���(Z-���C���~T��֫�������ֳ/����_V�T�[z����Э�-�|(h7�J��B&��[7������A�KW.��tdt�kVM���8't��5=��/*77��>���D�bb0'�xs]����M�/g    IDAT2����쌟���˵��t��QMLL��+紳���ͫnT��4=5cë���R�s���vLS��ׯ\ҥK�ss�-L�CN�7�]<�O&���6�sc�������smeU��/{z|��mn�����������.�������W�Z]Qf��TW��M%�
�����ʢZ[���?�1���~D��:�������W������oJ�es8�pD�K����=q��7�5���435��Ͻ��޾n�][k��_ZTlxL�#�Z_[v�9q�6v6�Y_���e�9�^���Ȱ���wjxlT����Vk*<�5(3�zZ|p���e-]<︫���͝]E�'�u{۱��n����v��}����nm_����V���⅋��T*U����ƈ&z����^9��k�n��t���@�P/���'�TF|��v�nܸ����1�յ����ڪյ�����9U*eSL91���X��֦榧���{)��_�+E��_?�������_|A�^8�?�������˫4<����5:5����U
�w��������T�8�J/����7+�B��3Dz�����ΖN����@��[�A�i�W_��D&�o�;̖�0����>�^!K��Y1X����~{�2�
C�)� ����3	��z�٧��Ohgc��>@7��P`Kq�#��gk����#�.��o��܂�ww����J	���G�4��:�8�:�ˎ<����U�^Uuw���M15n�@�MG��=�����{�3?��z���د����7������"(@�%+�h	 ��ېi� N�_{Uc����~��Z� v<-���s���Ä}��e=��36���7��t�����:����q�` s`��U�뻿[?�C?d�����6�6�P�\?�1�d�n��Ly[�A;�;���
��nܼ�G}L�^=hnm�U:��.�b����N�s�������A��Vi|�kB�!� ��|���4��ڼ�XY)2��1T)�ȉ)������|C�.�P�H']y�o�;4�|I+RCT�@G|h���2O*�E<�x����_�p��O+](9\���Ei�l�)����1y\�<��`��AG׎I�YmU�][��A�h���{O�S�z��n���%��'N.�e�ʵK��:y�:L�Z���O;h�	�M��;8F��=�^Jz��g�!h��F֣rr�l�� �:��[��[��#Z_��].�\.�ݩX�����.y��p_��9h -�\a��ͦ	ݶn�\T���"��>L�,/q40��i��g:옲��Q&�P�����rٔ�Fi���z��o_U�1����t��ۥ��^{�i��������������~�c����z�;�[��Oy�ۉ�B3��XP�C��+�Mج���f"�!��D�8��nUG�������DW�#.о�տ���}��횊`޴O�8 ��=D�t��`�ԑ��\�lln�`�S!�L�L�q뺭�O�:a�����B�BC�͸���z�tQ/^ҹs/ikm#8�؍|�50�4Av��v�WsoO�ʘ�t�}�@uTQ��m��bQ�w,T���L������=�����-�ljiyMc#:�pL;k�Z�v]���ן��g���տ��O)���#?�o��t��o���5>3��pQk뫦��/.�uc冲��P�C�0�T"����;����/}I�׮��Bg5:3�	���vh�H!��R�(=�3�F�O����4jz�s?~���ҫW��q�j�`��/ho�U
].ThXЭ���&(誛��o<�=��3������}-�C�� � �*B�ѩ	MMOilbLW�\1�iltB�V�Yn�lޗ;�f�����'@/]R�YWynJ�V]�W/kdvN#���õ�[��\�ܱ9}�㿧���驯>��~���I��;��T� V,_P?������l���QWk��>4p_�EҘ4}n�|��ֿ0���@wӍ������w�C��#��������	����+�5������VW���UWus��'��S�XLI��=��b� �.�NG�b1P��g�2�)�X����(��]���6M?h��8CVY�<1���*��jzrJ]4��a2o��*gtR�rEu�hd6Zc�0XA1�:\__u6V.�ٵL񋅼�·��^������ޫk7��ӟ��"�o����Գ�i�2�bqL7V�t��kh�bJ�crtL�c��z�Z�����2��6wwL=.J.�(��~�V��46:�z���/��c�ܣ�'�yj������ۼ���W��.P�6�|fM���y�p1�C_�u=6�3L Ǵ��������Z�����[7����x��W<�E�������[��\�ħ����P�w�s'M�Z4��#Q�m��;��N�y�]�us�?�>w��������@{ʏUL�������[�om)K���������������o���y=��C����K_��ξpVO�q�T�d|��J#����֖��]M�������^8��fM<���G��C��֫J��dln�X��V:�������s���{ߤSgN�����i7�\�}`��_��7�����?�}o�� 2�WL� 2aw��%�'�8"��N)�E��c|tD��]�llh��q�{��� c_�~����>3 �B(w�2q2�6Cnl�V�R��{��C>l��Il�e��y�����X�##EkɈeh4:6�`}�Da?A��N�Cn�@Ǐ�}o>���ο���%�������:����YYS������q���Q���B����ڻ-m2��g�-]C�g���x�k��8���2U�ҟ~��z����N|����1���������sO���f�����=zྷء2��MK�9@w�O L&�L�J�%�ڙ8�W4gL~\���}U����K/�٧�1 ɻ�iG��{*T]!�A:"�f�55=c'���Ds3���5���F���5�)ery�ך�7��v����m�l�B��轋3��V{��;����ݼyC��V�����F+#�X^�.� U��� � ���pF'i7ZX���a�r<I�������k��.��jr|���R>�n�����b��`	��v�.^����p�����w{�M� ��~)���/�\;f!�+ ��+�G��6�\4T	�~���|������3�nC�t�k�LjC����iMN��ԩcb���*����r�|�1v~Kј��bl|ܬ��yL���	�&V*��-�Y�7׻z���lt���`(g�h`����`�b��yG����h�IY�Ĥ\�����>ܯ��v�ۯ6�0uv�ց�t�x��rل7�#\"YP��=)�ǡ�T-"�����Ƈ�����3����H���c3g��-�y��>�Õ�;0�)r��2eUFƵ[���l��ς�D�$���_������I&X��Y�������@C�.�Q��JqT�c�j�AH1b�$.��̤/nU���bD�s��$Q� �G�����(���'��Z���fk@7>�{���3)���P:��k��Ĕf��!�Dլ�)�%��>{��I,���x�-�����m+Ú�P}��W�}JSS���y=�_ԯ�ʯ�'~�u����������!5��JF���w�W"XfM���P<A�<��}&Hh҂f����)k�o���j���ʄ�W^{U��ʖ�J���Wy�l�|�);x��x6v3l��t�f��t��Q2�{�ps6�]J��wz��5/���i��nissS�F�p��/�
v��%;Ù�_xN[�늧qˤ	�:��fS!�=5�⳶�n�rzf����l+|�r��!�a
�Vݗ\�[�ԹR�i}s]�3�ګ�� �z��^�+Z�ݚ������������}���~]?��?���>�_����4��PQ[[�*��(W�ieuŔ煙���SZ�ܴ�E���� �:@�f X��g��P��c_{L{������*��=6��"�#_Ӕ�Y���|�����5���z�@��n�Ea��)�իW�La����i-��n���T�Eu��o��!��SOy�A�gj��5I���$\���ƒj���� �o}�~7��JI7o�R�I k}���)}���nO�BY�tA�;{:��YR���ٱ1u�5�1��hl��#G����w�?��ʋ/�7�w5R���/����&7���$��j�^�c�i�����D�6zI¦��@;�BLO\S«ׯ�?�I�E�{�}���ΖVW�T�fܠ���<�Ԃ�@'s�w(�!��n�i ��)�A����g�'7o�0���@�D�܌ �om���og˅�Đ����-L��4�4���mߦ����3��$�&����z�?w�h�=�A%}�;K�T�����n�D�5��SvWJ.���U)����������G��;�+�^ӭ�U�L�)�����CY�kժ��M�������仨kƾ�AhL�+5?M�a�g���?��}��UmgK�����6�YÚ��Ķ��D/Lty'.\Љ�'��~�L����4��Dޤ'���m'Z�HO�rٓ����)��eιkpύ�^��e����W��%�j�V��3�qO�����w vݮ7��}��;,QM]�.�j�P1pH1�&=�Ij�U�~}_��iR�BA+���J�����n����qmo�\&a���.�~�W�f���Q=��CZ]Z��	��8g�������G��+d���V�U7)���6ַ,���G&�آ�]�c��S7|�Ͽ�o<�#�g�C�o;c=w?Mt��  #mg{W�K*�2���q�hk�z*p�ZELnxf^Lz��O&5:2���� `K�� �?��;��Sd�z���1���hk�ġه���!��͙�o��>b�������xp�HjÔ�k6��gē
�=#�em��x��n�R6@���'��Az%S����O�,��w<�J)o)�骜ƽ>�kK+:�d���V$�R<���̘�._�Ջ�596��uuu�2�B������wT)�XfF:y�ξrN�}�q��i���o��#'�0s$��f���uq�Ν}Qš���5����L��G-�~D���i��;�"�>Jw�������uyq��R�0�Ĵhl��A�#����IPyl�S�D,���X0Vb��m���������>���Y'�� �ad����i�{��N0�j����Q���	�	��@�W���[K� 	U���Ȩ��,	 ��2��a��3Q�����t�n4�ԯ��0y��k���7���<2;���RtDu��B�F,H�g���^�9C�f�]�-�>
�����8�!���g����y����
���������U׺�d���`>�f���ۍ)�-j�4���q�8dU�
9��߂�"��f�$!��_0�X�N�f�1���m�}0�_@���KƵW?�����$�&���!�)���?���Q>8GCUC�hD�t����7{\�dv|��/3�Ü'� |8,�C�yP ,��wΒ�Q_����Ka�G>�Q�qۘ~�_�G��{�p�'���5�as�l8b�.��(����.�/jckǗ�0�F��ܰ�W�z���T��qp3_�K�X*[T���O����@9�4g�ft����49�B6���tu�zpk
�����R�����4E"�@���}�Y�l�頁�J�<49���̘��&��}=���)7A[�l�W7�<c8��m `�a�S��= �g���B�
��3>:?��O������C}�C?�|���_1w�t��ƠWn�VMCKe�T�T3E4f$�Z�S������3LFiw�\m�ML�����O$:Q�R�}fnֺ2�� h�M%���!� ��N�����Pa��2�57���!@�Es�������; �������#�;SI4h_�җt��Uo^�It����!a��#�:a��0S�ryD���SǎS�У��=B�bɍ�l{獵O P�Z�+�<#�gn����'�A��F�{*��?��g�G��;���a���}��^ٴk��ʊ�C��1��F(02<nG`
..��8�9dٱ~Y�4C�H%8��>����W_q���	����޾y�!DZ�K0%��	�۸Ц�z���~F�&R.M
�{���.��\�K��99=�ÚK���PA[[+>C	�r��?�����c�~�Ψ�H���aJ��0��nM�REo�a������nRp�������v ����ّܼ�պ���lvU(��LE����޴h~ft\�������Ԅ������o�~��Ԭ�����=z�#�a��SШ���+;*��*��:�*�.�=3��6k����-9C�.��d�7~�7u��u�����n�|aJ�k۹���:�t�{ss}C�##:y��_�C���g�����+yh@�����
�^�TydئL$�l��q9�\^�˯��K��B������������h�hDoy����|�.���µ	��{��[�̇��Ĥ	0�l$�l@����'U���fv�]SZ[Y��Ϻ�x,�*�+��������5U,���%
y���L��|�v��Z l`h�/ܫ�׍��`C��sB��g|���wq~��1��;�����z\�M%1��u�ᦍ��F�5�v5:=��M����3�}UF�>�766X��O�i�����_���N���� �0�ཅ��P腬�AJ�m`��yg�gt���L�6c	�I�o�[����T�f��Rqlع��fM[�+���Qmk��X��Z��^���؈���kW��e�G���Dۋ{��Ҳ���PI�^D��	�&�l�UH�igu�`N��
(渚bN��$kQ8�.��\��ވi"]I&��D�t���6�Z�y+��!s�����BL8
�٧��������NؘJ����Q�|/�^�P� �.��=�^2�\e���wh��ִ��=���;���D3G�������/�*��Bo�d��f��;���Ԏ�U��5�@M4??�W_~Y˯��H���{^Q��U��xfU?�t������(�y��RqX�ZKm"�0Z��Ra|T��aM��=���\UZ�>%����{�;�P�`�я�4��i^��>A-�Չ��u�ɓ��g�I�&�ۙ�Ce��������'h�6��g�1����B�x0���a2Q
��!+�ô�����������ѹɤ���5wd��X�<�T����ks}��9�yx�� /��)dŕש�w)[�X�����]� }�4��#�uLՆ
�؏�{�ډ�����ͥ[�x�-�k��I����29mlnjkc#� ��:�đQ'0�pq��6�c��X�I)�L��~�C�s��::=�~��f��DO*$3j�ה�g��h�Q��_����b8R��Z<a�i<Ya���d�c��z+�O��GTY���k��H3HZE4Y��ԂFƦ܀;�cw��z(�t�~7����eT��	���8L��tϽ�m����=��Y�g9�}Lf8���y*(�/���?�m8� ��&z����-���� �����F�e28�7~���{3��0m'X�ڙ�g���*�np4c1�hl��L,���JA���|P��}\��x�A��Ѱ��hZ.�����&�Kf�|�$�ЌAe�!���ߍ��y*��O|R[��J沾@0�6�+�@�ĘB@4Cx����N�9c|�v�!t=$c־v���m[�ǆ
N]���2���Tp8O�OhmcC�}�k��XQ:�E����򔅦���t�оf��u��wiaᘲ82v�Z\�aMC:�vՍ7�
��ֺF&ƽ��9ԡ{P�3�&��l�^��L���Q�9-�,ꙧ�ԥ�^�>���}���R�[.�*ã>�v�u��S��>��"&�]6�v(���p�UбA�4��_<wV�ξd
k�\����qc �A�4A�8H=Ёn���/���7L�9�������K��(�~�(SBg(|Y#4'����/�ɧ���ġ E����u�ms    IDATs7�\��ۙ-S{�i4S�;Nߩ��q:��4��Mg1b���ܲ�'�d�|Y�T�
���nK{�+���X�;���i̇+bq���U�OM��{�����ˍ�Uk s��TK������3bogC���?W�X���6�i2E����
H4��K�JK�ҝ����F�@�GQ�L)V;�P�j��I��f�Lb��$2�φ7�E[Y����ɓ�2�>a�3����rs��ݑ}�E�̭`U��u"2��!_p-�A���x��I�vK���pӃbĴ�����"I�U�R���$/�@�V�Syޙ}�TLoZ�AƘ-�180:�� M��ՃRגP�PR�PQ:_t�{�i�ƚ;�&�Ԯ��erT}&�4G|�0�f����1��ܜΜ9���iժ;� �8�l���U(�.�����ZY\
a��g����r��x(Y���������!�5g�p�y�%2iS˹/<���3}K �\4Pq4������֍�M���n[�c;�c�7ݨ����+�[����]9/1Yc��:�D�B�U
4���� $@ۿ��e�6;�	��&�%J���?��Ąi��TJ[�Kj@�v��gx��� ��*��� d�fGe�� ���irvJ��{�N�v�@�⽘g2ܨ��E9=���wu��M�~@BP�QĆphd�������������`J;s�p$NX_X��y4ԘT ���q�4i/�;J����0�Y9X�����]褜^/��h���Ĉ��!��d~&��S_W�gM�*1�!߱�H�TB���5��cuM��H:u\������ƏUr���1V,�ŧ�Pks��=�e�MKL��){����g	�����B�,�Z� $�>}��@�������q�D<������h��ڳ�xo6�@b���yIcFA�!��?�t��1���#
c��F�¬�m�g����Ո�ť܁�m{z�ĺ8^�W�١�Ӱ��ie��bbn�6��Ǟ���+:�٣ǵqM?����E�@���@���*k�a�S���9�M�4t���&�5:9���q����u����lm��p��q>�u؁R�|HkA��
�s�;ʧS:ytA��u�����.�8�����!�(gI��O�{�ZC�M`���8�?`PO��q�bNf��3�;j7�Mo��q��z�A��13�JjxfF�ϜRyd�zӛ�o*��if|A�7W<���R,dԬ��I,`��a�������Î��F���%�p�d� 7�� ���q��pD8H�g��icuE˗/LGbE-9~��u����a�Z_Q����&�f@���!��QP4.|��4� �I���NY��Ę���5gr6V�e�DAW�0%�C��ɘ�O�����|�@I����s��ACF>,ң�M&C��h���=�5����oz�2���7y�� jc�iZ*�y�FH��Vw_�dΜ�o�Ӡxm|�8{6D��fr�wG�@�4����7���ط$�1P��ȁ�&��$>M�Ɯ;��p70� r/����"��#�N/��Ķ�\���Άfp �4Ip���hb@3X�I��9�M��=-�8��ኒDE�����8T�[n�8$,�A8ۥ�j�q�GG�6���6�+�&�?/��&34d��k�{2w~(�ɉ	���}�)���bC4Rȉy��s�m�El���p�
F� �x���z./�׮�T��:������)G�7nت:����aφc����W&��R'AQ�TF��<�t�6Ams���k���EC�2<1fD�*Z.T�4.$�����Pi�D0Qds�{�Ԃ�R6���K��yC1cA�KD�j�̽�.�|��sF|x�,L�A�1Bz6,�����M#��/^���)�8~�S�T4�.t4���{�4�7�_���k~�|&P�؈��/��G�����b�e����X�9ԡ��`�X�����RdAe�΁�"�M�֬y����P�(�ތ�1�궘n����]�`:�UᒌfK]�'	�?6S̙�of�s����s�Y��	���4�P"�%%uP�*14b.;&�g��+�@�qEXݨ[ו.-zvAnm�h/d�n�����$�i�*����FH4
��9&Kkk�E�(����:�Lh����� ��p��f�,�����sYSuA�Y��|fn_|&.,�A.f�@"�V
v���ȡCSQ�GeXO	�[���ybZ�T�t�f����:��n�h�xh.~{5a^�V��	�\R
6�c?Pԍ�rPgˊ�*�[��`�I�5 �)0���,��������|�1�3�;���)W(��;rt^Ǐ���nu0��f���qC�����3 7ލ�QmW�LGG#{<P�:t]��4�l�����衿���2z;(�Cf,�5�'vg����AOh��Ɏi'~�N�}B�Of�m���519럛�9����b�\#�\�T�D��$HY��<��27�=p@��>l��9W�gT��U���4��[�]]���&gߜz:S՗&@�(y�e0=���=55=m�. �]f����b^=2V)����`[�L8�d$?_�{�4�����r���)�l��%���^{*p�������F=�[�>#{l�l�  @��XQ� �����a���`�?\�����Y���z��_t� �7l@E��� l�s5����@`�i�eY���lC3����WL�.��G����n��y��\�x��=��BcC4��A�Yz�u\Ǐ����n�$�f) g'�;����:��K9'D���<�3���(G}���X�{�Y@q2��j*�8`��z�~~�AGf�g���i0{�v�f�K��h2���_4��hy���w��Qo�/����=�-�����nΝ{z"	���H+�e�D+�d��Òh����e}r�J���T4DJ �$E
"	�H3�:��7Ǔ��{޵o7XR=�s����Z��>���f��{����M={��k�4�q }�i.��L_�lcŦcԑ4�á��\�.��Zz��k����]������?����,{�D�s�KX8�L�`J�Y�e�6����F�lf���c�-�5�5� �aW�Y���#����6�Y;��j�/�d\!r&������0�#����u�:	���� �2�g<�,_���?�ݽ]�}�m-m������':>8���V[�z������^)X�:�ߨ`��s��P�{����]�VC��B�/���詺���f���ʰǑ������c��h�.����~�\��}�����_�K*6�tys�ӗ��	fΨ�<;!��W��p1��E���UI���o���h�g�y����x"<���ݲƉ��x8LøW��ˎњ�\�pw�N�C�Yo������;֙3�ᙵ]s�'�7�����Z�kO79K�䭺�%:)b"Qz���'����T�F[o���77|�9��e�@�N��h�Rأ�����q���ۥ��%忳��M]H�ߙ�0���eU�3�-�¨��������`�*2���sc�
k�8��0�P8����j�ȁ݃�k��R��?�d@Pk�7�Uhw=����9QC���/�@��hp��#�����-�H��:>|���֖�	�1���er�e�B�ͻ8=���Aԁ,@<�	
јeV�v�MQ������V7��kA�T��\r�k��Bib#��-��Ӕ�G5�Z�/GG���cĘ�`#	�IL�����{7W���I������rӎS^���Ì�1�/�q<ܑI��(�}�+Ֆ�Q$��>�}��]�*wZ.��㤉�t�~���6������$�AUZ[Y�}2Ԛ�<h����b��d��l7ژ2mI�T���Y�͹��,~ �g��9��u�+C�e3��'���D���#�w��`
T���� '�km7��X��,9#�V�t����Ҫ�z7}��ΥޕDn�Ǐq a0]��j�"��y��S��!%�yA͵--�o� ���)�in@&=�����X��
U�1&�xB�\8�"����.`�R������"BH�b{�B|�ga��G�f�_��24
����d���!s�1W`Su�������9.����i���(�,��kSXq�b�C�fp\�S�|�	���k2M�*�@����A��\����;�E�C�_������)�!��l:�m+��1�W��$�:׀f��������b���
MvɃ����.Δ��U�`�{�B���f�{��)� By7�<h�h���������M�E���Aa&ӏ�*�Yi5��<#z�dw:�d
���Zֻ�������p@N��Q�Q��2Q�R3�����LI� ϟv�{��1tօq��2�i�6����Ξ��W=�#�����#͎�U�B���MH.�ML�%���
@}��!��ǘ֕c3h�{Zٻ�F�Z��gOu��o����8�P��:�]1�IB��:���U
y����w�ş�������D5g��S�#V�}��!/qn-��9�	��{"�-h[ $!�qO�l���|}dkba��hZv�����*/���u,!�y{u@l
>��PA�⍏q�Fv�����{j.w���n�����_�n.=ɞ�Uňd��_�����0��ě�}4��?��5S��AFrU�?|���fC���������'�fa,`'p���A�R&E���Լ�܁�G�N��db�� ��|�+vN�њ&�}��&�V.y ��!�o�۳:�Enhj�'���U���v�B:��j.�Q�C�$N@#��M�M�I$�r�s�'��ȕ5��Pyv��h�q��򂥊�[6p��}ݻs_���o������`/��3@�k�Ʊc��F��f�/
zq�-�6<F�*-u�|��Ʀ����u����-}��齃�Ҽ%��=�z
H>��p��c_��匟���h<T��֓Ǐ����f���� ӑ�=N��'���	<�ù>c+��f&3�=S��uC���i0"��f��Cf�n��<t_L�o�j-���勉��+��߷�14��iQ�gYG�Rb� *��L�Cƫ��������@������J��z���8s<�S�����͖�e�M��P����-�*hl�����_�%�; [7z��S�����)���8�}���^8g�0��;s�We��RiQ��{;;z����Aq���}�7�kd�{C�s��7���4��mh��C��'c��+��S�>�����=Fd��Yc��jkGk��*ךOs�X k���'�k�E�������tqq���M����.�L~c�7�j�,�˅��{I��x��Z.1Q���A#5���?�g���%�.r�]8;J��������h152� o�S!����4,�[�g��P	��a�A�7Yl�5�C8Xi��Br����!_�{*'6;��XXC�B��A4���-�~L����a��\���M�F���]҃�͍Nw���T �[��͠����􎍍C�	�:���Z�ɔԦ;󀮙��p�������E��|�D���Fs	�C6Nn��M���[:�.�i�	0;�РD5kS�ظo.�t�ц�4J4\8U�� f�L�����GTo)�v����"S�㒚�f����M��kLN[j�5�0Ed�r/4(�3�L/��������[e����Ʀ���Y������3E㔏&��"X��4L&���A\�0�>|����] Y���'�St/��R$3	G�K#�#�6�D3���0�g�M�x&b.^�f��.���V3rQ[�P�f0_��ŕnΎ��K	��(M�r9��2a��+/;�(# ��ń�Mbڃ���SU{c[K�~>n�}]�kN,C�U.�}�<07�!BV����F
�'%�B�[;z��'����z�K�iSc�SJ,�_����+���zQ\�^�u4�#��Y�7��%M�l4�S�}ޛf`��Y̝�i�݂����3Me�T�Up�0gS�<�i�P>�F���L���-�ie����f���N��9�j�$?���A�~��U֓Q�9#���w��´�Q�%U1�Y^�g�z�<����81��6�5��45�<LCr�
,s�b���!���c�z�������vG���5Z�T��{.坝;�&3c7�)3=�_�C����Scg}_f�����T�%�S�c�z ��k9AU1d�3_^�y��1DS����1k��Uã�uUAc�S}�g����eD�1��s�AT����R��wM[�µ��[�JMշ��v��jY��c��x�|*R�D1�~�e�\j�|H�Dş=8t�|8?���9��ߡ�]��Z�i���4��gk��<�����4��)�2�9���:�'H�����-7]�=<<��Ñr<���b1�dl0cfFb�؍oaD�:�(i
�����2�����2�ۿ�뚞�����Z���E��b��Y<�<sF�)�(d܈��L (׹�pd8�o��hh{yI������Ah�g0D2"Ȧ����F������Ч�=4w�/��-�P�|ܿg7NN�X]�%��Q3�w��2�B>r1�{
v7{h�l*D�-� C�h4A:(p=�d=��F�#h2*��U\��cgWؠ�yO� #Ů�C��	C�	qs��v����R��G�z/��o��>��De�v�?��}�6�EiR�yh=��F�2�<{�%Ь�VB��A3���?����'?�~j4��HM�  �F��Fz��,���%:f$�@Vy-u�z�豛B��4
�-9��/)��Y�0�|��{``Fk�e(�6D��]/��l�U����_���.��j����{������s��߷��j)�V��Ԇ~�D �p����ɀ��Ƶ�,�￯w��E���~_g��T�UH����v�3��*���c(��2\��-�9x�L��lds�����/|]���=�z���0�8�.��@�x���%�u�4��N�$P6A�1�����G����A$놺-��Zl�5z�1c�|���ch9�0��h i�{�����U�p5�IR�Ϡny{O˛[j�;F�k:�@a�vB@������\�[���# ν��w��+0vȂ�g��	��W�
��Ģ�ɚA?�i���$�I b����`���f�3f9��������x1���:�ʅN;l0S�Z.����/
\obl�ic�FRHGS�|��v�]G1Ht5�W�<���]��f���Ta�R@���!&]����F�����'�h3#	���Ȱ�]]ӝ;{���m}�H���z?�y�n�����lt��J�x�5q���b8t��f���{��y����u
`�͟�rm?��k�	�!i	�a쟓�3�s&%H4�q�A�l7�l5��nNOt}�
�x��x�Q�j6/����gၚ�H2�5h ������-l5��6����n.u}v�	S*�ꚻa���ه�#8B��PN�z��=�&_f����0��)�C��ޞV:Kf�`fY<��F?��p7׋ϒ�0�0H�QP0��M4�6>��*;�AA;�-�籉��|�Z3��3꼠��.~�N��g$5Q���T�E	�F[��u���;�]�k�YÆn�l��<C��{}�s�|�nAa��9@����\���ƶ:kkF����N�� �g*���f~�3>+��A%�!�T�Yr�����w8w	��t8"�$��,l�p9�=$t�d����)�����5{���ֿ��27�}~fÌ9(Qa��c�g� !��l�P�����K TC�4�r4�)ohLc�i�SW~mSݝ]�:-F7�9?���Q��-x�FL�٧b"MÖ'c%5��p�Bm�NL�'<���ֲ*�uW��*ӿ���K��NUq�Bs~���M�H��D����	�dL
�DxXWփ���[Z]^�"���Y��Q ��M]�z�p���{��$����{����^L���+Q��P��$ܷрqM�2�~�6�l�`d����pձt�    IDAT*D?1/�$(�����lju}]��B��X���G�>W��>��/i��h���!�5���tA�Й����3,�U�*t�-қ�>��u��Evx��+̣�s$$���7����;�g�l�����56���M}��z��������kevNB�����Ȉ������~��q�8���9t�PY��#�4����t<ӌ�֚l�p�N�M<��lv�]�
�DJU-`v������]��O��������f'�R�B�^�X�i������H5��(1{L��(Ҍ��>��T�fpQ�j��[���\khm����ֿ����,��A��I�f0h�6m�Y� ��b�@?�ϘI2��Ύܻ��G��ln�6�� �-"���R�y��h`<:��O�0���`�e�� &�oAe��~��L�rA=��"C���I����6�5���0O�#w��1������jjgsS�BA�cD�3��C7��s�2�6�� `T��|�`c�����i��Ai�Z�&�����u��E3������l��z�)x9An�g��kT ��d�C,_�$�V[����vv-up��!��/jU������X�|���CScC�:���e�)PZ�0@������Yd&�85�M����m޽���r����ın��i~����ۭsLF��Q�Ԩ��[[W��C�}�mmo��Po���S�M�5�1�m9�A�D��D�1����g'z��`~6�M?������Uh�:>��ŧ*2Ȏi������ɾ�f �4�0]�q@e$r�J����Hu��Y���;���{�n�����9ۑ}j��A>��FQS�#��S�q.��z=q����$Ɍ���_�^W�����'�MG�����
�M��(�7+X�<��Qpe�Ӌ_׽��u��}+U�0x��$/��^�w��h�.05��7Eg��:\��ft���7��h+��6�=����4����H,n
o���)X5��1���7���(���z/k0��i�D��+Y�7�5�ݸ�s*�O���9�+��:�m�:k����Skrhv���(Wĕ�e�љ�ֿ��ר�-�N��h�8�Ly	s�~�>A����Pn���ߠ�r�y�.���O�~�f
�v�PBP����
��)��д�<����&*|A��j��86��ɉz�@6t�^{�R]�!���bl�LQ,:Mֱ�N�P�y�;c����`[|���B�'��\+7�q���28fX�Cj�s^E6�*��"��c�zt  ��!,�^���7�lm��.h��#�����"ք9&�	�v��a��`F� f3�h�sA���w����Y�ߦ��M(���)�0(����0�������쪱��s�9vg���4FӇ-��	T���9�U������Fi֗K<��(XrŚ��[j,-+�607���Z��g:���)6�9�������Ƒ��}�����z��;vEg����bB�2�rh�b��Vę"i�h�,h'������U�.��K�лY��6k2ip�����7ݝ�CSj0g��Z���5���[�TC�"8�9*���m��J�RE�i_W���_p�A�'�Ĝ�{�.��x�a;n�2��f���!+UUh���]5M��Ҹw����ຨ�*;XS��C���vLC >�����v�ы�v�wv�] �?��؞C,P���;<��0~�B�j��X�I&V�"y��&��}�fc����DM|k�FB<|r�QB��g�  �b<{�7���kt�����7�V�\]v&��䦯��?���@��͠k�;Ƥ�P�p"ť4�)��`A��&9
�o	c�����Z�w�{i�TЧ?���^��S[��Z*W�ZKï��&ruj�i����?ΔJYۻ�����X[��I���_�j�5�����=d_�䠧9-�&׷(H�?�d=����zxa�̄��q���3c�pϢ!�ge1�����:������Ҋk���S7��k�WY�G���K�T��x�	b�7�A�����f���4ߙ�պ�XU��|�D�{�Xm��{��7�󄅼m��5���Pj�yz�A�^žkƛ#k���nք-u;m=z�@�<��Y�����횢)�L��v�=�ila��}���Bo<����k"y�Q�.�"b��V��VI��>�i��{��,4
�R�Es� �feK�ͻjl�Z�E\�f:�?��?�S�����0��$"I r�6K�`�2���3��ad�F<5�S����V��of����v�~[O��Z?�6Q[c��|uÉ��7g%O��p!��YN̘�U��������3����Q�]��g���1�3����6�;y
�//�p�����"
�?�k_PP	��A���;���䉪ݮJՆ��/���ժ7uwgO�/��O�RN�3�913�l'C�i�bG՝]�~�V����^�:Vy4���ڎ�s=P��$Ҍ,>�����yf_�<8;;��Ϟ�X�)�6������Bs�.�'����ce�}�����DE�yj�s��|�a�`�\v�}"B�S/[�R�TT#������4�Y����`�G0@�&:�� YG&����D������������l4���i�ryiU4�0�<�L)�Yc��&���e@a0�P������ݻj���8�̑��`��TO��fOT	�����[
h�m�KA���C�K-�@�P�z��?�_�9�<��n�a�F�5��<�7˭s�cj)~��h?p'�&��G�s(A�*�x#h8х��b2���3�AS�B��D�T`��k*��,�&c�l��d�&��c��0�l.h����޴�3�nx��x
��"�[�Y��5��55;�qd�`��b�C4ϓ��YlI\D#��p�ɰv�����iVL�#H��S���I�),$�AW���*�V�*N�Ƛ��/�@/�.[*����� e�+{\�I+�B� ǟ�
��B��]m��XR�����s]izu�����-^Z�d4������Y�1L��m��}S�2�$��X4�fp���&���b��[���	ai�263�]=�ץ��N6�0��;: �:h1�褢,s0d3">���T=v��q8��:FSh���5i�yLv���<f4��
��r�"��rx}v�I��.�4����6���
���#t������S`�a�U3E��K*�ַUi�UlRIG/>S��FEP�\�!(jYj�	�:)�g®�h5)0�b�a�����{n���2(I�������k`_�������?����~@�|h�o0+��İ�/���S���U4�1L��UЖ��$';&�P�f��Aߢ�T��	�~ź�+��6�*�r_������	�A�*���-������T�^y�2y:oS(HA+�b��ZQ�����7�!b�����.p�cz��aU�l9ĝ
Cߠ����`��MHc4�w��@� �鲿�\ߨY�"��9��wS��%�&>ۣ2�_6\�w�!�����'��1X�E L�
�i'<�t��'탩���:�ť�P��r�����L7D��qMs������_{\޸`���|���E
�}�Zߩ)�B�a((GM��=m<xh#�F)��~�#]쇼 qX��6枂�n���)�m!��#l�����&[*Y����U�ah\h�AU6e�Èj�q�Ce��)#�5�0���б?�,�u~viT�)7��v����>�'�`�#����ɸ��4�K�а4�C�����M5�+���.������L�^_���	�p1"��Z��nc��?����h�0� �ոP�M� k��u�������2��½�k�g������&�P٠\;	�	�&f%�3��f���B�?~�啥�(��(��1\O�b2�3�
j&�*)m���`�b�@3��p%W^룭�����#S�g�f$(��'� )\AT�v>e}�b
ÞR{E�w��}O�ZW�jC�������g���<S�U�l��J�3b �x��H1�P���5{$�VԙPD�T�i^�K��Vފfdpgg���'?�^T��Bi_p�kg�@��`Gc���'�>Ǟ�Gf2S5���h�[]Z����^_n�f#{�"Sc)�^4FGCk�p=�H%�NAC��f�n��7h��� &-YX��ZZ���/|A��er�-p�����HKͶk��/tr|�B�`} Zw�)PYj�a�yfؒ:{�U�X������)����M}����)T��S�M1܅���t�`˃0C��9=~�����E[Lh�&��%}��_V���˫K�<Sq1z�r�Y' �� �~H���X,(�����ֽ��'5���Wg*ڠ��O}̅�)����n��2~f9#�̌�f��*���@�v�����Ғ�;k:�M��k7n�;��	��C��F��g�����`2�����w�]�A����d�>��G<?��a�QW�ͣ_,�E�Z�� 1��4xFFH��7ʚA�k�����Dk�i��bH2$�&0i�LC��*�`lf!Wz���B��|�u�VP0���b�(��0:�X�� �

2�]��g���'�ql"� FAkh9Y�e@{a�+��يɺ#OJ�7�v��.u�}�ۏ��8�<T�̘>��m��[���
#��!_9�S�2�@�H0hL�~�>*E聨���l��3�xq�3�IbP��%ϱI-uUk6��nn�?<���T�$�G!h�u�Dá2��R�^zQ�-t��s�O�V��\_R���f:���QW��z�P�ۦ\�wŔ-���#.G��������4O��CK����<�\�j��I�f����=����3��Ę�O)L��5EZ�52Mz�F���h-����F3Д�.�S�˔� �)�Lb��'.���UjPJ������%b:]]^Q��p�W�PЈ���H���F����z�f2g�.EGY��,���xM
�l���bTP��T�f��r3����O	.S�������̇&Z��O��v��j�f;����B�X���:tuow/ewƁ�I���B��'�aCK��LSG��Kk�ޡa�y#Tq7nx�V�Ze�ǘ��kk��ex���` -cP�nP�U�W�0-�b��rQRht�Z�Q��5��~t��F�s��Q�+��Թ ���Ix��r�o��ӭHb�#!`^c��Ʋ��e��@��B'��5�8
�J�=.��p	͆E
Qe��R0�pS6͗f�\U����c�/�$�ܹc����SƟ�"��5�����f��<���{�!�h.2� ��m�SsK��^���G�}P��� �}8C�M��Z-4����X0��!��u��huL�$3�|��u\Ch]�0�����s�`B���v�B�9���~J5�w�i��#�B���C�>����ڱ�?�@�y��s�s ����=�3MZ �X��#��-�$��mnn���+��yEy-�4��7��b E	̊�e�;z�Y�m0�����9���!{� �1���� g���V��Y�.�'�+��3��w�}�צb�Ǉ:���&��)4��P�5�9-�(` ��E�KnN��B�ȳ�uڵ��X�vm<|��Ʈ*��6����oK=�א�`��D��µj���Q��q5=�)U"����Jj�A�����q�!KY]]�af�lM��n���w�uƨ���!)���c��}�v�3ƑHx����5��T0$`�d�D��Y�vʘOfn�na����K��eh�{O��;���լ��6���':��c�{d�r�U����PL3�F�g��I�PS�}���!��JS�4���-����b ����t#���D
95g��TTtF����bA�u)�B��8��Y���ժQC ����@���Pgu��%�l����c��W��es�iZb��T!"��e�P+�mt�v��{�����{:��������08�<<1�Q�8�v��H�~"#�0?�T�nhu��6<V�
��][LozZ�b�FsД��s��w��|���#J��N�ڼMy������L\�a����_�K:���������z���`?�0��S)!�&�p�E��c���.�ʫ���� �hh1�9�!
�
�&j�`�qO��줙���H��0
�m���j���]���������"4���u��֑n�ƒ�>����Ͷk�����so}YB��žƳZ)��@��T3��L��-����U�9&�kd�d��b�ϐA�'?���2�Ó�4�"�����۔ZA���Q���1��iw,�@	z��[��������W�����Ab^�H�d�i���3B�C���#�j��p����:�F� ��d�W��������l�ĝf�~^��)s�˚~7����$��O�����5�YCh�po~�9�/�z�C�y�ez��s�O�����6-�2��RS�r�ך	L���p���A҄0s3��s;���˪r��+v{:����	>��P�0��.��h�h7��t$�����M	���B����R4��f3 x����&�6�Ŵء��|�9�g؍4�1Gp�1*I�k��I;H����.�N��8,A��)Ӽqh���I��bŪf�>/+W���h����I�����NS 7�4A������2E�0%��<�k$r��XX�������������
����^>S��F%"[�g��i�����S�1ϛ$$,%H�w[X(�C��yB
�F2 ?�{����6���A�t����3�� ��6"��_��Ί�8؃�:�b�"���	8���S눀(�j�cbtw��i��騴���ږՎQ��鵆W�:=yft�ht�%d��Ԕڐ�Wj6��4�\�F�3�R-����;�o�h�RV��L���١�.
gf��7qٳ�!�3dñiZ�����|-i�@�����ۏߺEu�՚�0<Lō�V�L1��pKq��Κ��9���A�{3��u�E]�]����:�Sn>���VC�I�U�k�<�7{�;�i��ll��{Wͥ��L(��^���3OAVg���cs��H3�v~��-�6N3��3fd��2+��.n��ߪZki{���J�����Ot}�ʴ���,��9d	���A6N�>�������l��o�q�&飛�Zk�Z[]��14sAwg�Y�^��P�fQ�K0K���Ǡp[�;��8Wg�k��4̂����A3
��%��eN�4_<ۜ�k:�R�q��E3/�l����uB�aF�F�a�:<�+"�!�vY����ֈ�"h�V�ٚ>�D8H�<�`�` Gp+�����\�Q����ʒ5���#�t�$m{]�_�F��U��T��'�� �3���̢���$���|8r#��F��?��"'��N�z�^_�Z%j,P�S�h�)�h9��]�$U�a�����Ȓ�D��T-�Ş����Iu�*�7�^��yՖW�r��KZ^[���J�O?����^^���AZ_�V��#������y��A�J�D=.�ըO���%Q3��}�]Ֆ�t���������o�ُ��2�P�"(�PWj�:(��%G��������U R��W����gΗ�{�¨
Wn�Z���ૡ���6��#9'h�9�}��D����D���Y�>�qHM� 7��j?�����	|ow|K�O��<
��a�E#��!YbP\�h��#�����֮�B�'��\��˫]�[1�T(q�C3x}u����N���p�����g ȞF�{܁n�.t~t�=b�ݟ��?�5ͪ-���}�<b�{��+�6�Q������{."'�e��4��faF1`��)���*��i)d�16�*���-��}Ӯ�췕���)���:qA��g � }s�`Hn&�[D�d�c
[��$v ��?Ћ^_�[���÷޳�Z��ə./���`���8�^�|���kc#�9u���v�vϓ\D]o�h���io�h-��0�{4��    IDATf�M͠i��>4Ѡa2�dR�1Y3�A�8~m��rtϛ�M�F0���N44F���3�b���f��2�s����A/T��⛆uY����f0N�l�����F�榣!�^Z�A3zKA�t+q�d���/��y��hCÉf�n?�nl4�h3�e�8ݓ�7�o4���������4�>1�Jv��z���ȁ>����7=-0b���8����Un9��E2����^��qO��[{��*�5U*u��%��t-
��)_O�i'|��dpa��UX11�h(q?��N��IovSٰg�A�lכ!��D�1&�Yf"��3?�	�e�a�c'��ï#'˔��2È��p�����{S!����rn�2���T��Y�b�b��z{Y�FU�&��C�����X�#i��~����$���f��7����FjA�ü���� y�v�������f0W�i4�0�����F3�!���#RћEh,���!��tL�D3�i�L!���2"����d��I���=S:�5� .��m��'���!͠�3"���A�#&��Y{#&�(+
(��G���- $@ۿ_Qڹ0������*�,����F�c����J��S��4�G�fRvkLS}�/�)�q�}�"c��TM�Z�`h�V��4?��*���ع�fpu�W�?�����k$M������E:��&4g�e��R��P����3B�ͩ�AT�j�ӽ�0�w{#�@�L�:��#[����5��i�BQ�&�����4���˳P�9�èI�'���%����R9��=��4�u�F8�3�+Ŗ:�n悔�e'�24��3�<{���pS��ѯ%�A� l?�+/^��x��kݹQ� z�1U�>v84�q�^s3�~�� ��19���G���e<F��:�閞�����ٴ&�R�F!P���e��΄M1uΪ�M�Q�,��H��u��`�=�P��s���Y��\!��b#���3���]�Zӈ!���BjvT۾���;E��zq�J�^htz�4�b�\8�5X<� 9�%&�o1��!���Y*�Q��g燢wwa����僧��:QSݎ~�[ߴ��]0��q��ͣ*M����f�Έ ��*�d�[b\�T����d#��g C�8y�#/�W��CImh�WQ1[)��r>��x.�n��b�5E15�����N�h"{C����3�E7��_
��f}�r�vֵ�}�hS������X��=��g��Y-��舸���݆)�sH�?��Y������g�Cv 9�u���a����~_ե�ypO��o�ۿ������D��羊���=!2F���R�&-f��3r9wt��V�}��K �A[��1G��K��x^@�t�4�yr.ϿϹ��rÞbYh^+m����O���,�F�q�eĘA�g���^8+��v��h6�#�d`�^'�{��y���V�=u4��z�pvXF4�������`�Z����]�jkgW�FU��h��h̀ä d�����s���j������>��/>�9��!��&����dt����;e�&$�5�a�\���H��ʹ��9�����cogqdV��è0�S�U�\*��@��]����g��p�w�U��0y�|�"�C��r�������fb	���������>y۞�ӟ�^��f X'�\�g��a�v0�k�*��f�_F5S!�'JM�-M4e�޺�JS3�|��Z-VU)���������4Q�[3m�m�\E��X���%l�&+.�S�b�p�Maj혅	Jvȅ ��^���__jvCN ��vF���6��_�~cb~�$���a4��p+�/���yh�_l~�;�x/��1��cí�3�wkv�}�aI�d4&t��T�K�R�#�6�Q����+!�oPjKekH�>hp}���q��A����N qS&�źm���9�!!���[�$�_Д��Z]�P�#S�����r�lr��1�12�}�`�:k.X8���<2�x	��Yh6/�Q,N�L��i��ij)����;5'�n�3'3��r��u�Q���.P�-|��I��'#��o��4����:w��\IS��T�u}��]�k-�4��p�������l�<wv��V,v�]o2L#���T)��qFT��yю��F.�u5ַT_]Q�^�p1�ŋ��مJ�����d\�g��,�.���Z���S�DE&E��GڼLOs�vzv�I�?�R�x� >!�8��)�t42uѓm2�| �TH�Z]o��,_�R�#e��<���л�c��,�=D
�uM�iƸ��{[*/wU]Y���]���P��ǚNn���T�b��9�������" �D��b;4���)��pT�6xCqS�������{n��NώL�)%d0���훮�ik���*Ek�p��7+M��
}�f��\ĸ�AUd%�1�L���X����L&�Ȩ$h�Ӹ?.J�{���)��:*hj�s�x�S���La���t4��-��i��D��U@#�����J��w�˃W�:���@�����4�}������m�M"�M_�1�o��ʄ�·�z4�4=x���=��ZYO�':}�B�f��]yg��f0Fco�zC'�F2��[:pj�1`@�ǡ1�l��4ձ��]HLOM���S�V����8�L���/�d��u�L*�F�.�_~�	O���@�*�G��g�liigO��ju��������ts|�ܸ�*���n�p$�,�}�}a%����T�����w�hSޅC��@��}�}�kn�ZM��o}K��#Û֖�=�&n��H*;���*"J�i��g/�#�x�0�&�s �^�L1ʍ���rHp$���q�fe�\^���H��"3�w��^'-8_�"���R�=���U���s��	��9���������GZٺ�Vg�{��ɩ^��Lg�>����u�)w63�lf�fb�ُs�xO d�#���B/{bŔ��5���A�b��X��{_����ޮ����;���u�я������<�5q�Ŝ�b�=1����"���o�����@O�6��D0��kl��b4A����J��a�n�3\y�dNQ�uV��p��O`F�k�ua^�����Ξڍ�N^�����֫�Wz���Jn�����M+Ŧzd{.f�.w�����ή�6��ju5��.�^�U�5���м �ɐb`d�٨���H�G�o������+���^N���0o��M��b�������T߾���忪��.�.t��c�Q���ȧ)���$(��+�D�N:�292�v�=�&�(���U+�tsE�d���4��C\cӄ��2�h�Om��Z�nV���O�������}2�2X�3��� �uFӟ%�9�2j����'�����t��C�޻�����ѩNN�\�ӑ-�p]�h���|6&͟�����V1mw~��{�߃)(�c�켋f��Z�f���}������&@�ύ�(�#Z�4H���H�E�kQ�[� )��
Ngk!�X��O��
��L�F��D�h)�#�"6��Dz|��	���TE��]�'fj��:r�<�cA��=h��O�e"c�|��rԍ�����G�����7�GGq���S��Os`t��]�P2�)�Tm6l|�d���W���\IÑ)����c	��Y4`sE"��5<�02��f*���āh>u���ҺE��Rс������r=�%l\����Fý���"4Q�b1d� ��Zr��Zs�B��&���F���Pe�1�c\�d���T`eS�d�����Yi-,�s�`fdń�7?��YmyF��V]�JC�j[�抪�nX�Ά��O5�>�{��4߄��~�s�C\�Ъ��a�D$
����<#�4�|�{J6�RS��M5VW�k�ns�g*��3�Ω��S�1ft�(�4=���L'��lZ���7�����Y�LAo1s
&��yGco�6N�^FF�M�⯇
�����DO~�!��@	I5��A�{:j*�*tU�I�� VZY��[����n�u}p������=�rc��m�͐"5��O��?���Ầ�pZ��tB�"�3s��5ַ���g����J��>���X�����Yy8�Z�d���C�����&�l�*���(+��k4�<��?eMU{=��DaQ�\�Bu���9|�}�H��$,�!�pɴ₵�Lk��-Q��J=�2F	����e4��� �Ri�����Ɔ�k�ʷ��o��.��'?�����T��G�h��{ -7��}�� \�37Q����pc��9;�B+�4�p�,7Ը�P���\)�[.��|Og�/MgM�ȴ����$IJ��3D�v�M����HJ�)�+�y�C�p��x��M{c��|�ܞ3��S��K7�-(b(~y�ȿrc��2�{2&Q�psv\����[Z�����b��-���66��}G͵'S����n|������q:t>Y����Ɔ&s�'I8G�J�e�U�%7P��S�R�u��>���uVU�t�T����9t~�%��@�B��u�Q)�`��ZٯT�����GH���i8��㣎
��rX�ۣ�*!�9��t�~���~�z���4٩�D�Gf{y���M�څ%��'�\#�������Ќ���$���T��5���Ww�:�UK5����?�P7g���#�.j<։�)/��yD��ن�H��k/D8���D�W�g�5�J<g��B�z[k���oh�ζ67��������#�*�ab��J32Ǡ�?��@.���+��z\q /�� @��A�l��=��U�҄��|��r�g��4ꔩ�H&�4���iT*�B�����h4��z���5=y�D�ZC�����z�����|��~�f�=�Z��+k>-���b����w�~���++�Ԛ��~�RWGǎ�Zj�����F�Z2����ñڭ����ut|�8���u�<8pN7
�J�E��S����X�����>R������M��=���4[�2��R>j\/�f(�����ء?4�F�#T�tZj���JG��5�_���^b�`@5���p��55+U��j��.�#�U(T�ηB�[���T��gj����������Ϻ��tuu�F����NkI##�A��jL�]g�fk5�:<<���w���'O�(tyy���+��_���]�2ˁ�l��(1\��b�Mh�s��ႝ��T� �u��F63�y���I�x��{(���)k���_��(��-2HqoW��w'�j���L3�>s�
T�79��[-!ӗ�>L2�XT,8c�;�<�A7���e}�g�h�F��-��F���]s���	b�`GD i܆��c1耡L�g�0�����T��Td��7N�[ʣ�PS5v �gK���73��.Ɣ���T���m����l���ks���;���)'v[*"���J!S�8�����N�&h}�"��¤հ�*_Tsi-��bA��KkՇ&j�Xd�����Əu7�8�#u��9��C��$zVБO���"�w}mM���Ix�6R)��ZU*���49��"�3��eYf�<�ܾ���E����$���'щ�8�p��έ%U�]UK*�k�x��/4>��lp�C��XX�7j�_l����4��j�R-�!�@� ��b:�Ä
� ��*4�,�:{�L���qB}#���q2�d)˩Iӱ0�M���S��=4�>�>ǭ1�p�Ĥ���ш��F21^���,(\v�
ҧ������j1��M�gLuc2F�;U4�[1!�ƙ>�!S)��6��Y��:ۛ�ln:Ts���#�_J�7�On�0E��AϠ<��؇[dU�8��:#�	t�#��P˂r�e5�w����5>��S�Ύl6SYp3��@O^��]���_7�o����e��G��'��һЄ�~3�V�yS���펛s�cS+��pg��2]����8Q=��|55�u�ݱ&�O����`ওc�T:�.q.�KFx㐺�q?�%'5V7������Ma�r|t�����%���B	C�EtL�;����9�#�\b��ρ��bd��1<�5�������Z��F/�BNOS3}���f3h�>g)�`:�}��a\j�А���j��z����`���y���N�RĜ+-�b�l�	f���@�5k�);zQ�m���d6҃��\
{�uNMf
��&-1״��jukK[;j��F���t��n_i~}��"L��(!}C�gl�4��,ܯ^[on>���<[�k�X���Tԃ/~Q�5�f�j���w�����'*A�uv�	�~��H�4��`̀#�A�k�ĮH�`�##�l�E>FCK̚*�`F�p�c����׿�l�^0���F�q�M9��7�9���k���3���&U�n�J�!҅�JS3�ą��\��7+�g��N�x���Goim�J�n�"C��T'O?�K�3YM/�a���p��`1c`��럚A�*b��s�L�9���Ɨ�.ȯn�ʕ�Z~���vwu��VW���o}C�~��@o-�!R��u�[�U�����Hn�Y�I6��, 4�T(�됳.�x �5�H�=�C/����2�3@z�^ĉ�*�כ�<?w#���1f����ZM谹?��H�7=����u=z��)�G�ZY[��ɑ��xFk�; �����]�U�e߼�@�[;�S�hpu���/t=~�S��v��I���V�m�fhMk��F��e0�Z��N^�e���g�������J��q�L?"����/����՝;:9=��'?�OE����ʘjo�`�%�I�?L��Qk{o�iL���ӓC]_k����щ=���)��@����Ɩ���N_����
ͪ&��z��ڝ���lDdUL���NNO�b?��Z�eT�%�j�m�[���6l�Z�		�\ƨJU�Ƴ�OOS�s��=yWUh��Wn�O�4 ����lg~L�xz��,�->5����kd"Iu�������eb���C}8ƺ���&
��uP�4T+�UŐg�o����87��M�� S-��X4�F3h��2�t�f0Q$���q�L��h�h�N�v��I7Ns�k�����-����LH�]��jC��������hP��BIG�Y���M�݆�9���_��D��� eMcx��2���m���[|�J�jjT��V��t�B&��ř��|�c�k��b���I�
�`�
��.Pq�`�-��f(Aw��uC�4k-����U��p]�����1����#��-��j���������� C�䘉!A�V���y8�Q����f?��l^���7�8,&���B_�Z��L��������0�J�v�r�n��b�^Y^Q���r��|���"���k��^�A񭁎�:pNTL�*Up.t��+�2���ş�
�M��q)K�U�jm�:s�f��ًϥ��M�yM}���M6�Yl�Ӈ?�4d$t�~HS��eoz�SAcM�g�Y��O�FH���C��*�%�����5����ə�����3vK�������.��s8����ZSueMK;;jo�k2_���BW�^�\B�f���Z����E�/:�C��(>o����0,�#Tz1%�WA�撪k��ؾ�&hpy��ϟj�
x�]'ʕj�MT3�y�C�Q𩽰3�F�������V}OL?N�i�P~.����4h�F@o�����_��E�s=���z�b4���oĦZӔ��i4m��Zf�߿�2U,C]�<L�W�*v�j�mji}S�Zˮ��g���r��zP7��6�Q(N�kr��5�x��aD�����dc��o�(�km5w�j��k?����߳�(�q����߳K������"�a������P�lsbH��g���o�x���^�wt��T(i�����/���6T.�xH9v���0'g������,�[)XpћG�Nd�%��y�b0�� NG����m���]v�svx�ӃC��<���C�����@t(��&r�|�R�Ǟ���#��E!����d� �U3�����ٓ���4��몶������������vѬ�O2�5�k���\�`F�����    IDAT`�2��r6 O��F="���#z!_��ɓwT��u|x���@y�K�Z-�+�,������ԟ��w�&k�V8�[���9�v}k�n͠T�ǧ�Ǝy�y��V�㨐��={�L'�G��L�U�:9:U��R1�qMh��y1ʫ�������;�U�.��:>x��g�L����"o��.fudmBō=��b�ctt�AAk���H:���,5p�O���c����ԱHˏ�������R�Yҿ��o蓏g�'��IclG������#�����]D!Źm#��jM}2zx��{����5����$R�rj3<h������F]�������{�w�fz���ͦ^��F��l�g�+��/}�����e���f3D#րح��P?���h�T]WW:>:��'jck �|��0������Z�G<=�#���Om�aIs}U�&����װ�`��y�k*n~��0 d�@c?�H]��3(��BQ����Ւ#�~����Y�_��]��u�|��g��͜��eMs5��4�����#�#GMؕ:t�n�Z�	�h�]��������_~��VM���7t��@ե��zH�����������ً}��7K���P�Ӟ����km��m�4*i2��s���__������������_{��2�iusC���7����׍��?��_���Z�����<{k����5�g/_*W,��'z��/�X����J����������C�Og���o��hF->��"��`Cx���Y;�����L��@%WE�Ӽ�)s.0�1�5���D3ب6�.�<����ͣ�7e��:�f��/&���L͠Ք�F3�d���B����ڙ(����c�հ^�!3�U?$�Y���D����:(5a?��/��cp@s0&�s�+S��#q�=Â��P�P�`X\��A!�,[�tfc3d�zY�6���&c	(rp��d��F��y�H�G��~Z4jZ�vX�ք����F�����(eQP0;{��<��R
uO9I.��ȘW�KG?$�ќ{o�2�a�m4��ڶ�՚�}�_����"�S�8č<&jM��F�c�x*�^Sy���)���hy��b��09ӱCl��)U³�i1E���_	Y��K��Yl�s�9�YLg��Ҁ"hFJ�mS4�����UkiY�v7(׎�����\��c��tKP�ҚsG�d�l�a��m;�Ur��I�A�[8�"H��P��u�7w�X�i�����'��|��x���`6�p-��Jo y����Ḁ́҇mP���]5��[
Q#�q��<qLE��ϒ"�x�q}���3M�Aaʟ�1,��4Q��(2Ť��/�v��*�_r(�l�����ֶ��0��6�;9Qo��t}��и��ANSq��o��4�ЍE�V󙲃'eO䈢a�܇�ɵ�ۚ����-���h_}�T�����`�B�Mz���u�{E��fM�)dFi�9��+^R���a��4���]�~&Þ�Tw���G~h�O
�ȴ�Z� �{"����v�x�����퉇gf�S�����~����v�U�7��Q,�6�ܡ�n�{����J����.�.ust���vw�O�zI�FUs;"�RL��61�C�s8�@_�]lJ�H���_x���N5>�w�2���6v�j����U�f}�������8�B'��@�=[.���wif��a���~��~�أ��ެ��?�٫}Qq[^YY��H(y���!Й�$M��&&������������g����KS�*��ڝ�V76�76�=����~[�yY���X@��ވY!� ��T�Z�����j��ƫ�K���C�NO5��Y��h-��\R��� �{���4��z��yN��$w$�$��:6���&r�Š�O�jL��d�������*��*�����|��K4�u����i�V���Z��)4�����7�r[��O����������ޯ�����>�����~���������vFk�V�����������7��~���R�T�����_�������?�G=���5}��_�����\�.-u�O������ѿW��PгY�%�<��g̓G-��[ư�s_K��,�`���\/>�H7�?�#�Uu������;����T�?��Lk�9�Z�7������ym�6�Ұ�����v&(�{P����de��zy����o�`��5��f3r�S�ř��jb�mf̓�/���E���.� h�������������?��?�O>���-e�kk��_���y�]m��T��5�?����~��Z�|�]���/�����`p���K�l_��z��wt�������S��ί�M�������z��������_�����_�O>�T~���Ѐ{}���nh<��ٹ�m;_��,��:�,+*���Ʌ�>�T��?���s5�V���V�����w��\3�J�j�(�%�U��b��އJ2�ى��X~�aә>�\�ts�\�>y��掾���R����}�=S��\ȑ��X�z|����[Q���1��ɲ��b*�
6:98��O?��/�8�_��n��R���]^��_������u���z��s�,�~�LE���aش����O���\}���ܺ�JY_�ů�W�W�_�7����@��?�����}�m?�e�o�T�g6T�G��������ɻڽ�P%���Hǧ�μ:z�MmiiU�;w������qm�����U�z����_�w[�q��10��1��f�C3�\SE�Q�Ej���rE�Z4���3�v��-zv��fB�08�#��|�r|R({��S�ݙ���5�ڡ�i�A���U���X���j���Dl���s�o��"S-�%�7)�!2�r2s���˜�<�{#�&&Xv�b����=Rzu&ċ�!�Ɉ̭�5L=Ё|N�zE�ɵ�d7�:s�c Q���������p�����ê�L��x�2:I��BL<q�p�B21��Ҩ�Yk��G0�����4`�@YȦ�� e
����L�S�Op��`�Ɋ�P2���T',u����,��ꖚ��K�'�Ϥ��x��\�%sd�ef�����:���#5������7i����+S�L��W�6���|������#���N��;0�T���]Y�����ՠ� �K]L^J�./-�1�Wn;��TUhO���\Mx/\(���sh0m� ǡ�������Z:P&Њp���b e�mb�R�ؙ��x�zʜA�ƋÏ�s2��Ņ����C�Y�޵ȼH~P~���?���r��h\�ۇ��	N��������'����∛�_֌xR�t��=�Zm8f�١+s�ޡ������=�B}��72T.�y+&w܇��]mmn�����+��pB��8��������"���}�3�iq��%g[�7%�q�W����&6�s�?���L��3-�/��)<�Ͷ�<��
k�D7!�����k��I��1(��H�ɍn��tv�ʔ6�@Ͷj�[ڽ{?��+�|��� ���2|�%1�n�2�?����?;���Hh'a���KYۻ�z��yd�������qc�,/�g~���/������t��}u���F���D��?>����h&�?���V�W��;����T��������3��O��J��B�,^�&@)��0
xBޛM��t��p_���������w��u���ٽ���{/��I�H�@(	U�tD@Eԣ�P)"�{�����{2)�I2�����}?{��z�y�u�,=���~���.�����t�WV���@�"ۑ&�.��l���xdW�"&�nä���[��,��9EǩfN�Ob���H��*ժ҂ݜ��th?�6i�{	����\C��Jc�ҍŷr�o7��o?����:�N���-֯[ǡ=����PQR�W l�#�~�0C}�/η���;��O�&4�E�x�	������zT�6q�$&L���3krÕ���.'!�6�piQ�Tՠf��LZ�\왙T�E���%k7����#���}����K(-��Le�I���PȈద0��������OR���&W�$�����ۻ�s,L����;�jm5s���	�ȭ���ucM$���&�&u�"�#�a��==}Oc۵1L�u��I�� ָ܌��Ӂ)�~�DV\p]�=|�ч:L$B���3�|JK���&a��=����ꁛ�`�n�� y����~vlݦ~��S��d���)��:t�Q\R�ҳ�dե�h_����W��έ_S6v4�-'����80�3%�4����&��oN	W.O�a����n'�C<�-�KIe�
pf�\_|֢�ٸ
n�uȒ�����1��I�!�դR"3��81���#zp&�o6EU������Ⲧ8yx/�� �D���l��*َ���2��*�%z��j32��a�F`i�gH��� 2l�1s����7sd�^�옑��ɓ���+�0a<���}[�������fϡz��u�-����S�t��;h?y���6�\+�,Y�m��BiY�6�k?��}?�%��\Ɓc�hik'��@!IA���.fI�oE]�</��,�q+�]�t4�bH�Z�0N���1����Ǟ�K�,dg֔4�B̔3^��Ն#h)}W$]����L�H�� �����C�-�u��4���r��n�����D�����n5��n���3muj&ʚ7�r����e�W��	N=���d;�|����ʰ(+�CQQ�'���j#[ΈX�1".��8�P{Ү�Y��d�!ϱ�e�-ϧ٢��sW^ȥ��f��9��{9��Mi�X����
�t�t�8}�}�~�b&M����boc+�510,�`��%������:2�r���X
C�nx�����4��Jǐ��B$m��w8r_�*�P%}�H�5F3��-C��R^�5D�l36��8��`٥?O�â�	��Ћ\�Iii�!�J7B�3�Պk&cBQ�JP��@��'=e\%����ɡ�9IR\J�����Vq��~|�=Z��E	?B�9����C���$c;��Z�q�ӆ!��DLo4�fHQZR������e����|8�n�r��MVf�N������_�ѻ����l�b����NP<%��5L�6M�-[�jP�|�u5�������t��=����+�hH<�L���S�N�BT���c��Zo&��b�c��C��a��S��-3��Io@��f S���J�$�4�͐r��a�e���{e:5L��#*ձ;���ě[L�L�������1R�a�/��tc3$&d���GӪ�����@H��Q��+Fp����K4���x����8|�(��Wɥ�T��EVvY�����RZ�ZصgA�~Yͪ��\��>�:�*.a�L�]�nݪ+���rz�{������Z�I'�c��ڴI7!⏔�/[�� �X�����iπ�Bl����*�(�f�?��@W7�P��?��a�L��F.��3�nh�r ɑ	P��S7�F������7V�]����NٖE�9���Р�q��)/Ǚ����(D��h#���!�;T���ᇑ�Y�t��Ѭ����Uɨ!�U	�ȐG'Q�gw�t�2&4L�ȱf�ش�p0�~;��g�x=i��*��ٱk}�15�uL�:�.�E����ʢ��$ǎe��I���1���|���N=<�K�U����ìY3���剿<AwG��DE� (�i(uQ�m��xg�^��^�*�WU�pi�����0���)?O����'+H���N�b��Cc�^7��6�&4�e(��TR�N,&9�B8�"�����=2Q�4p)\ET����!���{�� ��{��ʫm�~��\Y�U�Nگ*g�<G�AA6��t�6���D<�˝�ͷ}���:^|��<Z<#�M]}-�'6�r��V�Z��~�3������))/��i���j��{�]�N��Ð?��#��W*!�.�G������7[�bǿ�;w�~'W]~]���7�7+lC&�)��"�U����2��<N7�a?���%6$q1�S\NAy5)�eJ{�F<�⟒�2iq��&�O�VO�x���)�8R�����6�a
3������������cqfPXY�[&9�z�;��|t6����-,���k��#W��ʦt$���~�t3!�&�lU+|D�Q߽�v�/_y�E��:����8�K��_[��%�J���P8Ơ��&L�^��|D���qƷꅘH��.����kj3n,�\-�G��Ŗ�\|�Ex��H&��mx<N��W��-��^�����M^u9݃�444p`�^�RFB��BZ�Χ�j9�U�m^L�Ի	 ,�AMY�e� 2i-�E�d#��7��_��@�,�R�yn��.�}�J#?��\FM��I��]�45qr�����K�O�,E�����C��&�q��(�A�!�o��J%�?yg�kGq�+9~�$_n����O����Y�7���6|��$aL�(�k�9���&ߪwD$#4lĈ�E�Q3A��sSZYAYu%���C�\4���!N[���S'ȭ�&�p��(.)ק���lX��y����0<����Y��340���axp���]d���$37���1DR6�f[��(�<G�0<�J`):�����Ye�C�&֖ʂJ�n6����MJ�.�ȖR�{
T�$7��֓457�?8Da}-Y�Lv�}AU
��U�O撆��)�Z���A���F@}"�aNĨ���3X��O���&2=�]���:\}��q��>m��

�9����;;���N�`�nW���-���ԏ�Ah���z3�w.�'�����w��;�����+V0i�(:Z��g!���u8o�jN;c!���6
KJ���lX����!B}��M�;oa!�|�vAl�Jݸ'�N�S��l�顩�Bp�;�3/><�֊FqK>�ɬꋞcM�}�w���pRZQΩ�v��e;��%�����"=o��"��< ��LGH���+'�X��PTL��,٩&����z�9��3��8y㥗����(����E��紳w�g�R�'�X�as�H�U�ݎ��/��#֙}>gr����_V���.�+=��@,�C�3�چ+���+/d��y���N>��O�����;n�Y����P��;�g_c3����Xw��b���j&�Ji_�\���0�u�4�OD~�����F�T���ƿ�v��߰�?N۱\(rQ]�p;��DU�b*��T ��|���?21P��R!��L���\6#�]�0R��M^4!W�fP�>i��NNb������Rь|����,�A�>q��x�W���J�T�aeo�҆V����5b�/�|=�ʪ�1�Yz�T��������~�;o��\i���7n��!�Ρ���֮���QWWEmE���e�&&�ށA� �ǎe����^�n=C�CZPdy�4��Hqq	ee8�īo���*A;��> ^���`�BE��"�r����S��7a_g�PĠ��t+ã�l1�&M�s��H��b	y.��L¨��r6����`�Q]�9�C}ݴ=hh�u[dƛ]H�Ы���p��!�� Iͼ2`ҴHQ!2@���$[!R�9�;#;�8��Fޏ��L�PU[��?��������|�2w�99���P^^J0�'$y�Be�DcsQ)~�cdx�4#F���<���t5~��1<�L�L�FGG�6X���W"YuU5{���Ï>ԟI$�Ó�����e����c8�������
�ڈLS䤁�N�fE��Q��%Ӊ�)�� �
gK'�i���M���tM�7�ZI��G��(v�݉���h�#���fP�RIl�9��h3ND��t:լ���4	*[G#�T;��1�k>�4���� 5��D�c�Gh���u��K��m�N>����US�[@ow����ݼ�!Z;;���#���`Ddx2���Ҫ�v���b�|6'u�	i�lc�ر|��+4���[o���M'nr��Pr���X���aǓ�%�����\��{�-�����P��}]yEd�av�$48)ƌ͑���r}�������T��G���Eeyfi4bAT���U&оAL^d�SPRLgG�n�κ�M    IDAT��
°K�w`�Y��&��	��y%B�B����#�&��-������@�K����ܠ_磏<I(W?pIY�gNe�3��ꢵ��1u�y���9x��F������ ��V���y�z�t�}�.�z����$��?��}����p�<���zz�qeeS7vu�FQUU��ꡃ�t������[,����@����D���:����]��ع%Uڰ��>td'ϪԪ6i��+)�bı�|I�a�vw�n�e(�uY�w�H�v�p����~�F�r2�0i�~}�DT�����>:E**K(�I�pk�G2�4�d�pk��+��kHw��2DQ7��p�3�K��߻]ã_|�Y½=�UOenݍ�q�|���#5ԋ;!2�(�"�q�))�g����)�!�WQ�XK�"�UU��l=�+�ʹ��ۙ1k�o�Ī�Vav��W\�57^�i�ϣ������Ͽ�g��[og�y��	��߃�b�/���w�g0���#�����Jpf�[�G^'�oi�%�V�z�5��4�"��tN��V�c1�$w\<�f��'9��^�lX�9�ס����3~<�N���ѣF� )@ֿ�Y�z��hnVɜ\+Z~�f�����@���x
��a3M�	Q�J�j�3Qd�U����W��H�1���+=kˋK4�>�d�!ܩ8�HP6������VTy&9�E�d��>�԰5,I;��DgdSZS�;��/� K��M�u��ºMq�����s�����hk'/7K�K�~�!�|���ҧO����JKy�ͷX�v��l�:��TM{NV�4��j����]eऌ�զèϫ��Ք�����E��n�S��M&q�x�}�=]dz=��TQ:�Jyb��5y*q����~H�S��U06p����y���"B���tK&շ��[Ąʊ��˙<������֦2//*`\m��z�[5R#O��R� !�	�b�0 ߓՎ_�a�
XD]Q�nؒ0y�D��n�񻬺�B�D:v����!6oۇ+��??��@��s��"/�����9��̛5���S̟9���<�~�%>���$�.l�,j�O$O~":�$-����lP��L�v���ԯ���Ŕl��I�!E"͠� c2lK$B�����c$|Ct���a���}'ZNp��!�LOAQ�O������ɰ�C�$�>!6^w����$�.�LK��x�4<Q��	�%�M	�Zu1q�����?�|���O$� 7���{59�ly�}*�v�$�,.��A"~EY�)���T�Giu5�d��mmMPP]M����������/���VYU;��w�p���������6�}k��3h�wK,θ�2�}�%��ӗ,�6�>g(bő�OŤ��5O݄KeZWȆ�F$��.�k}.G"�D�n(�f�C��߆Ϗ�zҫ���7�g�P�UQ��~�8L�rXؚ<f�/Y�3��feh�&h!J3�:pC**�NUC�|#=m1�M���I{=4�(݄�'%�.�p_Ý��)�~����bT]5�=�ꥉ�C�(͠L
E�#��\�#��?�h�C����G3(aՒ'1����E^������n��\oA߰���d��r�U�!Eց�F%��I�8�����d0e`x��L/e��*s�pt}=���ݹ[3\f̘��ISٻ��w���������áR���?p���>J�k���!&��v�NL{�d�ld������)����m�x�t8�"����A�gJ,{��4bL5$7z��D>&q�@$����Q�]�嗑�������l�f��w�$��ݍ��5B����-jx��s���F��X�X��	����J!&qrҋW骫��5khm:�u\ȤQu<�أ�ꖌ�p,�@����"��u����DXB����h�#M��=���5���g��Ү�]|1}�B|
�o�>>������
�6}��l�-�u����������3��	���-�78����h9|����|!��,��,���^��fEdi*�����ˊ'b��i4��L��U���fnYu��PC4�C�kA��'�׃�+[G�����j�� ����?�O%s��c�it1!l:^� /����u��ihL[Ӵ�� �\���̙����}���c[WG�`�/ȶ%��ekh�	[��aV�TjƝ�D�}2��OF�)J�jXx�"�k;��Y�j�_v1MG�9w�rz�U��h�R�X����ZE<�}���i��,���Fʪ*u2�r�/��=-mZ$�d����ST�'�P7N����	�Md/iN�T��N��"�\ʦB%��fP�/��0�� �v�П8qh?��~\Y�U�"YV}�}e瑓���/�"�ׯ$۸]v"�8Qç���<gi��D��0$�S:����4&�pH/⬜\��u�nQ�y�]�Y�3V�<��u���t��I 0MG�E��D(�*�vC������x�d��;0DQY�c�۞\p��̟;G�ޞA��n:[ۨ�8�kn��y�k�/��` ��?���7P0��KOg�eW���o�Ƴ/���>]��K�d��%i�ІB<�"r$qYZR�-$e�E�-�K)����lD�Ԩ|F|U��f��'�=y���#:U.(-����[�I�N�J^^���
����.� �WȐR|V.OX#��I��{d &��dB`&F��w*�ۉo�Y������^N�1�S&rl�v*�NfVV��0���^4�+/k^>-���=H_8��xhl��+ϴ��]m�)�=����r2��+�<}*ǚ�s�mw��P%�5��~�[��}�YSf�0zO>�WN[�X�e��`��7�7�k:�E�)e�w*��OQ))��`B���5��P�(��|0��W-rwk�]���}��y�S5���!���@��St����r�8���UVj�Bww7��eTT�������~� �zȦQ<�"ۗ��lL�H��H!o� 9$�V��1�
_!7�.D��
�(��b���ڷ�/7nRP��I�8���ۻ�m���lb��d�3=����~,JAlv`we�{'j
Q�_�����'���1S&c�ppݵW������˯��׿�p['W^{�����'���us���?�����f��+�������--m���rd`�)"�v<���*���Ւ1���<Fu�`y��b�PYazO�|���:�N��v��wZI�q��z�-PR[��)z&�UǬiS���f���<����i<JAa!a�b��x<^��	Ps!K`<;D��e�>Z��H$��Đߧ�{Ey)���&*q��&pƜٷK%��;�)3�4(;$͓�M0�{���,3��c���x�,ƉP?��Y�f��ab�D��P����������������];w��ۯ2m�Tn��v�Y����'Nd���L�� �g�y���.l�eT6L�~��q��#˔DJ��ޫq�oQ���d#e4�v��H7�ꢶ��Ðg���J%ɒ8���hoa�]�VW�bŹzN�*FT65�e�Bl�b��*@Jp)�pL#�,�*M$
G�f��7@�:J{dd�+}[,�#���-�1m�(J�ؼ����0��IuE)�旌+)a�+�1ڛE�'KAy�X_<��0�h"��|L4�Ryo ��pK>����'�����n45�`�R���F��J}����_|��CML�;_I��?�H$���c�s4B��Mh�K=�������wY�e���(���[�����	�?���#dQ��5�$��3Ue� ���������K3�l��Tһ�	Q�N{Je����������^O�$�F���~E_��X��h��>�򥁕̾�S�$�����Ҏ)$'˫��ʊR.[}	���f�?ש����� ��,:tz�gd�H�ݯ(@5@٠K�����c3h��$�o���+/`���呇��ւ:4<H� �mqx=n��I]&���oT�׺�����d;�21{��.^ʎ�;�|�g께5k�eU|�u'���3b��ƍ���Vi�-Ӛ��\>��S�|�\����B>��S������u��L
�Ů��ף^Akc!��H��k2M�&"=Y0�^���h>̚�c�?!uT�2}���T��_�[5�G�o�q��f�q�z�YIX�L��%`ɊI�~⍓I�H�Le$�����d|Nzp+a6��X�o�jH2jT-K/捷ߤ,;�[.��lS���2�����)[�H� +�`�Orb����nW2�<��%��K��IS�RUSCwOe��|�͜j�d��M�ܽ��;w�wm�����K���*��
���|�g_l��ބ''���,�;���w��C��ي3�P�{��9e0���n\	��Ogi��庼ՏmD&*��[�"2,�.TxE@6\'�����Ză���E�Ut��%�g̨:��[���W$$�-��̀lB$�A�Mq���7��w�d�4TI��.�\�i_�f;J�f�s�Wp�i�x�ٿ���/Yq޹x6�O��w�8��!�Q	���%~�`<�@D"R�����`��ǈ�_�3�C�p���:�>�<�������o�aB=۷����ݎo�G$��{�c��I|�ɧVT2i�t�}�ym6.Y})�7lP��w���5��K�+f�S����9y��^�I�$块�A��vH�e⫍Q:�Ji���F|n#�^9OE.	�N�1�����1��0�9����g%�W�:��*���E������?���S���P3s�&L�\M�RD#�E$)�����n.�r����{��cǓ��i<t��S��`�,v|����a�	DUB�q&�Aʖ9A�b"�7nf�zd�+h�`2Aݘ	��0Q�:Yy\|�E,�3M��ۏ��SO�n���K���[pe�����l�9�����/���o����Y8�ŋOg�����O$��+�'�.9��TT���pP�4�1.=�ÔЫͅ�P�¢Y��fP�A����<w��\
V�)���m�r|�6BmǱZ�dy\L�>M#~��T��h����n�V>�`-���@IaCCC:�J�;�KFV��2����Xlb;�����gR6N	pł$�!�%Q�9ř�OGb>�p�¨V����\ɖ�?��j�9�i����n\v+>ɠ4Z}AZh��|��߈Yp�錟8�m{v���a.�d'O�-ˌٳ�-�Q���X����F�_=��_l���cf����f��/�+ȣa�������ϫϽHj �����������%p\�GI)N%b�h��g�3#��AF$�2���Q@?rvF�������`��\��p�.�ug��g�]�ǔ)S�=z4��s�կ~����S�k��4�i4��"�QՍ��T_b��qB����:�G�~��D���./c�9�pp�.6�[G2f���\�$�iھ��T����|��E�O��O���`$I+ͧZ��x�N̛GM��<E�6f�̣���%����R��(�n��Glھ�������f���^�-����7�|��s5KO��2�'}����joe=��d���ɐ٬簼�z�VG�靠*3����"�yЍ���Ғ�t Њpx��,59��:�h=t���?�j��뫩������(/��E0��_=�ֽY��4<	�J���U�I��Whdk�;$S��)ep��x�C>�
IS����7ЫC��� g,��W����}ٷ����[{`X�'R�%�93��D��'�i�T� ��(����ꨪ�V����{�,���+��{wޮq4"?����M�y��/�2a�eW��5���x���ko#o��1g-Y�9gLf߮C<��i<�#����q�O��#+��l+%".��)u�T����\B���/Eip��3��jD+b���#DB~,��y�L���2�A���_m孷^S���93���b��YL�2G��c-����ZN�u��s�)*b� ���u���HL�l�+!�sa\�3��DUI�S�|^�-t4fRMu%El��C:[O�*�����~pu�y���S�m�X�])��`*J�k#n2��a%Օ�I�&��pgn��W����a.��Jn��N���ϖ�{X��6�t����/*��ޠ����.��L�C�^fL��혞eIg=����4�[�͛��%b)OCyb���C�F�¾F�\#�Di �C�����6��3�w3�ni�顀S�?I�E&���v3��jur�.����)��h6U����t��z���-��%4�Ah���V̱���D�9e���nv��ɯ~�K&��@�� ]�}�ِ����R�J0��˅�����ͪ����mhH��PQ�2�`K<β�gS_S��uQ���iG���X��d2"RP��m��Q�n�V�R&�v�d�#A"b<U8�Y�s5U�̟w'4�i�f��_z�j�G����7��;w���Ysfr͵W���tuu0w�<�P?��s�t�-�׍�{��T�6���L%ȃ#˫�l��$�bNU�������I�R��6J��р��6���OJ@g2�po;��v��ɦpƼy��8w��dge�??D� 2ܴ�����A

�G�I�ltԠ+/~,N��Ƣ

��WhlC\Z����Q�<K����̜5��_����l�<��Ó��koUP2"ø'��$tE�4�����d����v*�*���P�ɹ+. /?���n���K�����>����`#�Z�Yv��\t�*���]�\3h^��̜Á}�8x�����8]6���:B}�8��q{�q���s� Af=#@HE�
�p/�eëkv��-�T;	�5&��呐�Tȏ�jf����P1�Do(��T�WFf��oN�WI��C����2��fg���Ճ;#S�P�GV]�>?fë�=���_J~�Ӂ�REI���'v�X��y����7��=w�F�I�tpZ}�_�y�_�.�؉r=�H����`0JJ��6}�0G�ڵ��ͥ�{a���p����E���å�\��夣����M7k�z�woTĩ�ߏ���������7�+/�LYq)GSW[ǭ��ʆ������Ry|nu�sfxu��[�J�2ti���q�yI�J2�.��ߤJ�dj.�i���&?�J��H	�-bh���J�O�@eU5�P���"�̘Jqn>�Y˓��N����;U��O��G��$��)P�	J�&�����$��
����i��xYi�p���^�]z&��w>�<��Ǐ�J�HE�d{��t�������b1��J+�^
	�2rD�����&�����1���0e��|3y�JT�O��a�f����D�	���w8|�(���:Y��w�w�Z[Z��G�(qQd��{q���g �l�J�.� "�%��t".� =�d�#��c�@/���8��q��E|p��xO,�E<�����(ʲ��n�$�EW�a�ZN0q�d��'Ϙƙg/�MSA����g?��#���,8}��8��p��(V�G%\f	��K:�O�,r>ʽ���u����G����: ���eK�w����|�^���o��M�a��	&�s��.^��v a �b@�O�6�����AUެ�d5˖�˶ݻ��3���[nf�̙ddy3v<�>��ͼ��f���n
*�����o�^�uJ˪���8r����x28�����9�y�ѧ���.�k��WJZ��G`�
��Z�a�
���3��3EG":ds!�B���)$!��%�1aR�,�O�-Eb���_y��?����ˡ���Ӧq���Oa��ށ ?��9u����W�������7[ii�B)��1�DEvll�d��a��!KM,J`�__�n����Yu��;t�u}H(ഥs���K)������j3��5"�"be(.&���m��on�s�G�6-�3��;�<f̘���-�2v�d&N�ʙg.ջ�n3s��I�{���jl�kn`����{�O���TRUơ#X�j%_o�'�t�h�,{�Y֮�HV�J�H��&5�A�]�>�:i��7�B��$�t�\Z��H� �̝>�sͥ,��PK7�7~����d����RVU���᷌]C����C������?�U߹���*���~^z��{��    IDAT����{>K3�ʀt��x����$`\��b� ~�݋G�����
�w�t�\~v��	�v�v�s�Fm<����@$N@bd��͉�~���q�.�CU�\p�E,8m!�?��KϿ����q��|�n�}�}�(�]^x{-%U���O�e׮�<���'������؉V_|6�m<���l�l��j�Ǎ'����JBI�E%�@f�#[R�F�Dڒ�c7�'�Tq��7��/��h�#�3o�N�@d��`w{w��Ｅ
���j���9�ܳ�=k
��cӖ]����*1�v��<���=��'�x��{�����`S�j�&�#Rmt{�Y�Ikf�Ô������c̝6�	5Ul��S�V�~me9˖��QP;7|�'� �lU՘;�IĜ�/�cY�R�pfd�O&t=���٪�2On.�V_����Ee�1��+���oY3Y��
�J+x�'y��תfx����"^|�Y��8��x�/���q��LH�"��l��(o�,F($pD�`��R`��n�u��P(L:��?	���&0�������4�E����B���0��q�16�2���Dd�F֜�@��j�;��&=��=�7 ƔS>�$s���Xc��0��>]��0er]�����l߾�3�,� ��_}�-�v�]R�O<v�n�\�7�E���O&-D�j{�	��..��1�pL��X�3�,!?�˩#��5o��A��t-��0�z�)�D�WX����T� �#i��d�>P"����ӕA]m=3��bԿ��;w�bƬ�\|�J�.����^z��������I���y����x�Q�U_�/�g-9����{�~���4l>Iav�b���B^����C/�J�WJ���M�U�
�t�gDe~0�Ta��D�B��$��R�,� ��Z�62�aE��̜6���\�����(�棏���o1a�t�&ANKf�l%�@D$v�lV��L�N$�'�Lb��G�BA5[Rr����d���].\����Y��FF�����hw]'O��+(+�����H��]=hk�G0��ǕL���e����iÕ߹���*|� K��IYe�ʁ���_��Tt'�v�f��e�{�������㴳��3����'2�S�Ҥ)���;UZ�أ���?S 	v/ј��X5{Kf��6�v�2�*Υt3aıR�l��"�U��!\��'5��,�Y!2�vo'��V�dZM�5��g/���Dr���\u�U�_x:�f̢��Q���E��s���Ȑ�m|F3(�~i���ăa�~^p��L�����?����?��};����ªy3���)�MG	G��+���`�9��1
�C�a����mG�
�((-e��DM6�Z{x��Ǖ�x��._��nQ���Ͻ�K/�����_�C�ǟ|Je��?� 9ٹ�y��Yc��󝫿�?��?�����}՛�����"a�BUdr���Z
xe��oü�2��,H��Q��$'��c��jV,]�9�e�];���3O���2m�t����w�rFWg1�?�~���Y�����������������}/����`g��&�"H�*�@����������J�5� �\��"~|�M<���(J%(����S<LWw~��^����E�@?A�$M�%4���)(���L�ܯqs��+'���V��H�㑸t�s=/��	S��s'G����/�W�����m[w�{�N���r�N�ǌf������d?u�B�lYY�  	�b�����n�,�4�EI�#ͤ�{�!��_9.�!%�0�0g/�ϵ�/ę���0����?�Q��r�z�-�u�*!�󥥥�_��ٻ� �^~S�N�&���5~̛�}@vn��B�(шl�%�Z��{KI�"	�[K��f�sõW� ���^���	N�3�k/��/>��C�|I��NF2�5*�/�[��C�j�?��o2��p���E�T��覨��QŦ_�j�n�k�Gq���}hh�����?��N��럳��<��G(?U���;v��[����y�f��Jx�wx���x��O�/����',�(�H;m�r1�2S��e4��kL�)5�I���!�|�&F�P.P&�9�%�����3hk��@�I֯y��6�Wp�33C�B��ƛ�(�k�n�}��;��_�������7x���(()�)�4���p�&U�fe����H��
,̧EYA>W�����V>^����^�/�ɍ�]Ev2�_�2ep��&98�
��ٌ��gi)�:h<ن/"��8٠�z���ŕ��p,�ߜb✙�Y�����\k�����[<�����#\v��̟���n�]�����u���q�W����ދ���G~�ή!~����,���`�p��ɪ^/Q&�V�(,��˸�F�",2bp�s���E>���^iI�	A?�T�˗r���9�����Sw��ȁ��1c�,�C~�J��������u6����E8y�|�sr�=g.��?>�ڵ��
-u�8������&Q���Je��u��z�y�n�+��8y��o�����3fp��j#rl��s��G�o����'�Y9T��@O$������t�
;m��̝���|������U�.���݂'ӭ�������o��Mm4L�����ͧ��ש�8�y�`����*b*�~�5���K��)�4��	�-6xۼ9�`d��g"�b��J^�p��dD-��c�,3���� �a�y��
b�3̥�����������tw�c����>�a�RmE����mbq�KJu�5��h�.��<���?X�~#�WF>P-Y�{#��'��E����^�ڎ3����ǲeӗڷW�וe%̝3������G��L��NWg�������A<���G��^���D�N��ݩ��X*�1-?��Ϙ<e�p��%�%�tKϹ��s�e�U���(XM��cGU�c�W�X5n,ێ�`W/��"����&�?�����(�ަ	A?-5���(G����TEZ�,5�c8�I\N�q�f�Mb�_q�n3%��?<��e��0�����%Ū��p�Ŭ�;uڠY!b�k�!�l���k�*�Al�k�~�m_~ɘQ�L�<�Ҳ�Y�xՕ�D�I���l��5�_�,^�;z8�ܢUr�K�����4\�Aë(����t\=i#!2Q+sg΢ Ӌ-c��g+�m�KϑmJ�)\X
��B) ��
LN/;7��������v�${QhK/��l�IΚ>K�1����UL����?̞��x������_1�a������y���Ǚ:}*���}~�㟐���=w�����)'7���K ���W�ݛ��Д͢Ա�\��[�92}p4�] �V_0��s�Ԑ.TD���4�B�>i<g̝NA�xӢ���������S���T�kC�Xf�h����ǟx��׬�ꫯ'��L���lپ�=���\W�r��4uN�q�J�s\�
�}j�@X�<���>b��I��P���FJ�v"]�$į�۫�^X|�YlN��6Nq���vߐ��E�pz��Р� yn��ws̣����sf��z�g���~�������휳��_��{�Os��v�?�яnk�egs�����r��=�4C��ʫ�f�����F��P:�zS4T&-�	p��l�5��(Zuk*�^:X���<'3�����p�w�%��e��y����3��4���_���+.�@7=�}���'<��\z��̚5���~�jF�}�.���ߵR�mRhh���d�<c���j����x8d4�����/Y���Ӧ������,7���8z`/��m��m���M��S)����������:n����L����n�tw1(�'�q�'�0�9z�����tu�vs�5א�륫s���?�|��̬���}7~���&37�_���D������~�0�����.�����Ó���[�&����x]�d��VC�[t�:���4$���gVͅ��5
ҤM��� ��'ma�x����/��+/�đ���G��=�77���:�����;�_�����_�����q��՜F}̞o��>Ͽ���OR`D�o��H�Z<c�t g��a��t*.��Q�c� �`��n���_~9O>� ��Ւ��.>T��GB�
l`�x���76���O�DqD��93��0���������rgp�u7�-,!Ce��M�%��>p�_���|�s'.O����+���}���sx��y�kx��Wt���Ń�t�����<�5c��/aH�6~Ɏ聈=%�R�A)0�7��Qt�5#O7���y�4��8v���.-����\�z�����g����ii<���+��\���z�),�<>3g�a�M��ƛ�$gn�8�

�-*�[naǮ����?���(T(Mh.���k��d�����fM�P��hC�(���w;�c�y�7��_�ղ�BfL�ĉCi9v�b��йEY!�����:�St�<��P����[ڭ���sO&�Bʋ&�jo����+�a�/��{��Ũ��y��{v�?>������ڛx��6o/��1�����S����<����%���:�[e[� *2f��%D�,#�F`_#��,`c�d6I��D�X�ѐ�zS8�)�l�r�MW�����'���(���A��l�+J8５45W0LG{;MG���9.M՝ɂ��m��_��!�%j�nGD�Fܨ�Z刺E�B�����
�Y�f�:ژ4gF��l竏�P��B�[2�,_4J��%�t����M��͵��?V%Đd�ڝJ��0��3fp�7(�Y����X��?q�r��p�w����������?��h�1��V��Z��b֌�|��N^}�\�՘2����E��2 4��� �A��1�ڗE5!�c\T#a��=��	�H��̛5�ic����Zvl�������1����w����}ݝL;�q��G����-\z&?��<�ؓ����\�A�)�2)���������@`|!��+�=s:'����!U?m�4V�y��hܽO"I�ݥ��p,���OW(̗����0��@\H��e��Z�ĸH��}�����z|�(���]?z o^%E��,=�l�NG,��\���u�~&N�O��g�k��l��P"�ÉS��8JAi�1���[B)���iU�l�%��U����DX����eI��v�x�&����G��VJ���hc��]��;�����2��H�p��	�jjN4�0q֙�X�|/���/��P��DwȢ@8r'�?Bv62C%��&1R$�������3Ǔ�u������ގ�)���˖.������ޖN�}���:�{���d
A<�������R���9���i��!���ΞfΜ�C=̘�*��}����?l|N�J���\''��9�ڡ��'�V�Fk�	;��d�]RN����`5e��a܈��]�ʱ0|�25n�<iG�\#�����r3(.���n4��ʟ��4}�T���D}�$^o���&�>ͿH�J+vL$���x���QQ��5�j�S�����W�m�h�T,̅����t�8�9�������>��	��0o�\�L�Ĭ�7��ޞ!>]�����H�+�����4:���W_����I��N����m�����n�p@eR�JA$�+a�	��������ɓ1�sb��,��M�HK�n(�`�Ij�7����N��2�7�t"UPTB}�XfM�I]M=[�ng�gr��E��ز}'Ͽ�:}��4773e�.�d5���47�W���U��?����[n���~�8�w�NY�qŵ$�F�=ri��E�YQ���$�~!C���-��Ș�D�N�D��������s�p�U����utp��n6��X�����2u
߽�*��j4磏��c�<���%�(.������1x���y��wU�&��8d3&$Y��Ki���0��4$Yy�ՈQ[W�UW_ɺO?!9�˘l�MG(�[���c��4��cqszZ�'���2$c�(�|<EvN6�
đ��ŗ\B��qd��2i�8N�u��>�>��jjf��˸��+��?�\��.��������+	x��?�
�WSK������v�u���{�g��k��)iH�wTP*( ��:*�3Ա��GpT:�� I �=����{�����|߃㝵����b���s���~��<�ǌl������37sm��X���X������<�gp1Й��JI�ݳ��<:��E����O��=,[�׶��ˁ����	X�b)
%N���������ǒ�AX���s�������y�y�?ʯa<���9j0�F@��e���`�2i��<,���z����7������"~Ʒ^{�����dQk7IE:E��
����~�h6�x����A��Z��E��������+d����{�A�ρ��O��|�`X6�_��o���7���h����w~}�E���>t��[`wy����m߆�=�(l��Z(%³���Mɠ��U�e# C���&��=�*��=-2��1x�PD?s��8��?���=y6���Ix�%s��e]M-6��^.��bǎ����õ�e+���/�|������0 n�^+��E9+?7QEP)e�l���]��iKG'F'��������F<����a��S	L=$2qz���i���؝8pzc3����&Ϋ���ڏ��v�.Ŗ�/#Y���\��F�,����T�@6��s[��#�Q���V��'?@W_/}�i�=>�8g~z��q���9��������݊~��_���f�9���KyH�`�xU�(���rō��D�:%���d�/�6`�mw�de��rE�����v۱��Ǡ!�%��܈����{^<��3�����d����>�����^��j]��U�lhįz�O��7��e � 
Ѵ:�>ȴN�vI��t�-��{JZ��t�&|�S�����G��g�|
v�K{��$�o�������1LMMb6��U���D��9��v0��J~�&��&��}�9��X�r�~�]��xz�6���O@筁��ƽ_����`0;P1p�����ױq�z��]�"�0%w��o���vA1���E4���ᒰ�d!�BY�Τ����2?U���\ aM��(Is�8=t4���@:(	��	�w7����>�*
�-�ȣ�&�]���/���G����Ma!��!#`:z�q�����G�� �I}�Mf��$9�Ys��h���/��Q�PN^��a�g>�)9���L���k�j�����I�L�`,�a3�&�"��Hph�ͶF]� 2�r)���-bٌx���Va��u��7���Y�{W\�;|U��h�����A,.�������o/�����5g#�H����ā�ð�� G5B�x�s�44EV�Q��*T]*���;�>�Kſ=��'X���)�pdfa1�@)���<\�C9��D9�Y�*�I�^.y(B,F�ۅD<���i�S@�ò��Ƞ���w<��S��Q��j��h1�����h�F ��,���p�%��=����W�))8���X=ԋ�cG1v�@�<:�dWt��yd�:��%
e�1��bG���A��B��$�XFCkZ�:p�׾���#W�g�>|��o㬳6a>CF)���}A A�4�z3��F,���;}�d
��7�����(tV|5�Ȥr�0
(��Њ���D����A����f[�� ��\�mA
��#:=���*��6����M6����iQU�ߴ	C����bx��W���P��*[I7��AYO� v�?��� J&��Tf)��� ��x�4�%�l+(���Ə^���Z���8y츜�T�]���q�͟�=%�����#̅P�܀�� ��f���K���&ǯ����l��~�N��0�`(��6�;���F-�����= ��7#���K#��T	Ȕ5��������A @�>�,@�`����S�1f3m%���a'Oz�I���}�rC��J�^QN��͠�-8aZF}	�D�F��ę �S��    IDATx�$�AB#$NB�l��>X�1��[��P��:�=x���L�D.��HZ���%b���`YG���=��_Z������C��߰~�&�p��ql��,����h��[୮�����Z�����v�)j.�J��m2��g6҇�@oa�lR.'��dͭZ�
K��%7���B>8�b$}&%�\j��{�8E�7i0�!�,i���Φ�f�e�*�	N�7���/�MM���FS[�����&���;��s/⭷����.�m�߁��"����]������?�u�0���B|�����/o�����
��6d��e�-j տ�Ҳ�)/ʔ�(&>o�V��F-����S{y��3KI,u�.�x>������'#�I�����r�ٗ�S���ˌ��_ۉ�Oo�m �Rܪ��w��~���x�w�!o�-YI�)S�3Ω��\V���9h5e��V�����oދ�ǎc��Ϣ�a���u���%'I���
r:r=b��P�����0[�R�sesX`Л������k>���V�.��o�?��o�#������1�7�f�|c7L'Z��`��[�s�.���wc��~���FƆ�� .@ѿ�1L�"(,ȕL�C�bp�� >�����F+ST*�M'��;�;�k�B	YQ�����О\�L�֞��~�Z�����w�
.��⺵kq�m�Ñc�D��07�e�V�cw`Ϟ=�e�,�b��F�˷�+��7���YJ�8�S�X��)�M�:�H��w|����K/�TB��?�����K
��o��tx�TD>3J�)�&8�:x��%@�H:�`*��A/�<y]�S4:i���{Q�P�`8��>��@�z�9�}��er�p���o�eW^��`�|�T�m~�Lw�~�P��qp�!<������:�H�<�P)��s^|ě�i紒$_���O�$�����y`I�C�%34�B1h
�A���ԇ�D�˂_��S: �EN�%��j����~��i�p�019.�2#:[�����^چ|�>	!��;�+�M3+��7He�T5���rRi+�&\r�U856��N��~�V;6?�[,q�� �'�������T<[{7�;��NOLa&B�R�Mc�Sg� m�]E�,�a�T��؆�P_��N�hŁ�#?��_�'��P�؀�c�E硠� ���c�>�����D<Dr|/�G���X][/�;b��&F�d��c���1���we��יx��33@�7!�KJޙ� �7S������A>
I���3!Z]�e��O��TΒ�c�����", )�N�����.�t�-�Ͼ{���	��4�RZLB6厕�
�lJ�n�lp�������+�J�;_Ş=o	Y���lڄK�߄��v,LO"��ߏg����1�(vf]���X�r%�< J���n�����011	�ǃ��\y���������;p˭���<����t�`9|5M�
�1� �ʠ��-�Z9����`�F��P`E4�
�hmY�;�%�\Q�pKȢ�2g�Rr�Q���L6+﹎��X����0*�$��2>L�j�#����S�e�Y%F��_6�,����=`w�EͰ�ƶ.��?tDd� X+�QD��qA*'�+r6[�F���~�����Ub��g���p��Im�u-�G���6fN�B�ˍ��S����[�ޕ�pzzV��U5h�m���A`vK;MDpt�4��>�d:���V�>&�&�݊�'�q��w���c0[\�a�KާC���B�?>�0Hm��-`nrgZ��l�B4�<M�l�u�,� 	hL��8�ь٢�E�J3���'X(dE9�Ϥ$k��G9rI�Кhh���|2%�!f��A7�Ŕrp��	w�9E����c�ԏ/��x�O�c�>��)��l�b�3�}^�9��br�l��M$c���������_���'��ꦣ�}]mЕ�HD�����E�ECr�w�Ac�`6����땸�S�#"�79����r��9���wx=�9g9�"����3֞{>FF&���A�&d��VZ�o��W�L"���jn/���m@��Fg�a��`�:���2 ðJI�`���H[I}Y+��&ʓ�|0ށZ�92��(I�g�8y����$P�<���ۘ%^�&�1Qu�u�:y��71���w3�^8�5�5w@���d�?��֢tk��C%qv"F,C_.���T�\����v�2dY�z�LLN����hյ��(,`t�^���x�7]|!�j�&���p�2���=�Y�t:��Ǐ`xtTH�\ -����'�`$Bo��p���"·b�,�	8jj���K�̦��0=5!�R4Gϥ)�h��4V�:���v>�lbS�Q��!�.-�m6�f27_(K�3�U(ӢD[]����h1��y��5`��{�_6�:�d�FŤ��k����Ȗ�`3��P�<Ȝ6�SW��Ec����|�j�!�7r�@`3h����O�����^-!�D߳�ٲ��Y.U�� Aǡ� "����9��������鳷������;w�N� N,f���؈�'�"�aF.W��0��+�d�Η^B6�6��_�V��W���p�1��`j�y�8ͦ�aC�@u�EK,V�Y���#������+Ē)�x�M��>r��L����`A����Ї?�f&Y,�y�ɧpjd�]�A��r ��xc�6yQ��(�����I,n�XHE�es��YVCO�FB�dT3*�/�N�����=P("���m��m;��LR&Ԅ��wHZ��03-�p�G��a ,���+�:?�������S��r	z��tJ%��k��$��
�)3��<,�.��|��O��cƏC*��B*�Q���Tj3H��T "RÊ��b �S�p٬p�����[���g���{����
v�G������ӳ����±�'�����w� .��Rt/�E(����v�ڋTV���]��f����x~۫ع�r0�ꪆFg��H��V
V6$J��h�U�%�_i��`�ύW2,�Er�E�������a�;��P %��V,\�5��`f~o��&b���ji�\:��uF�:�{��Ļ����/K����JDE�J�=��eg"��i��[�����i�&\r٥�$���椙�����%�)�`a|b�pn�Cd+��c��e��Wa:0����*8N��6`�L@����z�����7FrA�>��|�>	q5����iD��28�~,#��J�P���vx���U�5��zq%���.������-��y�p��%��>���3W�l6#�cVI�&[�@�y��TFAI�P�T=�R1])����،x}�6����fs)�}�V>�������;p��Q� 2G�ς��ܳ�����f"��~"�/N�Æ\:-�d�t%?���s�(��g3�a�[��?�Ռ���?q����M���!�PS#"�Ӫ���Qt�E�IN���Ri��F8�g�E���hC�������&�j�126���߄�6��	r"[Ŀ���01uF�J��x1�E��Nj�[�u��M�1�������K����Ί`���*o�0X�E&c�ޡB��Y�"�ŗA��Y"��R� �K��$�p[��ɰ��yNa4r3C�(�_#q���^$Qy7=n����XUU~�颌����_#D��n�S33����Gc��(5���P���.*�K�V�Bģ!ɥ�9q�gnºu�p��qLLLɟ�lȶ�6�vu¬ӈ<��{��M�ܻ7�x�FD��5
�z:100 �V	�������ӧGH�g�������zW��_�J��lڴ$C(}�bAUg?j�[$�1<;���#r���68�Q۳ɼ&T� ϶RA`[V�Y�j��&��H�2{dշ�-(PHfsW)!+>X���@8�Bx�d�b0���g�o1�>a6�C2������Y���9rS8@5[aq8Ǥ��X�/���'OK1�����Z����-C�h,(� ¼,�u��y�o�z=��'?!�C����������^�j�х9��v>t>��>��0�������W`��1u�$vn{��F�8>6�C'�#���k׮ǲeC�J�cx�/O`~!�Ό,�$��O���FT77��@*������#�`��a�ԣ�s �O�C��Z�jĀ�`E*i��J�3ɡ.7=z��0�*�LH��,T�����9 pP�R#�<.�V�$�Z�>S�UH�|/']�T*��*g$���UNd�X�tw}�k���������G4AO"�S+
��ɳV��aE*������̌�~�B!�76˦�����"��L�dҡ���
Y��fS	�q8<^DU74J�Q��,�z�8���I��G���SԦ��Ad6#'t0T����CS]�&g0:6�߃4IΕZ�����vw���ˑf''155���!��>W$��"C�B� ��&<�h8(w�
%�ѳ�$��RɈ��N8=^�G��ω��
���J
#�1h/�OB�O�K?8
��8]���K&eX�w�^<JS�ɤ|��ʥ��^p	<ͭ��(i5�x�� 6N
oEFfYL���Ұ��>}�8
�\&�d=j
E�TW##�I3��+X���a��0�dBGg:�����D��%����$FGG�gb䠐˫�/���$ܝP<.m�+wX��r!CR+�U\Vh5������F߲e�b����B�iCG7��0�*�P��e�@C�(���#(g�H���b(�2P�y���N`x��Z/�zA��<��fP�w��zx�������h(-�b$_�w����ڽ�?�A����|os@7\z�"�&�S׊��	e��A\sم8�	~��o#0=+����^q��Xy�J�޳[�zZ&MD�3f��x���-�7���.�%W\�� N=&R?��b4Bᇷh2�X���/��'�J��p݇��k��+/>��{v#��#�j[��#᜔ͤ��g�H3X���ފم�PUW+�� ���V�t�K�JWW���[qrx+V�Fum�L�"<��G7n2����au�a�x�W4
Bk4���E\Kc�#������Ђ��Y�<�β�vO)⓵"�̌�DN�Y4�K�����g#H�J)/�|f���z��Վ��m���i���0����|�T�nق�'�ɡ@i�Q2:i�Z��n#����f��="0 6�e����ė����fqp�H~!6�(i�!d�g?w����O��^E"��Mkc=�kkd��/W�*���'�����}K��$]��l�u2�ڻj(�۰	�C+��cO�ȑp�}bf���R�_|�8p� �z�I��[*��u�S헩cz�6X�[�`5p���i^o������o7�^C��9�H�d�M۪���S$/��kQ��i���� ��� �JI���S��I �H�5,LԜ!�RyH�64�l1a�[�$����Z�+_��K�%����߀�M@l��)��[���y�TNjx���9�K�Gc��^���^-�+���x�7$�������[�^��5��x�G�w�;X�a��Y�u:�.��6�<.;~L�A5u2���e�+;0?����F$SI,��E��~���I��Ao���/���`�!�+������F"�2�O $
B��X��i��2&�� ���z��SF�P����5���(%Xm.��l�	7,�F���V��۸�n4�i�u�ƣb2��Y!ݓ�,N��� ��0�p8��R"#Rg���sorч>��6<���Nq��ʸrٴL�(S"#dH�^T�^�t(�T,$�/���m���O=��������-�1�ڄ]~�4��CJ�Vf��&]��Z�X[/���<��q%�������DM�5�j����lu�՝o�Q �,�yy6Ŕ�Ym05���o@򹢁�&'�@0;��oE��JT�v����@ OV����Y�ȣ.��Z�����(���#�!� �6��I����̡����`3�`�:15������.D���!�m6�\��Qȫ�S�T��j���"�s�}3����hniC���,s��P��̹b�w��hʝH�5u��G%�Ċ�>��ӫH�&Ul<	>a�h6���f��f��v���7����������bvj�cxꩧ�F��xD��u���V m���ƻ���r6�SYV
ȗ4�����w����&���Ø<qE�&'|�+Q�>��Pv�FMY
Z3y�п�L%������30����+���yE��YR���EQQ���{�1.N��-'�i��T�-���E2�C6�����q=���<�+�-�0�r�4�s����(����_���ԩ��2ĝQ-�T^�6�o���8#tѨ����%6P�@N�K�TpЦa3s�l`�K�b�%��X/�nvt�r��3طg�
�
����FSh��e@E%�{��PJK4�[�Fyg�-��:���
�͌�?��ߏc���‷y	z���xɀ}~�u'K�Π�! OH�)�]�I z��Z=n4��ȝ��d+ʻ���lh��<
�y�W<U>�=n�WȠ���ME�$?�N���ac~�� �!���w��J}��q�����o��m�%����e���ØQ]���x�������&#��n���n<��?#�C�/���!��
�4ڍ�&�F*E�r�r ǂ�QGu����k���/�ɣG�a��)DC����p��$�Nr����Ԉ���"7==}�m������,V+�V#"��J=�p���yY����h19:���3h^:��e�ŷJ�`w�$�D����)�éD*J�4cP���J��Mg��W���f�Kh����5#�EĦ�1�{�ȴ��௪V���� �bVy���WS�OJ��1)A�f���:}�Zw>t�*�SIt�tci���V$QL�`~���-���O�4���؅㇎�n4JP`vN�&ޗ,��L�s8����PY��`e,��ј�C�����6��r�͜o� ���R���K�t:�&�-D3y��uX�(����!n��>Y���N����r���y� #���RsW�R�1dc!�L��j�H%8Vd�pN���-]=�s`^fl�^<������E������{� e�����LT�L��͆j�T}N�H�M�ژ�MP�*��p^� �`�N=��Z�8zp�������<{��b�;{q��1�M*]�rf�In��$?�M_�56����33�$�q�U�`4�jI9���4�ҹUL�"0�]��
��]���
"�$�1�MFt�t����.;�'Ʊ}�k0�m��+���.�������ڷ��X�j5=�S'OK�T2�F&����m���loÞ�_����h�^���{�3lҠ���A.�t6%�JM"���V[U��-H�2� �N�H�㤖�䁗��x�*Rl�$��o��.P,� J���gP�|#�/���	d�Q�b�/J6��g����Hp�VPd�"�^>:�dg��f=������6?���/��&R� ���� К�[E^<Y&�!5��h��c͹��e2��/^�F���j�=>y����x�Ǳ�sp�'?)�k��8����صk��)9nk����LNN�f�a٭�B��s�w�^�8q\B���3ۭ�Ϥ?���*�O��</��\,m�sC�M�(�mB���F�WP�Q�f��W��&��Rj��j�q7�&��)�f��J0�rȧ�"��Đ��T8 ?+��$�q�0�S]\���A${�Sunh)S�����5⳷ގTF�wI�s:Uq� ;5�����e�l�mv��T�s�"�(y�tuw����l(�Iar������j�T�.rj�ϋ��^s�wށ���E%�Τ�N%e��������dF<�fqjn��j�e�Nϰ�f������Œ0�y1T�E�E6,�M-ȊǏC��('���=0�|p56�����ފƒN��l*I�sq��d2i�n����p�hu��_�3!�����9`*�c(g"@:J�+4VL�O+Bv-0��2�bQ9u��    IDATa��⑸0)8(�g�L�`s�e��!�+`�W���[_~Mν��C���$�`��ygc�Ib$D-ϕh#���_/[�&�	�p�f���3h����Ux睽�S���1 -l7|uu����h��G.����ocn����(�� �m� 3t����`��dG4�������PP�4y�Bvu���a�!Ob��)	�4�j��3��΄h<��
+�U�Q�rH��$����y&]=Fe-̶Zɑ4�<�e �MEPH�QʄQ�̪M��1K6��R������l.���\
�sb�pWW��rBa�B)^���wU�D��|��1���� L�zZ���B_o?�J#�G�֞�hkmņu砭�A�^�t/m}�^|^�CC��Ád2.>E~.<�$b��Szm=�l��.�{������m!��S��y���B9-�#%n���w�[�2���O,Z��MD���V�E>���`���G�����}C�1;5��������n�v-�b���`�ia��*�A,oq&�!�T���ڭ�����Q�҈��V�%R��g�J6�Ah�AT�(dc��̨on���F!���B���Vi%��A	JC�
�Ѥ�e��SN�r�"��Y�ˋ�Yi���;0�|����g�}�v<�O����w47�ʋ/�������?��r&��.�4]%ni�ey�XH���n�����Ս�0��M;~��m6/g07 ��fi�����˕P�fa�YQLgՀx*�:!)��軚[���,`)�Ո��4Μ8-[D�ӏ��ˠsV!C���(��l4���S(G��0:�w�P}8��Cc2��M�������Nd$I$�	�
I�N���	,��_��j�|��[l�lxgQ�ˡ8��h4"�ςl*�6�� �/�k� n��n<���xPS߈�]sZ[�%ߏ��SSTc=��C�hnD"��s� �_���g�b�љQ����O�,SQ�$�=���Q�6�jlX�^��l݊�Ȉ�5z6���j�=�h�(0:�S#^tə�hd���چ�S�152?�h%�h&�و�e�Q��*9��`Ezd�e?="��s����®L6ra�+�<r��<��q!�ڜV�(]՛�͍�������0��k�t8 �H͎�Ȏ�df��uհ���lr/In!�*�B�
0z��x�;�^�s�Sҷ�2��.y��{W��-���C��.�S#���[��㣘�v�&�N`�3ʴ�h���1'���*y�q�@�~�$m�3�c�߆�9e�޻c�#H����`�XdI$Y��Z)�f,�(���c|���*�3�H]�*-�A$0��lܸ�u~D�����"#�;�d�0U����	��.C�T,(��B2���Q���FTy\�3p�8�D ��a=EF�5Mmȕ��H�Ve��m�k�?7��m
�N&�_�A�X�8��ߚA�������A��y��"��[&�l�t�4bs���Pd�HH6�4yф�F�Qv��\F
��$yD�����Xs�%�x��ؼ�YY�ssB����'1����&��G$��<���Sg`,j���񺰤��tBds$~q�E�mSs���g�������G`��q���EO��3��f����ط�Ȱ�Z�
�q��q��9u$��SŜ9��os��a	���C�1��S��d��	���E_�����&�))R�4E���iRi؟
RP���h6�h������|I�Pds��QYI����8�u��3��f�E߆�j��O'����	��ϜMQ��F�
�Ӈ���M�ކ'�ق��^���������DØ��A2���AS}f��%�8�sc0P��	"'�⣣D�MҐ yJw���ϑ��̥l�����.���S�t:%���'���$��Nx� �H1����$A�99Ģф�Y*=R��)ޤ�NG]�ZZ�����Ia���쩆��%��2�lF-���0�M!�N!����͉/��Ҥ8��sNR!'N��gr9���ڕR	����;��$��xD�����ⴋ[r�i���Ǥ��B�MA�b���hAum�=���6�<~���,���	�w�w�4�'�%���V,C[k��׍�Ɓ��"05���d<AMN�H�JY�路�՜�Iލ��mV,���P�
����L�Z�O��&�l0Ɇ�J���"�#��$;�Lj�dH{����BH/
�N�M�tt�`�brb�dI6��<�]p7��b� �)2 D�F�0!A:@:��/�2��
��yhL&X�j��6�]'��ң� �d�d�T�dPxA�e�,�\���		�wX�HE�PҊl���֑�i�!�N!�&�l����5�x�w����6m��u�i�С�xq�K���Z�pY���Kq���x��g$����R0_��9��"��3� �g��" �4i�v�[E�ՁV��t�͂A�@��儝��w8Q�犓=��RWv2�b�*]:�5��p����ό�cv�T�fi�L�*t����@ ��CoB!�Bhv�D�L(� }�-�\i���9�0:�����ch���U�+�lb(<�hV�9.B�el��x*"��?s���ה�����bw�ӟ�Sӳ��/~+[��ϻ�_y�l�I�f����	�`h��_zQ $$���&�ؤq*@�"4�����6�@$f+����"�D�cT�}k�bj��Ѱ*��gD�*F����9��U�y���A�0�{�7��Z��I�R�k�;1�b�t3�=�W>[CU`v��ԃ��>��,��X��Bta^���
�p.d�B�Z�5���V��Ҋ�Í�F����BIq4]<�btV�z�I���f���;���L�fq�I1�8�N˹k�;��z�3Ϳ+�
��_MN����k?x���ڻͭM���#����^��kϕsk��۰�]�#R����q�Y��O�_Ҙ�A��l��U�@�&�
I��ko��W�����L����;�����	8�ډr�E� ���q�_,��\�pXq�(dniEgOZ��Q_�`ʩ={᪮C:W���F��*�F0ǔ��S�#81m$$�e6r���ppC�btl�PP�)ޙ���뛤����0ir�Ϟ����"���G(#T�p����8$-�Ϛ�@�ߔ7��qZmH�ȗ��Ƅ���cI���{��ŭxr�fy�n��8�� ^}�%�{�ߗ�?�5�9
�Ɉ��g�K.Eh!�o|����S�y��x�<)�z��d�B(��,x^�vU� ���c��2��V��{�2,4��נ��������a�I^5ښ�&3�^6�\(�SG��|a�Jf���]p����U.$�A<���ט+V0:1	c}��:U--P6
���">;��Ŋ�N,]�#5�1�NN�"K5{!�B�h²�����!2{�\��������z?j�}�'S2�� B����Bj�YZ'�L3Y��S��ϗ��Ƅ]Eo�����Ǜ;^�ѽo���kq�� &�O�gI7N��bja�/� g�x�/H\�Jif3�Z�&���K#�ѯ��F�݅V���phY]�G(E"%��RE�3�C~�D�\b��R���f��IA�mF��I0^�ބ�6m���%��"�Gێg_z���D� ��SU#j��K��B��$�(���%8g�g/���%������(^}g?���;�7�;zQ�xT*�d���`��5�']l�Tؔ��`2W��I�����*��Y��z�	M��
<����e��d1�r6�r:���PȈ��r@��&�ל�3t����C)�RRTs$Q�*�Bk8A�8�8����f�yx��'1>>!�ub^[[ZQWW/���{V�=kל�H$��'O"�L"57mVe�0�רg3F4���L���y�x���CL�P,��u�v�LO���F����ʉW�
���wN�$H�^8�u�)�w�'��*��V�v�O��B�dB!)<9�{�^Y��ųȂ��
}��|*�D(%�N����P�*��FȂ�?êu��̱TE%M9�B.�RZ5���a�i4�d��),5��[H}�XH����F���Se����}�+���n���ǳ/��ӅUg���V�����ѣ����O�w����j�>����G����'J3���(�"����i^���e%oG���-�`t�`��`w:�##�'����Lk	��a��u���˨7������F�,��Bs���B�b�.A���'ƠDb��?g7|m��W�#�� &�$5�R3S�ˤ���m.垒W�\&J[��[��M"��R�D*-�2��e��5N,�Y��6�4pڭ��#B�s۝RX�Cن�fU)��d?�(ײ8��7����[n��w��=��)\����.Y����<�Ǒ�(����̐?��*�o}/>���;�Z�+�sғj�@E� 3��'��,0*�x�a���J���SS"sas �r��}����f�n��>�yN��(�s�<0=ʜ�r3��Ao���G{W/��$"�9��B���RU[}���K����LCI���a�᭪B4�F���,�p�6���@cuC����܂�`��|�I�r�cV�	�[~N�yX,6�s�y$B	i99��;#���^�AQk������������:�{6���E�k7l����Ǟ@W�֝���2���_ੇ��i��*4+*�Щ�a�L�z�@��Y$=Ao�H6��R����5����L���%��Z�*[
����R<�8��ǒ�ٞ',��V'�[~^��z���6��p���a��i�N�S��͆�^T��nDE)#�#:;�T���44��6�vҦ�HœS朗M��Cm|��2E�G�$�(��tLd�TH8�ż;ҙuH�9D2�g��&��DnKe���K�(���9X��"����|����G?��w~�NLz��կ���_��06>
�^���g��Sx=.���;;^��땮(��寒��~�
*��}R�rk1+��R� ��
NO=ZZ[�l%�.K�ϓE:���n��F	P���A&���(�wnuK��x�	L������^6Ťs�X6���&��c^��,4�m��b���.��X��yg��������Վ��,���h@pv����U�'n'�n���V�r2�r`��4��3((	8�>8}ըh�0�M�q�����Q�kPКe����E��Ɯ�'���	����Ѡ����혚�������ٽ��_Ѵb���7�~+��o��7�9��}�É�'e�h����|e�Qo�Ƙgf��C6��s���,\M��T����:X].iJ���0�8���?N���-Pd�KP���lh�e8�z8uZGF�!��`��ѻ�,t�X	�ύ֖z�9�{w��#���<�3��Up�7���55u�������GB�����˗/��������Q�OL�'��������F��nX�UN&��- 9q�.���󣾶V
�3���0�dk�3��f,ԓ��4bT�d	�8#h��A�W������ѧ��#�3�]�w~�6��W�-[�j��~����o����l�J���"�a�+;p��!�T�Bo䶫"���K�P��?0�4ҷ�w�Rf��)���b����`F������(ƨh�5;dk��e�q{`c�O}-2�8�{'ґ �8��
�=="�M%��ƪ�~��_��E�J�|s�$��Q�ӃD&-w�����ga���Q��14�75��Q<���0�C��������kِ4N�^��8�ࡷ`s����5�~�:=��$�x6{�BY��� #�E����G)�г���7���.��W�avdk�����ة�ظitf3�C!Զ����3x��7���E�C$��ؔ�KN"�ZU�:�`	���>�!emE	��@s4;������M#�Sւ�LCֺV�M���FF��/ �p&M�V�K�CkC"�S����� ����؍��������E�.���<
\$��j��u�_��m�+G�`����O��:6��� �l�Z8��l�B�`�[3�f��D���fФY����[3�q���� �>�/I?���3(�E,ռ1N*�g� �n�tL˳�9�Ж��M��[�2௮F.�C��H�\n�l�b������4��UUaٺ����������8�q���G(9Bo_��߇#��+_�'���W����G� H�����JA�\�ްY+��\/� N8�"���_~���ވ��ŀUf�,R;�ӣ<D&%����F�eT�x�L���@2����������M�mHe�E|�MD�;|U0�4�,��^�>���F%����y���&��2(�9t&�d�~�xj9��%Pb>S�D��<�4B�͓�h��s���>�9��d5[QBQ$��xRP˜�0Zo���n������e�f�*�t��Е�x���9؏U�V��~/��Yˇp��w��ڄ�.�_��q��1��Z�g�hc�S#<�S�O�ĕ�;���8�ℇ����Y������f��d4&M����p�PV�@N!"�/��s���1��B�e����039��܂�AK�w��3�N�<�$�f#!$fΠ�ICW)�Ԍ�[��"�0�b�4E��%8=)�2YE�5%%�"�65��B`���*91/3֥��Nd!�vs�H��;�sxAɂ�l�����-w�-�Ư~�^ٰ�q�������L�o��m��[��-[��֎={ބ����"����� ����2$R��rY��l�T��4���S�Ɨ��Ѝ�͈���#˧7V�d,�y�6
.��JI7	���܊��Q�iiv%s�T���u����6�Q��avl�'O��|F�[�p�PR�Ȇ���� ��`u����hmh�_1f�<r�XJ��ܒ���GG/P>E>2�J2M&�2.�S���u9]�����E#�J0�LH�SH��p�������Ebj�r��ڏ|���o~/~�[>{�<S���W�r��ß�'�G�����?q#���u����x��G�P ���2j ����r6;7�Y�v�ז�f��|J�)yX=.��Պ2`n~F�rZ6�;4��1��b��7o�\ҏg2���%h��}���l�@�谣����z)6�|~���.�����1R�,A,6�Z;��ҍ|J��q��	+��U�Fw;z�v���M��B�����p��0�إI2�5���^3���B��BxA�6N�Y�0Έ����|P�9���1����b��	;�%-t�d��|����;095�����?�ַ��L���G���/�#�L�cnn_�򗱰���-ɏ��<=���qJ�+3�A���9�"�N�:�.'�3��pZ���6Q��&��>RL�P�υ���
ő�zoq�&�,fl�bS�03zR�O�ن�����K���uhp)�]�B����/x���ȋ���ъs�o���(?��kJ���c`Y:�;�I�i�@smf����/c�����*�j`�mP���aD�O���N��xZ�F�6�^�F]��`X�U�a��ĳGg 2M�t6/�h���	omF&��_Ӏ{��ul~f3^|�O��-����k����+�0?����|k�>p���z�_,R�F�
)�)�Oc�@��1�ot�s�@�H��f�,~N��j����fjgaQfȘ,>ۼ����@�Lf�l�,������Ӓ��t�2�v�W��و�'Fp��a�^������c���{v큭�I��]}�r�~�,LN�n6�}W_�5k�A$Ʈ=���hnm�������?�	z�/�2�5�Sׄږ6d�d���޷� �;�;��=!z�-P�G ]h����b��R��i�4�l�����Z�[�~�i<��V��~�/�7���y{/.��"\t���O�Aǧn�4�<�n&���(jj�rp!���bw����|�)���t���2��u�FR�%'�>[����ϼ. 4E�JyaaP�K�-�k6x=���;y�_ߎ|<���ۀ��A�Ѽ�w/��4�բ���>7�    IDAT�\}9�;��Sx}�[HW��jk���N�G�6����l�Œ�F��11|�|~�+Wb��� ����� �f;B�"�:=�^r�4v��yZG�Oc��[�C��݌��F:rBAn�KD��I}L`9��J�T� ���e��qV����`�T���a���`��Q��t���)0sF��cg�qzj�w©<^���z�f.!����)�e���F*���u�� ��4�$ղ䘟[D6�ZJ[s��n�͠A}��>��0s@K�etJd
�����	���;w����3����_���zt����g��׏�Z.��vX�N����8�l:{���"��e�x���b~v�_}V�Y��S1��w�b���(,�5��~p5���5�j��H&�w� eҚ�k�&�n�_.�����!.[,�ΫY ,��pw��_���B&!���l٘4���k�h�<l����
lD/�v~�l\��P��e$��-0'�FM�.�&�V����F��o�ȱ��}�Ǉ��߽�BY���?.�C�w�y�l��e�Wy�?S4E�G3#�z�%[rｃmL3��BKB$��M�����B��CpL	�`��Ȗe���Mє/�># ߺ�Z� 5@ʿ/��`[�G��}��O{�d��O�-�^�4� :)��T��O��MIv7m�R��c�V��M�w$��J�8�6^7��y�H�baί�L�b3��a�*1?��ED:���M(�Q���38v�(����?4,(�Jo�-�fn�ii2��*�:�����Bd�]RHR'�?4���vqm$M��s�9V�IL81$b9�-�F��&j�|5���ð�/Q������=?�lv�ww#��x���	�ֈ�������o������f�K�}���O?�K�������*>x�=�M�G�n�Flۺ?��������x=��.ϋ�ш%1��I�/�2Ӈ�	b�Z��4������`8�V�s,$��5�_�球�K"�#4����a���ò��0�"�#!�a��m�-8}��X^�itas"'7_���b�>�����2TẀ'#NZ"��?r�8�����'��t�EI�$_=D��1�~��I�[EwC�	��	L��b6�#ݶ�w"%�Q�d2�P(*�Sc������o�u7F'&q��?D�'��|�8���G?�۝���Gt�ߺ��g������-g���;_}��~.�G l��ѐ����n�g�n�ܨٌ��'�AM
��I����
�"��tZ�οG:�Г�,�X�*yQb�@��&�O���}2�b��p9P=r��������"�n������	�Ve��`u����@Xh�����q�梨$9^/�r����H���~���z��������-�S|n#���D�Cg6�leS�J>U~ a���"H�u�1iZiv�T� )M#�2v�[λ&[���30[���C?Asc���G�!��ݏ��:p���{��yCh�/��Eԟ9���Pz�t'�J�),6�4s�����kB-��7)��A��S��8�c��j!A�l&6G�T"����*�٠C�z�� Jڶقy��Zg�� lbh��L\z�v�?���/1�w ZW&�+g�?DWs�Y+)��̚
�d��"���Yl2�ޮ~���Wq��6l�tx�f�0������C>�Q��s]�����:Lz���u�j�p��9Q���j� �v{�4߾�ntv���z��|��[�ᑟ=���L\{͕ƣ��������ߴ����1;^��_݉��Y��ǹ����K�l��֖o�(���fR�ȡ�,+&�aщ�C[R���qPC�웂�(�R� 6��XTa����hO;#>x�q�y;PQY%�*껻:���܀�+����Ͻ��y�_B��%#3K�ω�ă�梼�\��[ZE���?Ǔ�7G�q�::Ĺ6H.�JCE%JKˠ�E�{��B�N�B\��Ó���2LE��mm-|ZZTJ�!e���C	M�ڔW�n�W̛:�u�82Q��&,���u���O��p�Ƶ(��ƞ������ۍ�=�4�\v)6���>��zase���zʨ��BB�i�q������N"P�Hh�iE���g���ymH'
G���4���MDVL���N���a4���.����.��e+��ނ���U�������W^�``w�~7ںz�ns�h4K�M�h\(��|\z�%h�lƞ�����\YM!'']t1JJ+p�m�E_k'T�lX��(�0�hƔ����;�<�\�\��Ɩt�E�.�dب��Pʦ4�4,[�J�`4q9t���P7��o�G"�q�7n�ѣ�$�j���ШLx���j�:A�}~���8,��aJ*�2d����dX�揲
�Z�Y��y�ҫqpL�L��
%^I<�N7{��QS�@�Kd�M��jE��*f-��'�t� �:֯\.�����Ãc$�=�8���p�7o�k;�����1A�sJ�`��a�ۄa� ?��� N> �����̨5�-�q��W�7x�}~q�I��V�wQ2�;�1�ф�c��cFefWW��w=}C�'�$U��7�z:�Mt�q�����}g�� ��ȫY�8���׮�!/ˊ,�C�|Z�ꑕ����ta��u�®w?BP��)�*�Yh��h�fTi�"3/������!�N��	���%?l�xnQ^e -ʈ��)ƙP�ހ�"�֩E��A��Gx��� CX0�7]5��#x��'�XWu��E\p���*�j���?��� ��)9�?Y|���4X�dfW#��i�V�Bx2�Lo>Lv+&"I5h��Ğ#8�7�ʵ[��d�Sb�MTɤ�z��Wh��-�f��fP�DxJ	�g��ݖ�j5)K^��(�<2DJ)9u܀b
]TE5	C�}�Q������P7�܌5�d�VDr�FG}0L�X��NpJ��`O+(�)9��j�PM�gx�Jb��u���������c�q���`��m���[�M��+.GAq!�ͣ�~��(*)��~����FHi�b��'��ӄjA����z���O�����J6�bZ0K$�O1h!��i��H�U��X�@\��D��!�Wa��GJN�b�0V-_����!��@
��*+��'�|�GCc�Cos���ɿI��7�U�0���|�f,]�P�#��B:��A���~�]�>Ӏ�VMz:�9�R��}�?�JqO�~#�%]�z����bKH���l�p ��z�-&�����4�dx��[�D���w��c��oT�g�Eai������+�b��j�l\{�ux������<��u+�̟��>���+�=Nv����S��25�ĉ��(X�1���7g���rR$�d��5���$�O	��+Aؠ$b�`1��?ҏζ�%n$�ܜB�[�3kjNJ.2�=�>�p<(TS���S����~��嬞5��lf�b��OP�I��������?@�z�t�6����a?��������]-4KR�Y���݋{t`�/�9��)�CE��kcB����������-��n���c�����bu�ګ�����ǼY�8���HKK�O~�;$�zx�^\~�u�����g����G���-(����xO8-DPJ�h����ʫL�?���%kI�����'��ZNˑ�A��x����j��ЀP2��m��\TΜ_�H�F��͍-b>�p����;xs�N�e7�DVa���a:W&���q�z�,�>�yr���3�+�ѕk��̙&<����`�`�xQ9�
�Cho>�����g�Y֦����-�b�L=�T�Y���P���/���';��m�ő����K&�?���Бϰ�wp��-(����SMx��7��Ȕ��.�
�c~<�ԓ�J�>��!z=�}>i�tFF��R(��� q&�_��f�WP�(_�|����+,uq�U����5�d��Z��m&b�1t��"2�/Q3p��@k4�D]���{�@UoEA.�/����a�w߽H�NMC��B+NCªX�bN7�C���"1btC�6��j8�.��Ƞ��73��ٲ?��9��� ��c��7� ��>ݏ�S�����.Ş6����B�Bɬ|�[�I1��]o��wޜB,]��O�����L7n��z�����شyV�^��_y��+É_y��
��D[G/�z�$T:�.��=}�I��`v�w�>�\�H�N2��[�U�ǔ�R����ƵH3+ɨM(V�,���0�kr��19�/�X�V��e�_)xOo^�uir80,).����X���r|���9�BcW���JB��ʵk����]l�&0r���Q<)�7����>?����l8
���ͅE�����h?z ��$b�Qy�ל�������V��s'�c������pA�։���@��m��Z�%˖���_|��Ƃ��b�ih��lō7^�Y���F�s�*A~��ذir�s��SOb��uX�~%~t����3WV"S��e-�V�=b1�:�4��JXE
*�k���TDRHy:��b��Hp�H[d�I���8�dZ��$>�,���u�?~DЈ��R\p�y����`w��Y�1??�l�*���w|u��fO�cd)Š;9��._��Ǐ�L]��=�Y��˙�͛6�K/�}����� ����y(�Y O^�	��_�&���gcْ%"7��٧���+�-��oRXa��0Y302���p?��U��zt���ס����o��T-=0�\8���ɃˡG�׆�3C��ӽ(���Or����)�ݪ��f9x�&��ȲNx�	�6`}��������D1�*cSH���H�}�]`^��8�+�|e�!M7�]0���:t�:�V��֬Dg{N֞��y5(,.©�'�	7kF��=O՝FSS�n�V���K���[6oC���G��op��\tpڜ������p�q���{�3��5k�_T���n�{{%
���QL���8;.<���g���)L!�����tp
29:4(?ۂ�sP]V
�=2�(�9�t>:xD�m�W��OK���GF��O��|F�9���)a�������H(�Az��k>}�b̌��3�~�;�72�ؒi%�t)^�ɽ� �:��a%YaD����%cR��%:���z8�f�[��=�hknB�̙������9�yh���g��n�3��{0��/�%N��\x.�N���w8-&�X��%e2�eÝԙ�b��0:x��=xc��۲j�Kb��F����������,!��H�R��TעD˱�3��A�I��W� 2�a�L7�	8Y���恠\Lv��7��)�d�D�UA�jN��` �rb�]-��*A���WL`[�Î����BCG&
��e@B69�SID���SHl�##QM�lۊ�k��g��n|��X�z�y�i���%������������E��
-��<
�ST�|h�b�ȉhJ%���"�!R�A"J�������Q�>,��eh$;���2>!((SOC���V�ŋ�o݊�t��������]y�W�Y-y(/>�<��4�Ȑ2����1��Yҍ8��mغ�,�R��܂Ύ�@͞;�O����x@ɻ��ɒl���G����E4�N{Ɜ��	�@Ć�-N4�R�a,�!z��Yh���~�9y;�܅��\����;�v���[�mCqi)�{�y��hκ�"l;�|�c�n	eq�f��vOp��֝$���MV2�cO�{ʅ��O
E?���g9���y�ÊT���2��T�q���Tz�h���a���hHLYn��v,\�g����(�R��	��"ZX�W=��S�����&�t�Y�i�@m͏���h6��+z�������py<���k�3���_����@e���p#��>Z��#:1,�&�w�!�!�Ǉ������8�:{��f$����L\VTQqGM3Y��[$�lub�ƍ�w|���`4�q�7����=شff�(���x|�f/X����E�7��y'j���W^��`psU�8!M��'��v�v#(�҈�1�r��P��O<89gD�zy�,�(�bV�P�F0����$�:�0�i���U�������Vi�=N�:�E�RZZ
�˅?���h�����=<�dj�X�b֬Y+�,�E%()(��;����&�������O���SJm�sYu5�A:�O#�OgA��Â4qc�d�H!��;�*M��t�%�M���gW`D;�7Y��H�5��'Z��Л�8w�(������o�tr��x�����/���G�~����"�x�iG��R�+q&�3�Yi�dY(I�{Er�W��k_6�|�R�#'z"*���HʄA�91a4�CA�S�1>���zq�d�������� ���?�C����^�����eK����?������|��l�R͢r��y�s�t��M�K01���5����G��⍗_CCs=T,y9�+)�,���ft���*-��t-fUW!���HG/���'϶33S\�Ҏ'`cn�Å�@@Xť�0i���F�hs�*e�t��R0mݺU�-���e^�����Oatl��~��D��:����8z�$�,0�D�a�fP��Z*7Lt�2�Tγ�?W	2�P�����d����p�n�.*{����r`�����<Mު�fb��y�:� ���/����J�eQ�|��~��{�0�r���'��2�ņ/���L<���YF�o2����b�̞�O>����x��Ϡһਨ�Ak�m���̧B��H}A�^{F
�f�`���v�	��]��ˡey�X3��F����oV��Ueh��F4���g����g��B��UX�fr<&􍠫�/��2r
��u�9�.Nw:����q�H-�z+Lf&'��3H-�hM2�8ݻS4O��dH��*������l�>ɦ�|֦~6��mDwk�i�Z�J�	����q�ԝ�=� '�V����Ɉy���l�Aѐ�i�UWwm�m.�6p���a��-�x��_� |�MM�R�8�.iZ3�iR8��8x�O�g��ZoA���-��*��^�d� v��3+�x�l4��J����Yx�Ï��у�ڈ��9�d�`�Bk[#"�QT������e�g4ʼ�+0<���yq�U3�4�V��F-z��p��1Mz�ƄbJ�c6	�I�є����(��"8�'��+�Ťx0(��i��jOU�*�_�|#�$�j�H;����Jρ(�ip;�0$�hiBg}-��C8w��t����/Z�Ysf��O'jaN3RI�*�*��DB�<օG�8"R����o�����#�O`l��4-� �k�Ķm�aʰቿ�©�>T�Z���Rt� A#��a��4�?ށ�:�%��#7+iiF�[���C0gdb<���Dqe%B��[��w�(�taVqV.Z��*�9щ��iV6,��b}�~0<>���+C2��}A�FP'4����M�1JK� �r�Xo��� 4Ӄd�5�E��r˵����#MD+�:3�����)M���(������x4�}�&�vu���Ø=k���M�2('ӄ�*�bEqI���|�g�8$�����?Â�5����wa��98w�6i��n�K�����` �W�~��\u��B���~�JH��<�F1:��8bu�F�u�2,Lhy^��avjR̅8�3j5HP� �	�2���fa&n���=� �����O��
M45�b!��1�t4"2�U<5�x�[)D�.i2���OBE9}��¹D �;O�[�R17	�No�]�����o ˗-��U���ۃ�,V�^��� O?�4���&�����c�G[��(��SLA�F@�ԡI(�o��LRE��DJ�4�q�Q�Ld�б��TR��D��~�&��� n��-XOS�W^��o���x����g�p���¡�����7ބ*�&):��9AZ�M߸�L���PRR"��[o�%�̵�߀�s���yＷW6$^G��Nz!var�_�y��	X,F��MB��D��3����H�fG��AĬ|    IDAT*)�tWT�iӛ�+#KL<l��ECkܞ,\vٕ01w/2�M��b`ȇ{� �sݿs�714��^{]��3���zId0H�l:�Ѣ_H1�k��TSf%�ozd.�Rjq�8�銖Nn~'R�gN� r�&�絍E`�?	`b�!߰D�x�2q˭ߑ�6�}���y���3Y��ߋ�7a��]x��ɠ���ä�q�_R��n�A��{�ڑ�v�d�IAq�^z2sp�E����	�<�(�TF�Y3P�p��D���0��i}j�s������H ��͒C��r���W�ynܬ!�3��tˋ��q�ac$�c�>���PPR�̜|�t�"I`���ؼ�,�hn5�����p�5׉KX �ɑ���|��?�+A�Z"�?��T:<� �U&R.yKJ>M����S�c��I�V�P����uM�y�l�%���,Z#��0����0�uX�|	��\&����C�Fc�_�r�q��)��;v���~�;Y{t���C1��Vl޼�f����C�D�	�WT�������o�__~o��hMл�PYS#(Kw[#F[O�����ߪ�*LL�q��4r�
1<8���1H���Г!!TLғtX�hJ�J$���ye�(����#��3|y���*�钂R�J:dss�؁k�\~��hl�b��-�t���nGi��ZGῧ	A��թ+C�r��T u�(5��y��r3�r�#=�T/ 1o30҇`g3T�0�-*��Q\\���Y��/�~YA��QO4��6m?��__��hs���q7��i�y�6y�W�X)�C�aw:��	��7��믾!9�ߵ	�E���.zu����:�*]����q���(�������t�	_v)�{o��?�ֈ�J�V��jOW��q���PY^�?>��;�q�����m���<������b���ϗ\Mj�k��Ԉ�^���Rt�[?r�H�8Z��j��xbR��/��/�B��ڼ4��M�t3�-�D�t5�;x�
)��$���I��z�D�S���Ѧ#r����̢]�,�D��i�g���rg����!���1���{|tL
1:Q�mvd���/i�o�!��a�
�O-=u���/���K��ٍ��� T:7��Ũ���Y���'q��D����QUY!��ݕ����J�K4��y'O7@�3c�ҵ��c,�l�0"�1���BeY!n��0mB{���<��K��hM��ͽ������9U���wx<�{P[�c:ApJ��J��,0_�&��~e� W���)�*)`�_�9P�ђ�J6-�]�e����+J��(����hqd���n<��3urv�_�`��%�'26[��=Y��;�2l5�D�<�ӏ֦Y�l\3l.���lTή����;::��_X��)zc�r�f{�qގ8x�O>�h�N��_�|�D����K���;h�A��53�= fV4�b��~� ;�LhQ6w�D�L�6 ��q�m7Jl4�����u��'#�[�H���Z�B���Ƚ2��0�	F�e�!^,�I{'-��7Y���*��bmO� �(u��#)z^
i'�� �0h΁4Մ��B�v;L�%���uc��}�Ob�e��Pw�Pw���'�DeI����%^����.622&��O`F�LTW�ƞ={0�7 Gf&-Z�͊IfyN���(��?�ġ�L9ݘ�d%��,��"1<o'����[H�E�6�mΒ���Q<���{�1����D�ܹBs�I��(F:Z�cM��{;֭\�����=����Y^��4AOo?#�8���b9H��%|�h��ڄ�d3�u�&��LW��c}�0���'d�(�!s���Njg%QɑVa���Q��J�FK`�}�PFQb�����P���_��gRK�w�hj�������0n���_�F�?b�E����O=����!�5� w��=\z����)�~�	����d(�
j
���8�ԁ�y����0oӹ��2M�1�4��G�)6���e0K�
��������9� T�?��*͠F�#��5����of**SD	�f�F�Z�s�/�,�O4�d�C��.�`[��-Pł��ӑ�㑥Ã���6�E�jH�6�eL�/I�~vV.��E���QP��kס��-��9+V�F~A���k4q��7p��	�q睒���?�	�}��aT	��5#���W�)�����N��C�!�V
!�,���2M�*J��6�9�����h*����8�.VU\���cdh��=2yްqN�����u�_޲�l�:��'"#*�8!�6LZ �gU͐�I�7'[�Xj�{�#	D]�p1�'����吲83������ێ��&��I�tj��6����B`rٹ9���ľ�>��Є؎K:����&���0@8�lƌ*�'�'�s�[b�]PT�s�] ��w�'�Z�ח^���[�ly5��u��*�__yE
x��R��	�t��܄����qHg���U�f�z#$DiH�P3؝���D����∮T��1l�Vþ�u#AJ�^���aɒe8~� ~z��xC���_6�;v\$� ���c� ��L0��t�u�3QZT���^��6����7������؟p�%����mDr|h6�-^-ϐ���uBq 2o�YP��ł�3��َ޾>�X���ػ� s��,A�}�H$���7֮^��dMͭҼ�[����u�nj�˓�U+�	գ��|��hnmǙ�,_�+V��`���S�;p ���5 �'�}ȧ�*t�	�{��ze���2��3��OS;�n� M�@7K�թ�v�e�Ok���I|��E`0�a�����fK�kO_/&��)-R6�:��r�u�c�[����]�k"���1���Y9�t��[�ttvadlB��=w~�G�z�=q
�=�,��A��z�����V�� �M���@A^<.����|X�z-�}~����=����,ڽ��N�I��ΐ�F��̝�m;�C�`·��C���T�t���"�47"5�?��C���((*G<n

�A����3��:)܃)�4%R�K�2�;�l��M���\i@�#҉���Ns������lX���$���Gd �n�9BJn
�%� �lǉ��gP�P?Աz{�1w�������E���!i�|�@�E�����}�������7���#4a�ю?>�4�4�������j>}�'�Qh�I��8q����MW\��?ݏ�I?/_�o�t;v�~j�9e3Q1gF��`����x7]v.���M��G{ofΛ��1ι��$7�E6?���gcޥ�&z1fIҐ+��tm�MXc��a�8�N;�.��R����8"�uJ�
E߯�H��6�2p�s8��83�cJ\c�>��� ������/�.|���h�h�֎V�2�p��Qc�HV*V�q���X�jj�;��Ѐ��Y¾`���a�^��^~~�����'�dV@o��k�ݤC{S�|u"���l,^4��j���o\!H�O���>���롶�d�2x�
1�Ø�Ea���vx�&<|ߏ�������w㩿���B�#a�����I����'���[~z-�*ɑ��6�,1퉓ɣ F\Rl��L�>L7�B�fk��4��7�x2��S}i �0�� �-"�6�\cDI���@s=��f6a���(��D]�i����WV�v�U�d�݊�HT������d�G� Y3�g�d3�С�2�������[���A�o�������2�f���Oa9rK+�]��w�Dtli�48m騩(��� ��2�q�X-�����RcbJ��KQPQ%T��6�,jT����K�Ǭ�R*��I�����p�`p�'ڸ�d�--0h�(��|e�F���'	���%��ꦿ^K|YSH���6������MM*5�S��
FiN��|E�N6��5]i�TTFD_S=r<.T����zh\���bB�
��e�I�G8�?8��;w�������8��3EP5�J�襥�X�jΜ:�d4��W@�7�� ���3�fVcՖs`�{��܆���i>S63���DiA6��v8mv�~���'#��#�L�l,Z���}�h����1T�d�'?�N�Q������d#̞L�M��bpp}�mХ�c���SK��!�aK�R+�,�#����O&�ʕO�J��Br��W�l��)'�)��O�?��?q��cF.��8��d�@/�F��D�������n���e����C���|�͸���0��rv'�8|�O>�4�~�]%�,݀������ �9�x�'����������T��q1u'Z�������Y�09��Z ��Q�E��>M�@a_�d>�g3(W���7�j����j��� ��!�*�x�h�̏i�(�%�`�!©�T�Xf�0�ٌѶF�cAx<vTU���u$DdrRB}�������@��Q�]1`Qi���AAN.B�	d0�/ˋ��Q\Y�O�}�g���d8�˄�fuﻹ�C��X�t	b*���b�P��'cr��CQ+�l��I�d��h6���x�æL���WY�B�J��iK��(Oq�b3ȩ��i�3:Lk��N\|�%�}���=�۬��fA�����Ç�v�ZY��<�,��A
N�}��<�=�2\�V�>	��//�$��3Ͻ�ΞnHϨ����8&CI1�S�ݚ���t6�F��aF����,��D�9̨,�;＇�{� �`��h��h�qv��C�"�R���av�|,[�
�}���1���[��&3BBM1cf��|�J�g���-��J�6MIĔ�&Y(�����g��H��n��*�!�\�ΘF��tH1��)8�&�3�<���C݂��c����ؽ{�o���ķ���ݚ�(..��n�k��&���!�h`s�P^V!�5F�Q����+�G~�+���<���j�3���cO`$0�م��Ű�4������t4t��(-���JK
p������s~�>�"�$������#
 �0�c�q�����󫥁$*�n3㶻����t�"���h_o|�=��&k��H,.�Eu3��̪����n��~*���]R�uj�����&�%1�!yO�Mm�r��X(�3�/�h���}��`$��$��	L�H3�)�����0<�8	�t� ӕ)YLŖ�f�J�����Q�z����FMu�t���
����b�k֬AEE���?b�NF��kG2��.3%3�i��Bˉ�PE&�n�!++WLhw���bnu5�;~�����o��Վ��R�����bt`X�}}���{qյ#��¿>=�o~�G�U�KbRGww���p���U �ɉ��nq����0�H7ZS{{\�,����0q��Qa�(SSy�^#D��W�V�q�4�?~��S�^PZB)|)�KiVE��mdb��AMi.F}�̙3ŀ����������3�N�5�Ӆc'k%.���҇��R�ڜ9sd(ȟ���N�###�x�R���x�Y��Ӱs�;Oi��]�����98y�0|��@�*M6S�^��}�NTT���+�6n>u���e���]���s0:1�X`��
\F\�m.��2�� �h�h���~fk��ш��EttO&r���4%BC�Q�lh҅����K���%��??i����馑w��	�2��>E�O5��r�}g+��h��#�����<U$(�CSz:6��Y^/N����p��sp��qEN�Qcf�Ĩ�{�!�twKsN�472u�gT���Hr9�d3��� o����f�<1�����ށ �*7��9X�t�F-��N�ԱCP3��aŌ�Hө�l�"����D����^�o�stM"��F����	]w*���UHOL���q<��������I��]�O/�gn"I�h�{�arhz�%��%& ��n�u�S�[��M�}��U��I�{�P�R� ��=��3JQ3�xM��9YSB���<,�=��Ϫ�.ި�<��F1��,�\�)���AaY����18ԏ��l���M�4��Ő������K/�,��V�Ď냼:f����{�Ǣ����ŌY�榐�a�s/��'�|&o��<�΄'�cC�8�B����� �m�������w�>��᚛n���AXmD傥p��9CiJ�C�� k-�M�]#N�_�����o�3���a�uf�vl�o�*D��y��� c���V�|�N��f��"]��d��&�^�I�=�0R{}��7���qC���DrS�k�Ǚ��=�r	"��Dv�.��D1���}���f���c�7�@( ��%�Ÿ�� S���D�i�Bb�]���<���6o�矏z9�"ر�|�G�GQ��/̡�<�$����Ȝ1K7m�>ݎ��n��A��cH$&QUS����k��A�ƛ���?�<%�F`�-��������@?� BUٸ뎛a4������F���!�q��_d-��]®�^�X�tr��QG�J����\�0MdI�D'�V�IL���[�Ƈ(qJ�/wZ�_�+C2��3"A�:<��d�c�����Xo�6J�J�j�2�墻�����bŒ%K�t�2x23�����g�^a�э��R�z�r�2446�_－s�>K.��5���Մ��Z���^�@0w�,h�n��y�g�b���`'�X�}�"�P��� 5����L��j3�^�6��D[�:\be3�r�Qt@ӱt$&�4=�P fU�=m�l��AcZy�nᴟ�y#V�X��(��w�s�8y
�ta3Xa��JOK�E��Y��u�],�9y�o��w�{?��i�m=i`�`i&�����ڔ�0�֌&��Q	����6e'�2���P�H�M5�2���IAyU�'���qs`��4�h��� B�j�^�F(W�CJ$@���V-�fo������N�n��c�� (.*BQA�4;<�C̟��c��M2�ݳ�3447�3��8x��X�f;���pg80�ۆ��#ШC0h��v���|����pYAW�_<���һ0X�Hsؠ5��KbzZ�x�]q1�q����=�`@c�Vm:�e3�1L��? �a,�K����:yq�op8�A��+uL�y#r��V��)Ek�)+)� �嗥&s)���B+V�=J�)V�lE��fP5�P�F�����Ѓ�g���u�0<<,E���ɲQ�C�Lq2���)�zn��Xr@$�N����7���55�6�]�������)("Q`�ق}�K�ƙ�����\t7���aD>��zdfM0��[n�y۷@��#4�~p?���Pm0��� f������R�� +�,���a�p��g�������q�V����$&&���#19��(�%P�!D�[���b�Fg��yi�8M�t T��w��R�=mޣh��i
MJ6�=T�
��H��iJ�]�i��?Iy�$2Ȇ0:N�0��**ˑ��-��-���72���^̝3G��]�v���EWY�)d�&|>鐷n�:i>�w�7'Gl�kkO����R�vt���T�B?� y�3�!�A��PE�Og�ۛ'b�4�~��X�b1>x/���h��Ee�,(�⑁~��/��AOkn��\w��`�'q������G�'�3�q��gP�c��^��9hjiD��`����%��n�Y�F����Bz�.�Ra
��h�=T<ɛU�j?]i�,d�9|!�M��R�FFI"<�ܳA�q'e�NS�����v�W���1��/IgK#�*JQTZ��yZ[۔}/��Q���_u���;PWwJ�"Meee2]��o������ԝj�J�[���K�����Z��4A��̵��ـ����;����ڻ{�q�v��a̩�ɓ����M�%va^E>
�i�j9����]~1z�!��� ��_�R�aN���	�1�?�h� Ԯd����Ĭ�	_@4�aê���1�GY"ʫ�/��:�7N�2��:9�� U��\`e�)_CG=�6�D?�#�x1�dp*O� �t3��˅2�f|hhgm=K��,^yVŧ"X��h� ���2?v.�Ct�t�Lj�p��P^9C
����Jα��!A�JJ��%��f��X    IDAT�*{12�QSS	�^���3��=!�+'��l/��4TUW���܂�>ؽ����|
!c6�s�#'�D�E��i�B��[�����ȯ�-[��P0�w~�G�x��2h�f�t���D�o@2F�3�(,+��~��@b�x�	��(A4JTр(�}Z�as?S�uW�EF�P�f��"�ʰ�S\o"k���h��M�%�d*"��0\f�)�vu`��z�J��ҋ��?0!��\u%rr�16:��FFF�����ރ�����F�$��t�l��p��������E�����O��/}z�9�ς��������Gp�_� N�i�55U0T�����? �׎/N���K��&@��B��5���1<擳�ț�ަ�(�rㆫ�DQQ��?<p���/��.F8�B0F�7�	��
�����Ye�1N31�)0���k8�ϥ���ti6	Jۗ������6�<7�^��KqD#QDB�����EC�[g���DV�1��PW;�{g�¬�
�ֈr���:��W\�l�WA`�>���̃>���V82\��������,���1Z-�n��݂��$�	N����o����AxJJ��/9Qn�C#�1<66��j
�N̞U��.ށ��|?ނ�zt�E�((5�%��?< %@ڿ M�K"��,'�������	�s���`v;�*�4J�$�>��;�@q*�D����0������|�4&DL=�d�RO���͠���1[����+_�M7��'I�%u*&�FZ"�ɱ!��u#:��ǏD`Sý�6-�Lz�0�,fĢ9g������<�E>�mm��������s�=#���++QRT���+No.�}q���EH�����+�)��)�^�v�OA���+,�(� �AE%]��wd��f��J�)S� <>�b�/\i��4�]�ړ>���9ՊaJLa������e#3Â�+v��]�?I����y]���mP���;3�������L��� �!n�b6nZ�����j���G���?@fa�_D�S� �r�yPz�Cr���v|�XPp�,����R�)H���Ø�4�|em�Z�l&R���*!��F\6��E�z�0t�L~H��A^R\�U˖��1��l|h�B�������ߡ�4l����)#�.R蔷a�Z�.�b2��P*�S�'O��vct܇O?�\���!�E�N��`q�����c��]g��F��D4���m瞃���E^�}ø���⍝�@o�B�qÙ�%����!$�#X�l.���ZT�U���B{�Vm�Zg&��EHDc�'G<@����M�B��TX(�5�.VH���M62�[ݯP]֭�<�Kj��_�{l$Bo���n_J3)���MyZX3v��&���F��%�h��X�l	֬^#����^9fp���7��=��;:���C&6�\�4\�������[���ѻ��{���	�(/�g�����L%Ҡs�;c\<�h@k�a�S���)]���ͫ��oǚ��D�|ם?�kzG^8�J$� �E�ہ9�8�/b!?��;ؼu���ַ���c�(,�-f(�#Â(���2�Z]�pg��$��$"D�h���S��\){��+&�3j�5�
2��s���cX����
N�ke#�c���.bl�� T� "�QCZ�;˅��R90o��6ij��
�sӦMR�^r�%R��>J�^�P`!Ƽ��/�\4 \��f�"!,^�D�܇~Xh�>>�h��8`φ%���b��������qMx��PP��D,�k��;�9{�|�o���1L�{�L����`3X���5sg����c7��|z��{q���Ôڊ��9���3p'���T����ΩFs[���q�|4�HSҙcf�zJ�R�)�"���ק��t)A�L�?�4kR6#f�ݔfP��
W��/���b�˜�6��H�P�(�V�_�A��J�]w߃��>�&���3���6\t��hmm�}�j��^�<>��ƹ���C=,Z����ΚU#���s��q��	'�л��YT	[V>.:��~d�����g�lҋ��w�s;�/]���a\p�%hh���EV�Lxظp@46����e��3��&<����.�Ƴ;��#�zJ2��4�����"����w^"ց�+SЛ�bC���9��q��w��,���kBh�
�+ma����-�e���ٗ��+����Sb�ETP+nDɝ%2���
U(���
l۶M�)����1܅]$�.4�B�z�p��1<��_bdxz�V"^wCӠ7��v	�{�W(:�pHд�"~�F����n6�0@g-DNa22���76<��/A���I��c7����������҆[��u-=H�K�;s��
����b^u)k?ǡ����߹�\w5L#���?|��(�1Gbc&�a���b	 ��E�,d�A�_�iD�8 �*�Ñh1�V�o�0��9�bz&�)ĊяҤ(�j�h�vu\�t�4��;�X����0��y�Ɖ1L(9��	���R��e�d�ǅ[o�Y��r��iq��i���+����a�a2�����J7��z�v,]�T��8��Vd4B:�؊y�V#��\j6GV>��������;Qej�9��ø���`A5|� .��Jt�w���E��ep�`"�a�\����h�g����ì�E�{����_�c�����i5:�G3���m�F�,$�D��o1b��f�o!�9�]�fO��_3��ٷ<���|Jq]�!I4*Y׬�H��L��j*��9yS���1�Ɉj�B9���:�1��b��K�q�=�7tuwa��Om���� M���J7�d����555�퇕�/����p�D����N�i�s���L����xD�1aú��1{f%z����� S!��A�t�j�<����"���n�K��*̬,A �'u}ؽw?�l�FYS::�&5���
S�'u�´"M�%X˫1�0⚔�48��j���z��G�f��h��ԍ2�O�=�%��R�G"��!��6!26,{aZďɁ.�b!���i��ɏ�'�ը�ſ����9B�L� C3T��h I�t Dww�02̞U��M%$��h�@{_?��:�'��Dr*j0w�Z@oA8�Dh*"5��jJ����@FaQɹ!� ���f���z/�/��a61��-�C�����c�I�����C����aeCȷ�cv�:��� ڛ�S��8�z5ϫF���Q�n��3+��1�/�u��Hj�p�"ӛ����jd;�%�Ц���m�q)Vo\�]��������BS�M��bZgw��Am4��E���	�F�NUH�Ѳ	�R�*P�47Y��+� &6��NkS� 7���SNj�`e���!B`t1��l�/��W^)E��`��L��!q�o�G__�L8=��%qZ�<�˗/Ŷ-[��p����E��N���oJ�Ʉߏc'j108�P��{3TiV�8ݙ�[��kG�q���br�W��4�9��8���q�E[�a�%YzV	�0����g���բ%�F� �Ī栅sF4HC�-���A��K/B��-ӭ��|WUVf���_�ս����ٳd�<e�23��������+%�»ރ������`g�06=?�L�Bh��3
XZZ������{��ƛ����6��VЮ5P�ϣI]�` �xbdTMt ���\�F���I�cu�Z���3.���K6��tOte.r�P
�3�`�Dq�ȼ&~�2�Ho6Ƞ(:lB��`��Av�Aq�8H�0r�����,��w`jzZ446w�u�'���_�<���V+F���j�M�����4~�ޣ<9��s��]����_z�{�P�wD��/\@�܄7�Ar��3G�rok/|�К�����9|����G�[B�_��_Ǉ��/�H
��2K�1`���>B�>��7��K���O�{��:��O�쐅��?>�������C�?(��j�9o���a'F��kN/���U:���0�s�Фm4�!�=���Љ&~���y�aj�L��U�9WNU���P F��lS�לF=j��,ۇ��e,,.��|������	<s���v����]�'�)�v@�=|��c4;;��>� ��ַI�Etv�Њ���77�$��,��h�����-ñ�Hf�HN"hP����g�	�Ã����<��8�B)��GV�_y��}�C���/���\+|�=���s8�4����㕗��o��o⻾�A�5�塇��ߔ��l�	������n'�Rч�|å��.�M0��aF��K�G�2V��G*�t�]_w�'͉?��d�_�V�G�74 N91!"�U�i�4�;�s@���luq	�T�j=��I_I�R��d��͛����t�|6GGF�~�;'ӄ���z�Νŵk�Q.�q��)��ޏ��=r5x���,Bv�0���2��~�%l=����,O��H�c��q��������_�Co�|�߀?���ٻ��E�I�ǋc�K�5�����Z����[���hvZ�_��NC)$t����eD�'m2�B�tuf�F�
��T��: 2�0��M�2�����I�O�R�?�<�֒�5�O&�P�5dF0�����خ���#�q`ukp*E$�q�g�1�r����׵nΜ;�:�4ъG�:�^|�950^[9�(�HB�%
����&�Eu�K+��qs��nʠ&O�t`'��tVȏJ~O}��v�9�ˢ��(v��^��~Ǐ!��So���؀7����waf�JՆ I�M_x�1�S}���ފ�>�6l���+HO, I)��P.���i���3ʲ9�stI5$�Q�GS3�������j��ԕ���ȉ"���-$ *:h��F���6���IS�1��V�^G��3�j%�rh�+���	��򘞞Ɖc�L��بp;{�x����:
!g�K�"�"���Y�~;�{�W��f��F'�Y��_��Yh���0ҳ����7���u��#��A8A<���;��Vp�]gѬ�{����`��06���w��gQ�UP-n���	o��n���׃x���V<{~��G�"�T�U �0M��P�Y�Z����U5��>�i.ׯK�����L̄���� k`�e�NT�{J[h�G�����p0�5׮W�(�S+��i��44D�t�4EN�I�ef � d�����L�$���µBJ=�b����;=e���Z^Y��ԔL i�Fpp���~�Ծ�;㳋x�[ފb����=�:r��}�[^D2����coc����D���N�����ZA����b�V�A������p��Ń2^������l�Qm �`w���Dp0P�5s��_ 0�A"ut��67n7�r�� Q'��t�f�fP���[5��f�@3��i��<v�]���	�^ͽM�K�XO^\����I�<2�I�fD&�C�b��Yg� *�b����vTkpύ��:�3#��.�@;�(��z�6�b"�6�<|�?���l!邉�31w����~��&Z�;��L38����M4L��Em42U��N�\k尸��A�%�$f������p�y�bA������0���ݧ������sh��x��^|�e�'��-�FC~���8�[������U���q��I���O<{��D��{aR�z(��h�(P��Aʎ�aq��}�P��l���T4#K�ҵ��X�����p/����BW9�K1�ٰ�9�1\��
�]�����Z8s�$���7�Rv�ps;�+׮��^�Q�� �'1(��ܴ��Wō�{��/E����~����?���
Œ	,��Шw��+�Xv�����u�/�&��7���H�����������O����|�C�˿� >��HSs�6x�-�;��v=���K�,/���v�}�]:�_�����|	#3��{hTBy�"Ϩ^?�lv�\ƽ(�j�hMF��l�����d/C"�]��TBb��uh�c�M�ۮ�2���jC0��ӄS-��(�&��h�����7�K9vT�0'g�KB�>�w���e��ʈR��@��x�(9�jQ��!�l�<�˿�AD8����X�9x�#B���Ie�4���K@%+�E"R>��T�o5��������|�?������":���#'1�Bhw�X����<��W�u󊴋?��?�;�<�w���^���i��u�k�
�6�p�Ds�'�,�Y`���a�F�k�ء��wG�.
n8�nn�S%���H���y�Ԣǵj�Z�mN�z&�;��Z��4d�R��kr��7>�N�̙�r�L�8'���>���.�b�?�jO��8����3�L+�A]D�y�Y�8�з,L=�@j��ڎ��x{ׯa���`������͠K������_�E̍g���><�������.a��)�LM����q���q�'Ы䰰4�w��_Bd4������ƍ,�<�v��գLN�P�p���UoMN�C��j�H_�ڢ����u�n������`��D+T<AӠ�^��j~-�1*�w���P�H�^�kĩF�41 N6A�J���φ67 ±�bx0�s������p�ڵWi],�y�l������3{���`rrR�m~��F2��'��Z�����`e�p��� �ʢXm��t����xA #	B� ��J������߀�y|���g��8<�0�+��?v�/���$:M��M>��,����ƹ��¯���F�o�����&�+�1,;�D �fqʭ�����"�O��A_.�w(�YɽN�Ow�4l�L#2̲���q�Ԥ���3����*>}4���nT�kV�5~��f	k���[�|�/�g]��P����D�@����?�%j���q|�9Kgj-^��=��d"�J�"M��Hsw(����W0�t���z���v���{LH7''�h�H�x�HDl����,:UF�X�1ӪHzf7�����8ؽ��{�������ا�(���(f�
G9��Fb}4�Ԗfk��ɟ��+z�׎�/e�)8�F�G�!p�%��Љ�]G-���Q0��1��c��rz�jj;���������ZY�LV�#0��(N�Y��!癘L$0=1)����Z��|� #4�/�M5�]��k�0�C�S|�w(��)��(�T L`��	<���
�N�_~>�Dcs�XZB߶�N^/�K_ݺ�"666�����?�p"���]�k%Hgv� FG����Dbphr�}L�Gtd~2�g<��6�q����q�Ru�~���l�A���ϸ�w��l7�J8qq�!o�m�m0u�=�QW��f�>�\gN��GtKy�[�#�&��G�i�=Ra��/�N�](H���n��fj��06��'[B�"a�t5e��z����^֯�C1�=��^�z]˽R�� k�[��Ǿ�.��1�����n��ԗ�5l2�3��'�3bݵuxZ��p��뼠ɧ&�]o#�(*��ʓ��
D��Y�}a-�z>5�Ծ�� �|&|�z`�׽ڛ�6x�4q�"Ș����o���7:���S~��f� [W/�w��!��h��N��S�����Q-���bٴI�~h��MW}�0��[��C��P�ȟ��4��>�bu����I���<���������c�Pn0}�4N�� ��@�y�O�w	�'B��F.���2�)���@p�δ�sh7�6�A���z��)݋�]�j�\}淛AW��m�|9MN���߃E��TL4�T2�O|�cr��ɟ�ILNf�?�k�/#25��Y�@���8�����6ׯ�Q��g���_���|�K_�/�G$�=�R �@��>�����s*�s�
���c�l�Xȯ�!�M� n�UM�)��q�4�sX�p��ϋ�̈́[n�D�|,jetK{�j�Xt���IY]��//,c��w�~�&z������=��5=aAL���cǑ5��8E�O=�,�ꓟ�#����yLN�b{����*���HM�F�CJ��u    IDAT�m^Ge����'����e�Ǐ��8��.�mO?�M<��׀��ɌJ���P]��;�
�x�1d��j�X|e'���Ϡ���o�a���8M&r��kE�9�����3@��䅨������!��wj�T`(�N҂���o!z/7f^C�Թr��f�a���YЍ��P�D�^zM���I�WQt`K�gա���'�l��=����jlt\��C������*�&�y�9�lF�Y�`a~	۹j]sGn��O"_*���~(���HS�Lg���Qowqt���\|�)|��2�������SȌ��r��뗙�T�C���ޅ��=����n�05��z���
��᱀�dbd(���\��7��+�V��ƞ��LX����,J�I�@:�H:7x~�~
��Xڵ����8�v�,�-��i�����y��dL�V�����r�e��q�3+J���� � �L��"������-�.]���cs�8u�=����G�,�.�����O�^�ǁ'�E,��'�E�����a�,/~���(�o��\X��sp���$V����U������bcSx�����z��fk���ctA�ۜXp�N-�O���Tr]��$ō�'"������/��u�TJr�㔂&l����0�z�߳Hj�!�\z��V���~�ڳ���ߏf����#�g������� ���k�Z.�jʆ�����5tE���F��- ��Ҹfiq�X�R��-��T�t�*jN�f��C�=|�j�b��)Twr�|�%x����h�2�<���4<V�l �q�����e���0s�4�S��z���¨�j���хX<�"c�8\#>]'�C|��ܲx#r۫� C�IK����4���jbs�L^�V��	 ?��3��~��p�>�HKOW=�{�}}}���T� �~���\e��U�4�Zcv��Z�LtH'��48N�ibLν���H��{황��xf�Ucس`�Bޡ��#�e� �̑&�0v"�'�S+�Qj�d
W=��ړ�F�I��ɳ�:~*ݞ�+{(n\G��G�Z�����1d��	E����H1���T,�!3%F��Ebl������m��MD��4����-6�����y�F�׆Z]R+yߚ��9.$�0�[��5�����[����iN
E����}��� H5D6��r��v�ǣ�	�0�kl����)�4��4��;�\6��X�Β3�޳{����i]� e��l��\9��w�'�_���K����E�]=���G�&����E���-=�9L�Czz���#Sz$���Vm��GE�fqM�_&}hj��N^{�s����+�7��Եd��!}>�?sa���G��"f�;@��:#�l>뮏2�bu�(��K��W���-�zmj�kU$���$��`{���-�v����G��� �)�s���@�V��r��=Q}��'�F'Ǟ�0��?r��a�{H *���e>yV�$��8/��E���)��r�)^�X@�� �R�V]��AӋư��(�����=/:��,�~� ��k������=��`��5ݮ}tZ�h�*c�FQ<v̠
X&W��JR�.�����f���kd��F"D}',���u14Q��'�v� �W.���#��O`<jcg�FSq9���Ɲ�.���Rj������]R�	��Zu-[ ?���D���hP�vX������R��F��Zǃ�cg�|�N��(jl�{59�tv7@������LF�Eş��M�G?}$,��q��0��4�=�ó��t��L3��T�ߖHܫ�L|������&o�����WP߹m����Ӏ�?'\=����2x�ŗP+��ЃD:�p<�ѱq�-,(y��:���6\�;��֯mni�ߤŸ&�,:�vD=������`��N4]�o�n���>���I�������;�:��u]����%�Q�ӆS90�v@�9�i8П)8'���:�T�f��3�.�.�M��n��7�L�{�%������g�����_:/^,1��#�0;��^��[k��\=���d��������Ǉ�"]it�H���~D�֚(���a��0����a!������ua<̘?
F�����Ɉ��8Y2�I|�ìG��Z��ɑ{�}!��>U��P"M�=��l�\�<,i3�����M�y���0�H$��սd�q�Sl�����Q:�	mr]�x`���Q�T�6�C���U���	�姥�G��P,.!�A��@�MG����_�^���6�GxtZ��v����W�+����#96���,<v��������E�6�&�W�YXBbj����:Q���~���덠Rq�:�u��e���_��,L��Q�	��'BNě�?A�_T&�r�\�Iw�������(�{j8p�b��y�hL���7l�8��;[54���ö��9�N�X˖��&͔�KZ�i}�������24���f��=� S25���81%;Cj"����=jD�C��DmwkO?��e��Z������;��D�+�p��������4K��b�O� J7�,�6j�&"V � �F;�mxCaX�Q���M->Ģ^TKXԘ��h�IK#c��A���46���h�xfY�yEc�WM�ؐB�'e�42N��0�1����j�}�V���W#�&��%��!��}�{I�hs��{�[OR��o�A�3���4qޔE�r�"k�����;ұ�_e�C�A�l�dǜ�pXa�c��9tHڔR��f���~�_�4|�c+�<��@2�NÃf����WQ�^C�`[�՞�Gvv�sG�f�/4�l������T��B��xl]R�Nv���AN�x:uP#-�o�K��4g�%ז�͝���1�F�h�Ƣ]`��{.ݐ&c@�n�)s�s�2�Ho㴀��&���
��1��r��j"��0�F�ZF1����ery�5���%�tSL�����_�9��ɭ�jY̱R1d�v�O�`������d��݆��!�^��3�_���9�y,L?��3w�����ˍ��W}{��-r��L`|a��i��o7j�wA݋b�h��H�F��m�{�2o�c
��XD'sUA^Ǵ/�^jz�e���y���:6Od8��d�zN����(5h�TBy��Z���F���'\�9D���kԑ�Gp��ӘM����v/>�J�}IWTz�rH�ќ�:�U�b�{�'���#�ZM�<�� �ha=�g�\�s�3��G(�� G ����!�z}�s����(�|.0:�̡�H�-Î$���*��!�2v�]����s:��N�&�x>�:�8�f!����j+h��O��L����0�5��*�>�FsGX+�5�e �#��RLIBa$D������￧���V�V�A[�e��a �G��և��&��<<�&�,����Z�"��
��6�q�ʅ�H��|��<K��D��Z5��b3����V�ǈ�?�eb3�3,X�AG����d�Fme#��_=��a�U5ה`��-��mD��ZZT�1����w�`JPh?�/ gnu��+���:��>��~���Zm�1ݒ^��0�!ņ�l�������̃��m�젦��|s��5�>�k�g|8H�v�)>5�օ9ӴRl�OȖ��@���/p�F2,�$�^>�(��H��q���^��F��R)�3����4�FzX��f���|H{���yk5k��xt1���:Lb`-�Fa�1�^t	:�1��x,T�l�a�̝h�쩦3fS���6��͠��D�[�����7�}lN%B�h�"r����fP�>�Z�� �'���k�P��&�I��Z/�� 旗T`�V�W!���)V�G�d�&�B�t�-ƹ�������fB+{�^)�}��O3	����\��̜(��j\�ګ�W�3�5_˝rȍ�Eչ��JĚ�,��#�͂��^5����ؿIg�R�6Ŧ|ڹ�Y�y�j�U�4!!s:e�~��Z�چ�zq�Y��p!���k��Evb��q\�|����E��M3������u���W �xvc�cFF$��m�a�48-k����Cj|��2�ܖ�U��Q��(�h
�I�ek�F�L^h�l\@��4Uc��jl��qNhY��4�5�C��.&c�h
�o�zŨg���zGR֐&��>��R,<`���z�#�,^w�-xpr8ta��R���n! ݭ0̐{�W ����/��$�\W�(≔�����՛[h���#��[(l��.�����<��f0�����:}/�s��F��t��~����(c�ȮC��A��e8�|� �HM��>��=?���/ .�1�m����1��1�;!c����w!u\�ʣs>+,~L'Y�	��$*!�	9��>�r~�gN��q�u���`�Z�����m��_��	7������V*Uѥ���Q���Ў[�i���s2P#������_�Q���b�Ԩ�.�\��x|~Nyu�P�r/>w�����v�o���~�$�12����;�\F�c	a��o��wNi�nK{T`|l.���1^��� �Q�᠇z�R�0�=/�|�D����B�[�m
�����)�oF�k�Z��2��}{����&U�fC����>�^8NS�#����[.��݁
�>��^�8�z�p�dFXX����ށk_�׾�Y��yM�≄(�,jMNޣH�٤vO&�>�w�k�{��p�p�TU���Ez6'8ԴRO�����P�up������B�?����?E�� �h��H#�<�P:���,�݁l�)�8ظ�^��bӗEv��VN�o'Ql��������#HC�5�a�qR������6i�t��ٗ^�g#K�^�Qq�~���&�;�:�!|=�_L�����x{M4��M>����W���+�Ӭ�Z�E��l6}^�Û�� 6�_å����o>�f_ �H���P��H)v��<����L
������K�7A%M)�z>�f9%�0�|د���|��0>��/��|V�#��~�%�j+�D`iU&L#S�P�P��j�{�j�ۚVP����љX�4������x~{zD����	ԏz�!�!ׄ�o����T�V(]�(s�t���
}4���v����ɵ9�s�w��{̈́��s���黇�C�%���'c�4��lf��ͦ ������{��+ؼq��^9��h���ܯ�ő�G�I���_<�����[��2Ւ�� ���yu#�ݑ=�s�0v�7� ��Q8� :�b�)``�);�u{(l���u�bX�9����x}�����^y�i��)����G�(���:�Z����폨xf#�B�H$�c�82�CӼ�#���@N�8�0L�V1$2�w�llޏ��-�6��b����铉� ��3�X,��q��s�{�P�l�ٕL�V��n���ˋ����A�`W`:KvE�5����݂,.-)��k����}����M��q�yasB�8��Қ��RK}��<��v���Ju�*�
t�M�aJ�R�cX9����	�����R�@{A�R�����Q���Z���̀���H<�xƠ�;:�<:���8σA�B��G�������H��m���DWƋܗ��Z����5��u��%s�Q[�<]��#D"x}r�g=�cd�A�����_Mtt,�{ϝ����k�5ܑ�g�}L���}��a�	|��{j����K�l:�w(������_s�F�P�!zt�B�u��9q�g�B�F�C�������(�n�¿羦���l������`�H��� v�LH @a�aQ��Τ�q-��1��Z-�]Em���C[xm"�4���fƴx��o޼	�VCc?�a[*�E4=�A8�:s{H��4�mF�D.��C���dqsJC{z.��@�o�eS���R���paz�oO��^	���0_�۾�����)
))&�Q4�qx�[K�Cc����cQ~��2�� y��M��EO�UOR6����jj/��'�&�
3�U�N�Ԁ�e��NT����"�H��S�oS����<��_a,�\���=�h���ӳ�����	d'g1>� ;A�PA1��J��;ۀӅ'Gpt��)�G3p�U�:]���ߥ�#Bp�C�&|���4ۆ�o ���6�C�]+���4D���ʘ�H:�h����6���	�c�I�%��k�Ӹ�8�5�\��
�m�=Qh�ߠ˫	�6���j�x�����];�6�>��b���T�� ٩Y��AP����N�=�׾����h�����٧��>�1Q�����sr�MLM!=9�H�\tN�m6�h�o�^�g#:����2�XM�Pj5��/�W�j)#=KTCR-C�o[�4��^`�����Zc�44��e0Z�oSUL�ɶ��tO�Dj�ddb&�\K*��f?�;N
[*>�	�ᕍ!�}���.L�]+�ʋ�hC�JG6f%�Ιq5-ZKx �S�xB_�c�0F*,���Z�,�˰,�jj�#�f��PP�bGN��ϼ�߂# N�������?�Wk�[�
\�;U�c1X�i�̭j��	fN�v6p�'ѫ`�C#�Blt�E�d�x,Tk�=��;@��j�����q�U�!�a��;��C>�]cx0�᷂r���VH}�i��H'�3��,�]�Ds�5[������N�=焄��?���*�>XX,탽vao�JA4��o;���/�����~A�%\�lF'�g�F\s[ ppl���0�k�7���O��Fϖ�B<������\���x衷�o���ϊ&=��F��`��-��e Ѓ'B8����1��1I��u϶^����&E���q����G`%�(v[�U����i�<���9 0 �#`s��)MM\=�
J[f�iHo�'�����lP�B��Ϟ�P���=�tDCbSf�Z4���?պ��k��1R���&~=�Ť�k�����X]��3��v77Q��6�I|<}$�	d���|�5p�ib��@+�"\�����b�G-�04+Q����8����+�'�Y��2^�}ߋ���w�#����/��ƧѯTP�?��k8xF��-.cbi�dJ���tPٽ��˗P�yhu4�_Ffi>6��{����(�+@�}�&���&pB��\L7X����̲6���e�<cS�����Tnl�E�A2�G�J˒�1�D^3��(K���@�BS7�b�0kg�_�J~�#�Xvd3#���)\y�y�8���W������b�f#�(�\�N�bҭi�f��|N��HK���\& �%Z@�P6d�����[A��#���Q�2��Z1��i1Z�ܸ�6�^Va�Y���"R���בP�v��5ݯ�6�;���Y����ܬ���MN�}X��r>oQ�yA`k��w�aG�2DB�A�`�K�&�Yfےׄ���(���ϮFMSxR{i��󗌴`@���;h�R�#�[����Y��!M�b�H�h� ���M'�G?o��2~&����#f� ��>,,-Kîf���%'��)�A	I|����4�z=h����/� 9ԃ_DGgp�5�G;S�
��r�h�K������m!35��㇑I����ϣZ(�Vd�B_,����UL.-�g���k`� ����|�
y4w�Q��ۮ!�I��c��{�A�l�.%(�0E�<O0�����������=�Q;`��gC](�,�p<.����؅Ҕof�����ڋϠ����L��q�}�ql�]sM�j�Us
c-c�"����2>�����nj�����d��}�.�l�-�o��s���]��k���a���?}'���9t���@Ԉ5�4�B���d؀"�A��j��>��Q:�^��d��;��yW�#{]u���%
�n�������ZQE3��dV<��ظ�X����p��[_��ӅS�K���N!6>O4�rg J-��c�j���B�hL�j˥%�f��'/��L,��P� �
w��*��oI��    IDAT!�
�j�ZAi ��A�1t�p���3w�( �E��d�1p�#a&i6��]��9��B��|^���q�+�����$��6��^��1FUX�kNa:�����6w�$P��$p�=���ٳ�GC8(�	�qםw��>���f(}���"u ��I��'1�{@:n�&Ji�tN:]x�A����O"���
�5�i6p}��4������rE��z'?n#�:t�PI5�1"5x��v(+{9X�z3wjG�7]C#�CL3�a��POW��F����hG��N��A�ؤ�R�`�4�T)<.�C�� �.B�QD�<����( j|�^�}A���ESj,���|�"���$n��6\:�����������(�G#�DT�)���xF�\m��/�W�C�é��W� �G;`��	 -�u-�j�"�_߇#,|�^t�l��F܂�����1G��CF�ڹ4����4�9g�(-2��<�x��Ճ'�
?W���*��s{�?>/���,�iC��s'�j�y�k_��]�6���<,/)E&W�L3Z�^����n�$���:����؇����X
'O߆f��R���?����ب
���
_�£��'���4M;7���Ԟ��ZM�bra#�)�O+�<��쬿� 8@ǿ�h٘���'�x��s���h�=�����~�,�i4�x�bng�+�%��h9��Ӈ��l�X3Ԝ:O���?bqN���fs_f!B-2A6�Њ1#p_�T�Ճ�A�Z5�E	�oDm���%!POCsN�:���K������5D��W5L�f`@�s��q�%l\D��t���ch�|��y��id mM �x��tiAXZ]��~�O�ӟ��q��mh��q�*[�p6��h��#�Y:"�0�º�*ʢ�]B3�')Rv౉y�-�?�@�Qe�'Co/�i-��HȆ��<Z�2�v�n��Wh5!�����n�,JÑ�(u���
�����-MQ��s�!�M��<KЅ�ۃ/��â�l�	��i�l�9��C���"�S'#��G�@踫�M�15;)]��q56]��Z� ��ROh	�l�ٔ&@B�ú�,��� ���_�7��b��çN���^|쯿�O~�8�zT��z����/�Wi�"�fih��p,�H$L��W� w�
��� ]\G�ȬAdj��(zlVQ�I ��@Dώ���k�T�*FIq#x�Ꝧ9b���	��"��3Z�ғ���h��q�%���>��rZm��	؈��:6��Q�'��0�H�e��C�R1�_����ȤS���;p���q�������S��'&Bˇ`$���U5,�i�*s>�)�Fv�?�I�c��O6�f�0Qn_.�=NobI�Q�biDF�1����G:1���Aq�n\|	���^�$2�G0:3��3��\袼����/���O߇��8&12=_(�V��M�����	���THS��+�Z��SH��J=&���ާۻɋc�o(�r���#N�ٰ��--.)?��%����P�/&�A|dD`��A^��n.�΀��8
��p,�.5��*ڹ}Z]�L6�G��Y5�d�)�� �0����5�mafi�T�L5�0u��8c#��}N�ոS� 0��c�"������4�������{^�F8����ڍ&��tܼ����t���1dg� �PÑ��Cnk�f�jM��C��Df~Vo�d��}b�X�6��� �ש�|��n	P
z-:�+�HM�(w�ƍM\8�BA�g<C:���߮3)�F�h��^�h	����>#F�?���Q��!����D�RW_x���e�x����Wí�뮮���>S�V"��cvq	��T�L&���?t���Q�-184!e�Gm8f��B��>��ʊ��P�1w�Q�� J�L�/r�TI��@�4�Q�T���L3H7�H8�H�,D#�4�p2�P���<w�F��E�!����`M�A�����&*�i�<���	إɈ���uln����ZUQ���"5;�A0����BO���A�4Ua� H�c�m���D����G~;����t�s�K�!f�`��\L2���Ͳ��A�k3ԤG�q�i�F�f2���򛩕aT������{Ny���qXχ��D���uǺ��7�m��ИF
oW��'=яIR�&�qs{hF�ҽ���Ţ����)���ލ��m���|P��P0����h��7i{>� 53��̌���(�����%��E���I�gD-�[��:Q��ЩS��B8�C�o��d��ɫt!.��r9ή��kE������($u�=�=����m�Ȁbd��
�D yr���4�"�5��8�sZ�Ԋ2�����{��phJ{a����{ȩ�
VWK'#�����0 �O�ҹ�=�[X�?C�XE|t�@V(�r��B��Tf��������7��a$6¡������9:��a%b��M"�����8N_�eŝ���\G�PB�퇟M��2�V�K&P����h�*䕐�,�IYk��oWEq�������������"]��%u_�w/�{=��UћԔ��%�m�u�{�&f�͵�5i�Ȇ���:�}�9}fc�n hyp��1�J<�_�>C�?e�;>)�BjE����_����D.�D�MS?�#�Ab7� l_�N�=�Z3�I��ہ'���x��'�gyKs�z�(�籱Άp�ZI�7�̸�,R�s*�$������:��T��
"1���C����CJg���N P�׮א f!��I����4�-�}��eM���
�^�o(�X:�i@�"FF�u�v�F�O����	��Q٦16` :�ƶC��H�xJq���]]�C��
�n�_uv;w�m�����'���q��p�$"��"¢�g��8=��td��m�,�E��{%�>̉�_���Q4�}��c�Ya������'.\���q����z8�:���.�\^74-+���0JJ[�%)��o\­����������SȮ���
�����7B37�ɃP�ma��e�U���cj2�5GM&�#N�uG���[@�k���v>ol�h�&݈����wQ̑����W9C�-��$�+u���gh{�V�m��U��2���O�y��	Mٿ�������e{IőΤ�u&H�N�9�A�	~J+NM���'P&��?dpi�:w�E,��D�q�����
�͇��'�G�>%=()��k��ޔ�0��L��_Fz|�l�T��]8��(�]��������)̟�M,jH�A��G�o��h��fi�i,.�ɼ�L�$m����vD���1�q]��L�'�t�4Z�_3��������"r{{�)2��4mN��@pF'
��_��?���&"t��ѪU5A���u5���1�w�mx��o��K���\���9kI�f3F�r���ONa��4g�ZRD��[&+�[0�AN�.͔�.�F��{Hs��o0�~(��H����0*�>���|��.���ؾqŭuՀ�t���HL.�����I/B��u�o^�;�h��������bVlP��A_#a�3Y��}l�Jd'�2ͦ�� ���dޗ�����<-2a�`2F���{�ϭ��a��SnR�}h5�(���2.����ha;W���qcs��ʵ����<�n�V[���>^�������u�䗙ڛ7~h����n�3��xH�.Z�<��)
�I��<X�HF�)�wE�A��i�bL���=�G��x�}�dq@=8���Twn�߬�Q�K�ǱG ����HMLȑ��/������z��Y�3-hǵx==��5�4t��� �cn]��ͭ-4:-����B�ﰱj�������W�������'sNϞ9�p(�H�uȏ#�I;_ov�7x����_������ҡ��&PG�Zˤ�6r[������nǓ_}7�^1`2ׅeֺ�u�'c"af�r�����hH]��!�O���?J,�I�6�]>�^���4��U��fp����xl�D��������)��G�UtA���fp��;������27��Oz�Fi^t\R�q����]Oo���><��F/W<ȡ��mlt)�����Lcbv�XLU�X�����&܌����Ӛ<QS�$�F�\�X$0�%�V>�S�e^xR�Hk�K����:$6�2���u璠��V���J&��PE`ٰacZ@�n��-��cAd%��#�#ҧ~�ׂ�u�| �d��E>,r�1ߋjWw�j��؟�ߎtT�I���n�Hr4�#'N��֞
�@,���F�76wtȱ��C����(UZ���6B�Qџj��(��6P���k$���<&g�	�P>8@io��mT*Eӄ1/h4���",�vU:-�!��q��D�[G��G�TB�;@&�R* 
�ՈS�R�"Q>�<Y�8-ce���,�#Ѱk$3@���c�\:BF��P�b�C����J.i��)���i҆4��gF�6�S��I��Є�ߗ�	�7�l����H�.Ss�����B�x�������v'_��H#����,���vw�H�������lu��|7�&�$���(�m��}Na}����Y̭��N	1�W�8ؾ����r�0@x~��e��8�u�S��I�8[k����E���шA� �x�RQnk��'*FS���1Ԝ��.6�n�V�h�H�-�b��!5��zK׎�9�@2������AN��Lн/�+��,u����&�N��q�u��m?q���'��%�����c�S�ojA�X�)�M5�1OKtWK'�fM���\��׆3Yi��WP�6��d����è��6����>>��/�O���������gx��E���1�TЅ'�1�65�%>�4n��[_C���:)�~��:t�DZF}�>�̌k!��,�#����2�>K�9�k:Z����Ԅ�r�uk�PT����.���,:�<�0|�.�ƛ�����
�M����wƱ1�k���ܒ��bmk�[��.��LЍͺ���f��GV��c�]A��݃�&h���EsO逥�)ul��:c����k�5#Xe���i쉤��'Rfs[ӫLv�o�h�eg���=?�'�_���#H�/��!�"�v�y�<vv_A�Q��0��4R3KX8|�0��6�A����ҋ葾��8����2bt�*7j�x�kq:��t�yi#� ^��=�w�Av�#GAւ|^H�"XL�#�=� 冃��~_��籵��}��333����qFCY�D�R�d���/5�	� ����>�wv�G�K/��D*�&́��E�(rZ?Ҙ1��sH�e��O��
�WAi����"���p�쎃P(�\�Z���AN�*���v�p@ö�49�/(m��h�qW1t��8v�~���>��_Ň��#X9zZZt�0���\{��mT�1�7������ѣ�g�*��*۷�v�<
;��lF[:���FG�B}*�vO����7�'��Ԫ%l�� F��L����bG�+%^���=<��_��~��3�����"^���+��]Q��]��s\���}y��B��45?�G��>�E�]}� VKEK��h��j`|,��o?�/<����c�4 (�6,PEF�3�@Xo��ju�'k-Q��h���%��&6��/�k�1��P�����PE{�ņb�d'He���aY#���T ����.�{��s�ev6�1H� =��e�A��#��6_~�[kڇ��s�\=���$|vH{7�E�SǠY��h?�}ߍl��?�)\�t�h�dL5D�B��Gq&�x޼���W,�4q�N��C<����ǐ���&ͫ�v6��R��}�6��u�bv�>�7�/�q�Ce�p���Z�J�z'N��t6��|��&�U9�
�65$�7i�,�S�KH�G�\Kt]��(�����{�~��0�P4�p�~�tFwJ��R�XVzӧ�&fP��Qg�Kv��;�p�Ex:��M�u���a��	D	�J�*{{���[U��-xC��f��:��6�~+�#�������?�$�al�oagoW�'R[Y�gRi����`kk�-�W�	f��n�)�����ưD��x��\�y�s���!Mp?���c���ԍt� תa���K�b<��޻����ի���u�%(��K�[�6��Q`.-��Q-�A�Ք&2��t@]�{p�
��ħ���'����I�e3��٨ym̞�Sa��+9�d2�2�$�3@����Pz"�̾�M��{�&j�A�!�#M���rG:;O�_Mg�O>$��&/�w*g���LqSi죳��v>g�ѱ��s��F0J��J���o�i�E{��aD�g�L�� @d��0T��6��8x� ���<'K�d:�z�dtI>?Z��qg�����<�}�)�X�F|�f�p�]w"	KI��F���'�HH�.�,�x��v�����j����mN8)"u��<Z�l��3S=-��h�dݬ��5U�P�4��9CuA!W�cr��c�8v�,�ol��rJ� 3=���4�_��b�S� ��~��c������ �������/'����:��ٳ���)L�-!39g�8!���6�9��r���sf��6�����ǒ�Þ�=@��_��ىq�q�V��9�Z����8����nN,�CR0Z�.����O~�����G�n{���瞻\8�b��ga}}CfC�(�kB�f���O����.i���H���i&�=�f���~6A��σ�X<h�@�(u"��ފ.X������Yz9M0Im���,����ǲ�~k�H��Y̭�V��k똚��o<��e�o��/alj�𨌝Ы�]�G��U4w��E���.!��Ctl���Bu��n���E�YG��"�Frfٹ�4�4� ��O�n�N#I?�S?��׫ ���FR#��С�h;B�f ��P)����!\�pAFB�ׯcne�~�/`ieE�D��ɴ���Z���J�^��,��������t4�ߡ�釆�M��)̱;u⨬����/�)`	�1�5��xf%�W�2I}�e�9�>����l�U�����L@6�e��^/��f��<*M�G�q��Yl�l���?�}����=��#����!4"�)9
v6��y��-��?�x�Dv�(F���k�qP,�߬a��Et7�+��!61��#ǵgR/Xn���E�Oj�V�G����9�vK���m�
5�Sq���Q,v�h�7+��/��3�7�q}M��������Dvl�j]1&t54�>.^���ve�vr9�	4�]|���[�f��7Ѩ3�t6�+�Eû��Y��|���N��u��6�v��g����e?קӪ)<���&#|],֥kP�ؓ�/��d����v�Z>��Tc�3X�������$f����i<��y����LE��1�}����l����@�D/|�6�Ϝơ�΢����h˷.]D��%`?O8"��ɣ�,��-�T�y3�4�y�[U<x�����}���g����ŗ^V|�=wދj��:��ڽ�z���gO��~��簻�+��I ���5��vw�����Q�k���ޒ�L&���{AEQi�*6�XPP�!�"JU���b�H��P�C ����:��ɔ���p��=������zY˥x82���_e��6�Y6QZV�ݻw#��,��hT�)W����,X�P��	6��r�`�Y�f��(=��w�_~��+?��]��anA9 ��#�8�M�L,���(���[<�,)AfN�Ⱥ�J�`�����>�hnq"//�=@Y#S|�΄ԴL�bZ��7�W߾��p.��r�����n�Л�Ga�3���M�XB�4F=�H�뀔�,y�s�ֺ��!Ĝ��6�9�R�YY�.s�l@H$�z��`��q��1|� <2�i�:���~A�ݎG"f��rd+�r�Q]Y�gΣ��C4��j/fbj2)�c��G�555"�KIK�8��+d;is$�y�q��o�����    IDATT�5�i@w���҆J� i)q�p�<~��AGY�#����h�h���ɑM���_�6�]6��DZyVxa���p���#�7���A(Q���E8�4.��ꍈ��`LN�!)Ud�*��0�zX��WA��T���T�������t���d��5�Dk�/�ԡ64(V�(��-���
B�h�V#�j���� �j��Gg�k�.�;d �mێ���e�N�@�#��������gl�N'�CR���6��K�%�(�В�bɽ�ݧ?n��VX���2��L�r&�<�6m�*�(��H�'V%����3x :dg��/?�1)�
`�V�(t���
�3!-7)ɩ�U�H.�`�l�%I��I�����xmz�Q����Z�j�zG&�{D̑7ӕ����A�*�~�����CX��n~����XD��t��Y/�s��M)#�h�R�>�(��j�b��!����o�����$\~7V�}_��j��q��a�ۧ'jj�ū��ky%��V�[�Id�EB:��A�ݷO+W]u��=�����Z��g`�)pz����o�	�JO@ۊ^KkYA����#�R���l\1�2��g��ʕf��n�N��l�8,ߠ�(V�={#��:���C���
�q�׾��ܒ�v���Pd?E������S��{0�{�[m�;��F���RY&��JY3�`@�A��!x%cnT���#�`��K͠�� 7�*���<��H	~�d�K{��h9q��[(K�>)��6%���N���&��k�R_%��&ފ��$�fH�g1��j�Gs]Z�t1�;,f|���R��H��r#�7j%�����ɸ���Q�����Z�FQwl����iij`�)��"����o�����"��D"�ҿn�8�Y"a�*Xб��9�pm��Ö�?��ۙҋؼm�l	��bԖ7�M5����J_�;�]�M:	}��B�͠xA��F��y_`UI�k���R|��i�ҳ7Η��� >%�9yH��ĉ�g�l�ä7!��EK���ٍ痾���,�\��6䃮�D�R��/*�5��qpd�!#��L)Q�47���L"'��G4Z��س����6�^��T�I���
FUw�qF_s%N���Fh5��0����E����l�
�U8y�,֯[���:��'9pÄ	9�*�&�� &�����9e��ܰX�������?a˶�J�I.��B�嶑/7U��p[	)1!j�T��^9�کol�Ϝ��d�)`NYyp��)}z\2��5"�,�i(.���%{Fr��DU]Ν-AZJ�-^��O�}��\�61�t�B����ᯮ�Zm�Fm�-59]�Ü�o$ oK��z��U���(�'6���d��BC�z���B��:vcذ~x|���}ן8{�o1���ޥ�8�	&Q�BjZ�HV�^>E���#���~�����hp8R�X�G��!!1Q&�D�g�uD���`�&������Z�G�H�I�C%z��<l�٠Ŏ�[4�į2��@ERm��$��_;7���٬��"��,΋���"[d~�6�z�L�m2'��[���4"	�Xl�ң��y�a\��[�a�>����`w��j����ł����PV煳���l�d�Gv�����*�Z_�6?sV�HȤ�"6B��
�~�֠��;jfN���z�ُ!�@C�[|0����/��+�SU6OM��oh���"EC�Y<M��e����r�$6w^�H2�j��k�Q�P��;z��i�g�7W���y��A�(%��=+Ð��{�N����;�f'�3����t��3ߍ��nc�p����Me����Jy٨S&ċX��*�H�9<h���gBrNJa�gbr�:aڴǰ�H!���1Rr;�	�YkIj0�
wu9��!�u:RO�2�ܹ��x���2n���SQ.g��>�$���C�i>�����7�ô����<���Gq�]w���B:pj�Y�y�٫r����_��CcCZ���Q# �h��u�L��U55
ٷ-*�n�mw��x!�|�-Lf+�N�&݂������P+y�<��Q�g9��+��䐳���0�rf�&��[n���$Z-1%�x+�F3\7�ϝ�Ց�${".�J�Jk���sy�ny^r�sD�Mv��ss�3����{�ޘ��l|��/�Z�)2;vG�>^���٢�0���S_���'j�G��F�Y)]�#�CG�>y�k��؅��3𕗊���8�,^Ә� ����{D!���O�s�\�:yn�p#F���^\���"��&�K�N��։�).>��w�qqv$�d�P���,>gٺ�V���1�]��b��ј>��?��|�*<����0��;��K�� ���T�H�!�}ZVT�1����kF^��G����"�ʤ���3���lFZf�]Y+qh�p$��Fe�n��I�0���BU��K9��@����%�9>-Z�m�[�o�֑uB"B"�!��@_��h�8Ua}��,>��3'�&'���(��O��6T����Pu�<J��*�Y�FOz)�bn2Q6�Z8v�y�u�B>6�>�}����޻�l�kعu�4�6�]:w�̙��`���$�����0ex�4�A����y�n:x׎���<������3n�x3�z�~����$M�@W�.�"0ƛ��誯�.؊~C�c~.>�h�Ux�	Ѵ�H�W3(�@$�6�	)�HMM�wG���s0�6�͇¯�-�6�B��3�F���*��H��%K��=��!�
':�X H�%e��2�8�\R�Vg�d#:��biq�f#3�3�Rd���PU]	5�J�a��$F!�nCP�"P��зc������^|z~|&�Il��cTq��"1���S��u#Gb��?E}»0��fY�p�U�|hv5cА�{�(�������f��[��Ԃ��zy��)�0�V�Z��쫯����h6�����'�G�Y��n:t(~��+�.^�����A��9p_�ш`k�)�321x�er���b�Ni�ڹ=\K[ҟ۞�-ɤ��n��H���B������1 Y=���6��0*�h��7�Q�+�)�ە��	Qp*�]�c0�ʬ7�`�5��d��/�1wjYe��}�k��B��o$޻��!	�|���T����������㭰��!��=1A�A����p79tyd-����o�=5UB>�a�|�
��A`K����c�d��r���j�N�z�E>���0�v��
O��؄�lc����S�ΰ'�L ���oCCM�|�l8��G����FI\�[�+�3��R�)]8*�o�	kb��4�IX�L\�k4n����`]]��,>٬�`����$)�_?Q�*���w�1R#99Mi���L�͗i����RJ3�/�`��%͠%9K2���WG�����TuQr�"��2�����|$2C�R�� �Mj[_^
�A/ς=#	I�s�*�I�r���\b޼�����i�LA����GM]5����i"�@o��D�CBOiNff�`䃭��c�ijj�\J�K�/��kk������<\,+Gmm2�;��Y����|�ŗ"��#��x�@j�ZIn��"��d�bsKN�5��0�/���ϼ����'t~�l.���?D�-�AR�4��᳙��/���2��&Q�ֽ*j�PXxIv^Z�o+�zn	l�YP���Z��*��^�x*�x�X��LeV���6J���{�P]Q�>��Cm6��H��WF��Bϖ��$!��o��Gy�?3�����Q������Eީ�Z�ױ�x&���y�q� ��Hr�bJ�Prb<<--�{��a��f$#7׍���J���_C�_��&Oƺ�QXxT0~����QBCӇ�E�Fp��AHI�cˏ��{�_I=ʶ�[r������9Q2�ψ�ܥ�a�l�)���O%GOW�[���z�$yZ��)�u��c2�[����Ś��H�\0���l_N�Q�8=�m�@��R��?'��yH��+1)))�D#p�W���q�/�
iQ��i�5��[�ѫ�5���ǿ�O<rn������r�u��Xo�v��Ā�e�Tx�$jkj�P�!/8ʝv����cj��Q|�l�V����-ı�'1k�l	����y�d�K8|��2镖�-�q�:B��ѣѣk|�~܍5BT%��51E�hd�f�!++F�U��hq5��`5ǡ��J��, X��26-2`���F�����t����}Z��o�=��.�[?ErN��X��`X2�����.T���J[<2�����ޥ��2���+~��&'�N"�POS�ĳ�H���M#1<k�ii�-�ޅ�OO�}�Δ&a���٧�aɒ%r>������Fa¤�8[|u�5rJq��t�!���Җ���۶nŉ���I�&a��98v��?0C��&L��{�a޼y8q��lT$��3QH�U��]`Q<x�0�ffbӦM�z]r>r3�a7�|?���pLgAzF���̌���bq�H�3��EI���J���� �:���f�'ؐ����s�E�n�%�b�{�>��u��s��x湧�i�X��'���1�:�DBTwD�`�ä�����e�PW\$�~M�
FG�{�I��E�GM,���
��(����fC��&�U�	�V��	7f��n$F����}��g��(��+��9������N�ME
� �D7�O�;�f�W���Y|���|�zj�l����[����c�ڧ�<;%�UX�p��΢g��"Ǣ�E�&��H��¨Q����c8v�4j��YxCǋNo���d�~����{�Y�}>�[ΆD��		�kb�Z@��$-Ca�@ҧōT3cZ=��I�c�=	��$D��Ꮩ�2$#ܪ�^���^R�n�1��$��ԡ�2��ry�[�m��S�ܽ��W��h�(G��*���=��� ������������Pq3��/��wގ-[���� ^�ݎ���b֬'QRZ���Erj�(@a̨�y� ���׏GQ�|��'p{}�ݧ/���R6z�X�{�4�_��~����4l�(��`b�z[��z�*\~�������u�|��NnӸݔ\.c���#95iiiR�^>_je�:��v��"��G�<�ŀ�U*9�qҚ��Z��OBf׾�ť�I7�4���H�U4�Dmɪ2�ZX�mhhl���8Ut�]q-:��Zw���jn�`�j��1&[J�*QYY�V���;��o��_��܇Bv�|t��5�up{\��=萟�������K˖c߯��S�n����0���e�|^44�ㆉ���c����r|���hht�؉�hn	�C�np��b������~�x�T�h�{Ρ����z�mڜ5�ԫ��}�����y� 2����?����HV����z���GJ2�LQ�Db��lY+}���^��f��wTb�T�dn������A��3�������]&�ڛ�^�d�� 25�$a���F Y����M�(͠�a��_�A/��fP�Q���`w) �[2�9A�l&bN��D1X�Ā���K��
��7�5�)n^6$o�dR��]�ҩ!�H�p C�Ǣ��g�~��6�ÕW�@Jj
��y �/@iC�^}�����'�� Z����f���-*yj��������e!��B�߿'��z>��?�Cq��p��#Z��eѼ�V��_
<�.I��̨�p]�������V��i�����&�*?��&�h���<�?_6,|�tH$�Z��z��������'"5;W̲EgJQS����EK^��s��#.��P.��"N�IF���5����6M�+H�xzZ2��\7I�]YV��Q>#��$� ��D)'Ga�g0�7^CJ��ǎB�}��̇���a�����Ե��L����]n�j4&�zq����cl�釨��ıÇ���b����C�N���u8x� �i�3�y�-.��5�K!����U6��VC1�̇�Bf���'�6�|���h�n����EYY�H�x��b�g̩��d���_�D�̦1�>5#��Ò����t���u8~�	�qX�x��0f!�i9И��ȋCϩ��<5��׌(n�I���E�YfZ�i���"��Z���+����	p�BoKP&�~7��1�f��}��W(��=�*+���U�8	����[������:���B6k�T��p�7H@���M�q��y�٬�e�-x�Y���C�뮻��چ>C�a��9X�r����32P�*Ax���!�Á� �j��͛D�+#9B��JC���'����476Bo2��]|�"M��Y��C]He,���S�����A���}�˥Z���`Nǎb��3���ؼu�4��]��K�/~��
�����uU���3�E������LP��W�ek�XZ�Hu�����FCe0K'�6"�S0��[��}�1f�x�f�[�?mۃW^yQUii�r�]���+�X� ��%�(^D,���r˹��xQб@~�d�"	OKM���c0g�L����>}�l��]}�>�,^����K�QQ+S}Ѓ-�����q�Щc>֭~��z�E�3����u��l�Ԥh���G��Ry��2L঒B���d9{=>�,���57�����^�ݻ"�c.��
�ʑ���xp����I�X���Ω�Jv���Af,�0��\�Xx��Ҕ���Æ�ńAW_	/�i���N��8!a��XRSh�!%��	�=��_w��S���'q��!�^�<�;�m۶ɰ���M7܈���'O���3J/�y��E��%�LCC���лW/8p _}����:w�����֮��h�=��'b�ܹ8s�HA�S�Ay<%�"yo��h�~�H�����}'���^�p�x]R�M��:������=F
vsu-�22��(/-�����W��Acc=��I�ڬ�PR"r\�1�	��])@���Zt����Ö���?BN���j,�i� M�CA�8��F�WL$�a��U��	.V �{���A'9h>�<.�=vX�\��iBz>q��(�6h��k�ѱ�7�x1׭[W��r�������s���/{wᥥK������4xa��D�G�_Ey):���U�%�g�W��Y�q��HNKź�b�ϻ�ץ���2N�<��/.����fP�R�+�QT�"J��W^��'p��a�G&A�ʽIi��9��� ��,�2a02:��>R�	�����D$��hv���>��'
���*�!cM��MR��Oo�>)��4D��s��� ��(5"s�ڢ��~�4�9�7�L9݈����Cع{/:��˯��H�miFV�W3�B=n�m:Qh��v�*��rss���p5T�ɇD�=�]6L�dXp�a������	o�/���K˗c���p�����ښ:�U�U��?��/.Y*�wW��_~�M6k׌-���6o��C1��G��W_��>��/�Ħ�즜�>j�_�CC@FJ>��#�	���E��[z��E�U�5�֨
I���^F+y��?����z�u����ǃ%����("rő�6�Y]��-.���ZRF�R�Ά�m��A]��T���Ū|��f\q�5�?�7~?|̈́Z�̉�� 7�uFec��>%�z��2R0��	�p�,�/X��σ��!)%I�ܴ|�:��ۧ��ً/�_���7ߊܜ|��MZ=�������c;~�z3���lX�� O+���(�F`�.*����{�&[DM`�B6���u��o{௫@�.1�_o���w\(>�؄��T�U�Z�L5U[׀G"�LT|\F��a��Fh�+� g$�S���K���r3�&�?6�l�m�*͠����)�������[��M3��DmPqQ���)9��(��R���C��һ�D��sM���d��H�C��~�l�|�u��f'�1�`Ku��A|�C�1�/|->��}Ы���U>Y�˒�A�^~�ex���X��MlߺO�~R�n��[��3gEZ4j�8Y��?w����M    IDAT��49a�|�_��=���dt��eʰk�n4;9�jó����Q�bÆ���7e���G��)i�+��SW��f�4�X�JU҇���8Y��Ht8��J�/sz'���(b�*�N�p�6G��`pC-Yn4(��0h�pT�5��d0�I�Y���	�K�QS�$�\��-^�چf�_�[�`������U�!��щ�*ʒ|"��!e�ې��(Ek(䗢��r���~NZujD�O�M� ����[M���;ra�x�x�=N�O��|��:-F]{|�A\,�(~�;E�ܦ�8�ʣ(�`֧w�W^Ěw߅�d@�^=���J,Č3����aOM�����B)V������Bȍ��%%��'��'>h�?C233�!�WW_�f�S69<JKKE�ȉ�aY��a�X���I�5�A�j�ڭҲ�q��Yđ�����}E&z��i�\�P������55jK�\B�cQDb��`�4��Mեh,+B4�G��*��D�ٝ;V+�$�<2��+/����L����]hjt"��Bnōwފ���Ń<�ӧ��iXa��?���)99���S2�X��Zٲ�a��	��H�j�C����|Cǋ�^�!cǏ�M�n��]{�쥗��r�5�0m�4���R�8��Ę�X�(��r��OY�F�A�"�l¶͛e�!�6�L� K@����nCZV��)����3��_P���rٶ�]bQ��E6FIII�k�]e3H�Δ �{�?�F��i���V������EF.�bFh���R@1sͨS���8�s1�����թ�ӥ@��Y;ʥ}�?�x��Zdw錬�l�z�>?'�ٙp��`������q�-����
w�� Ν.AUE9Z�܆�c֓�����U＃�3g���)�1t�̜$UJL�S�N���>�����{͡����M()� ��n�]�܃�/��#�-穜�J(b��('x��ܻ���Q�!k�]�`KLFF=@��8$�R�Xm�e"�%=����-�`�_S�b�9LKEs�K2[m�9#�Ї�APF�ܫ�=p��(0�k2�R����O�C�x����Q�Z��K�
�I�[�*?-m��ah��ѯ?t�6�75�o�������kѹK�V֣��"*K/�s��<ir�sd��G��?~���gB�[o���wf=��N��7R����ګG�ч���V���>�I>i��V��|ޭ���[p���x~�|����+hjh�!#��L��{v����g`�����3ϡ��L<����L�W(�B`5�3@?ٷ�~-w-���kΦz[^�D/1�tL9Y��CSm�v⭨%�Ű�(����-E=����Li�����c*\v�hL&���"�k�9n�yo��!r:�F�ւH��/�_0��:D�M���NFJ�A�P���~���������]���O��xa���\Y�d�S���d����T7{d��x����W�\<��\Q��mVF0΁0!*�y�l��=<7�]=B�?��^�q��9iϜ:%Y�o��
��xn�B9��]JJM��1ce�����J\��+����x�7E� ���5K�AR!4�%%b� ���cǤUs0�W(�<�<��F�X���o��2k���h�o����_��E�����B�kT�p�Έ
h�"�5$����0�&�CF�� �ㄒJm7�m^�w�xt�J��_�!;%	�o�x��<5�q��l�8�'���;o��Jp��$&[Q�Ќ�g.@c�5������K�C�[���1�w_ęHk`4h0hP|��[��z��xF���+��*B��8��/�5z���[()+�{k?���B�k�z7���y^@v^�Ϝ�-;~���� �C���~ᦕjY�o�a��X���$��y�^�ҔA4�%�($�K���f&(���&� ߛK�,�/e�^R�\*ϥ�b�BA�{3��zR���j���@�hEf��@|
�m�h�Pk�E�V���D�Y��׏�1Ҍ�لn]:�*��;a2X0q�|��8�<
�-^H�C��@�i8ZT���bԺZ�^�Ƈ��{&O@]i9V���Լ�Bn^RvX�F��%�^bb^}c%���+n�|;:w�"�����%"7߹s�]?��w��n^]�B��-	�e�������ٰ�������2��=���� �~N< gu:dg`P�^�e�^T��ʰD��$k�M�¬u�4�\��o��o�����p3HևH5/m�\��f��&�*e�F�-?�v�'e�P#�������fB��f��d��l�������3H��P�X0�B�R<Tj�˱Y$�Q	�-�Ak���&<.	5�o�Y��!HMO��|scJ�\�������ҽ�^Ά�+)�����+��������G�1e����y�| �YY1�j��|�ŗPgKC0/)^"��p������&��ƍQ�PS�w��R�����g�NX��0uڃ�н��k��Ѿ!�X9�����;3�U$84��?%"�� }?[p�\�ƚ:�L�<���S�aNͿ�K���$QVc4�1d��ntJ3�M^bZ&�:�܅��kl��h���EKPW׌^X�5j�Y��q��5#¢�B��������I�B>���1�k���-��W3����#�d��
!^�G��}�*w��iTT��W�z��i�e�D���W����C��r�Gy�x����������.���4p�I)D��v��O>�|^}�e�<�����MM�X��E��$������q��o�|S�s2�Q��#�*]6�bޥt�S:����w�EnZZ�LG�5`�is�SANUY p�ί�j�	����9W�������ѳO��)<�=Y���n�Q�Ԍ3E��H�Lt��f�~fG��u#j�S��J�>��ͤ�&�FC�Yx����݂8����_�4t0�>�x���毿F���o�����Ec8��7���3�� ����X��,X�{���~����щ��$�~b�4^���v���|�x�R�RE���O��C�30u�=x{�{"9KKOG�}ѱsG|�ͷ(=_(�+��7M���_�O
��db%Њ��*>i�������-رe�x2��_I`�l�q�-�Ѷ6)��Ք���a�67�d�ο(%�Ŧ�>]Jeܔ�ku���}�@m6�{�����I��`z���㏻�v�7��醨��;��0�9�:�x��&�U�y9+�m���a������~��3M�N���x):����'Y.+��G�a�ƏP��(R��c����݁��-��Sg�!'��IMA$���ۂ�}\ 1��?/0�1����B��]:a��IqN)�M7ހI7߂]{���?�Ĝ�5�/o�u2222�z�{�ۿ?�L���o��¢�JP��?��A�&p�٦V�ڱ�ѩc�_�.�F��5Щcht6��KǸ533����gmCDFyy����m	���1�ǉo�W<=�v�����ݖ9���t0 utF3��v$'e�Gg�C����`M�FLK{�I6�u�����T 9ހ��z��t8��Qt��FL�c�gc�͓0����[�u��fe��ɓѵs��N#�jBNn*�yg>,���k�¬������٠SREɳ�
��O�,��u/�ϝ�}{~���B�x$���|2�Xv;w��ˋ�����V���hVUVɹ�t�R���㮩�b���|�]xi�˨(/��l��?��H�^�e�G��F���Id���~#dUzM�=焹��FdP�83Z�A)�G{���j�v����O�G>��q�F�D�(�R�u�"�6�p���].��Ff���h1~���^�!����hG(��B#TQ��FJ*�%'�L������o?Ƶ#.�0�����c���%�q�|�|�ƶ.��Sn�Q��g���f����1n�(t*�ƛo��!d���l�`���Fc��_㕅�0v�8\{�u�u6�����J\B PuU^Y����x�(/�@FV,�VL�8=�t�K����]�0w��|A��z��8de!�o=J����@�o�р���Ϝ�y�c�bT�/�܆�A�RqAEU����}-K�`+a2(j��PPJcz����m�Z=�,����Poc3�Kz6T1b��ѧ+SA�sI`6i���"���G�˟���];c�����u(+��K���/��?��F_�܉s�+p��)�Ǥ����:�}��s��&X-mxy�K��5 �d�ı㑗�!v��)Ͼ}{�˯>����'ބ1c�%��uF����u;�j�[�.N�*�{�ˠh�C����x��`M����={�c�$���Dɺ!�_��? ��IH�]HjOr`����r��Ʈ�03�r.��knv#�F?u�</T�ܻ$e#�d�*�cJ����l�!<(4v�a��&��x�lC�x�� �5�Ra	Q��M[j��&_7Me��㵸��a3�zl۲gϜǬ93��=ؼ�G���7��޹�RG���(�J/���B�=Q� >r.���/� 2��Ç##-E6��c L-�����p^y�M���f\7j�w�! �ԔT�ո[��s�O�~�XL�~v���6n����� �#�I�2�y�5�k�a�V�79Ee${*��RzPv���j��d`���T(>wZ�-��'АJE�S��3��CIGj**�p��I�5���2Q����R3�R'aB����?6���S�k3������`�%f�D�=��\��x������B'�fPȍ�f�b0�F��6�Y_��	��z�{̬d45��v���#8�$&��N<e\]�������������X��B|��&�z��_Ʋ�dd�`���0�X�t)k�1�+�s8����ƀE �6�?u���|�jj���جA��]e�y��T��ˋ����7V�PhY�+�u���Hc�p �p m欑���5�&�C�)c�e��2.�X�<�R#@��V'[N歱���%aí\77���M"՚�`��<'��%hts�JyT�.z�.,|�eX�Ӡ��I�)iW�66�4�FaT�a�Zt�PUrQ��Vr:�b��g������r��7���/�� R�͎!�.�5׎AiY%���5j\�bzr��HOMì�Gǜ<d'����q�/�``�^���4�^�
���-�r�h��Q��IdEy%�m�&PJ��|��t)ХK��лu�s�Oc����Z���<u�[��(�z|Q��H��� K0im���{��?���e��C��-�=?�\��--���!���o|����i]MC���N�G�~}������)!	��4�t��J�K��HT�A_?5q��P�mhS�F�BD�h��b,z5�D��h�-���"�5H�3b�KK�u�P���'�u@fj>Z��f&�4Q�ܶ6��m�O;�J��!0{�,�P�q� �**���I{j5��Ai�fL����T�3��xg1K�p��&��݋�7߂��ބ7����I)�"릟��b5>�����&L����|�Yi���Q�?�2X�%ŉ���}�HS�o������A��H�4���%hW�Aue�|�ք��xYsj��[]�u����:��B���C�J���:,v�C�bz��l�ڍ�!3�b*�4��P����Ȥ�*ޠ�!D}��:{�ϡ /��&���
�v&�#�ٰf#:w���c���HJI�����罿���?��HA�>�1f�h�^�.j��a��Pq�"rSЇZ�1c����O�ǲe/��_�aĈ�лO/��v�T��~�]
�f�#���&݊ݿ���Uhmkþ={�{���Ge��#�O��'ga�p��E�Ӫ(#��gc�c�gk�hï�����p���-��"{#���{6�""��x}U��.nt�j�*qx�d~F�5pZ��ktF%BC������A���$T4�m6X�dK�O����`����G������qn5*��^DU>8,j��^���V��`._�_~�_zM<��_Z�����{0x��HKMǩ8���<�'.x�7o�߇�����7�\��G+C�H�9Y��ܸ̒�L�i"��y<��'�P9`ڿ?��݋`��/��؈�?�\6��E�56��9O!!93~W\u5�w�^�.�����b���nQ�H�	�9��W�n���}��H�HG��sAΆ:)b�N���Z�,�����U#�A�"����(��As3I��ٞ _K}]��m����it;����g.��?����7 �� hL�V#���F��e��Qw
��5}
��p��p5��z8�X��O��������ֺM���t��E�.7b(2����������)�j"a��z

r��{���X'5�V�ð�CP��-��#�_�=?o������1v�8�:2����6`��mp64b��Ո�7���H��MR�N�1f�X$���5��ȑ�xl��pzX�z5��Y��Gi��Y�1���N�ˆ�CY�9;��(������@ _0 ��d�(vd�T������!��X�z^i�����x�h�"��g��������0��A��� ��6A�L�QB,ﭦ�@�4��?p�-ذjzw)������?�o��ǒ�ᗃ���U3��{ϝp6zq��qV��i����hl���A���߉xs�<5�@���q��#d�B2����r��Ͽ�k׭ňkF�+F��l����"r������DV��JlG_|�5��BEM�O��N=�aͺ��!�f<��܌�;v"�F_�PI�W�C�����bQ���r�����h�#����߂R�r�&������'�H3HY"�}A�h�cwĚ�����ʏ�	�1Z��Q��
����,��=ڄL8[c���-�3�	a���4rl���K�|��f|��ר�����<�wl�ǟ�o��p�R]�S'KнT4�cӎ�q��B�}��?���?y�?��(uF�)�'mGAw3R�q2t
z��f��o�E�N��5e����Ɔz<x�4L�z;:�-�w���E�ۏҺf�%&K�v��7�j壏>A����)K,�Qu�,�����ƕÆ���у������:<��6�l��Wܖ�d�c��!bKa3�R���LT�p�����Ae3��(=�����f������}���Rs��?�D�|C�3������x�n~.���9�*2�K�ANx�
��T�ۃ����a_.H�I;|��tN2Y�����4��#�Z�mi@�� �/[���m7��}C��Z�ʳE���To�Ν���0��Px�X��9�f ���a維������1��z���p8�z�12�_�|9\-.L�t�H��~e����_��w�% �~��B8YR�z=���?���kpݘ�����G�|,� |D��-I�V�Շ��	!�X �8�Њ��!�-��&�>��"/w ���dz�b���>�j��������L\���7pj�p���Y�H�-5�55h�t��~�D,���^,Y�l�Л��HC�."�HN�55LT�^D���������r��κ�8z� ���t��>� V�X��GN��)S��VV^�s%�8Sz�43�'&M������pX�"*+:m(
�F�a�b�}�`ժ��s�O�1�!�~Ӕ��d#JI��}�����������[�����D^�<̘>��?6Ǭ��f�o��_>��f�K����x}2��4Q���Ց��Q�{�{I�q�S&�T�Yx�g~vܢ�����)NY8[��ѥgO����B	L�%#�k4{(�G:��j��y�����s�:2����&#9���V��a$�b�x�*�����/,y�f<��s�x�2�����;o��!Æcǎ�8r���ƻv넇�?��k֠��9���):���t�yVDc��T),��{/�2�q��3���d�ع�砎�a߶�����c������M�<_\��
�|�$���    IDAT<5�!��w��!��뮻����P[[-Rd��%����&�\8D���l�m�.,�+ˮё��f�!R.R\����� ��pX���\pXC@�F#�B��r��Ú�wC�4�*%�Z�!�'#S(�z�o���l�f�;dfw�f��(���G.9�yl���NC�Y�*�@c%Ο8�D��|��/�������e��t�+8��q�f���ϕ�{������~l��3"1.�jƏ�uk����UZx���NJ@�.$��'���w���]�D�}��������	�'���{����?�le� �~ٳ��s�ur!�[��yy��)��P]]���Y��\c�8�� ���XE�o@��%���aFD�
x����ߝ���eiB���d@�=����z�Q����<����� 72�'p�`ye��G�E�t��-H����'�b��",]��y��ֲ�`�FϜmj @,�&m[ O?t?���	ۿ܀��}�	fϙ���W�w���;��׿Сc7\�X)p�	�_�q#/CC]����AD�~}q�]w`��8q��t�C��̔�3��q��aŊ7�{�<��������E�L6l�5�^�E�����5��������7�3��[�c��u��X��[�94���I�+e{!��p{D���g�`$Y���7_��q��,�`n�Z��>2oT��UH��@�-�u��o�;�M-Ͽ��*�
����潼�ZZ�0�����II)8}�,�N����$@Z2��0��eزg?^w=���60�Cb!s}�GCж��d�a����䱿����p��1�o\?v<���7��`�;8p�.2��tð~���R�n}{����X�j�d}�[x���G�Θ;����e�cvf���
�s0~�58z�/̛5ݻ�@��}q�b,V�	�0Q\|A�$֯߈�D+,|gΜ�����Qc0t�0?q����H�/}GO��wVI
�d@ż���1[�EBH#i{�XTU��׽�ᬯW�J�n9|�!�� [xn0�������0�1A"�7[�����ņ���*wA$
��f$&�X!pGg����=��T�Y��5��RJ��7<��� ,���Ft�3����	v�/-Y�����شy3֭Y�=��o�ިd�VM��g�>��^Y���
�ݑ�%���Ŭ½S�@�́[�O�=.5�Q[K�{ �Y�4i���=^}�5�t�Grr
�� qVɻd����3�r�ex���8Yx�v����j�/)������`��Wa��s��Í���/aLL{L��N� �{}R����3E�8]xu�6{�G�l�8�c�	)Ϸݞ,��%�
���
ݜ��Js(�c���#'���)�2z�l4#�"Lv�%N2��#:�
cR6��@(F/)���UaX�H2 ���T���fd�'���r|��װ�����;�c�ox��?~�z7���Cs�?k�+��?�ك��$���sf>���G�شi4�2	�?}��Ο�&B׼�;����_~���< �#���Fe#ŌI��8��r��u�H9~�u �-.T64���E�͎���y�"G��Od�n0[$�w>�J��;w�|5��	�ޣ�r�	��X��3�д�$^#¼s�Y��a�dd��A��L�k�3�������2���'�K�4�*��Z����A�&*8���3���Nz.�s��$�zc�����[�0���g�M��^,s�(������ox��vX#L�
	��ѭ��z��x��7�s7�N�'O�Ę���\�y�QԷ��c�^�44��x�O�y
;~�;�mA�yp�����"�Y���:�<��2�n�~���ԩ�t��&RFY�ɓ�x���������f4�8Q�n�3�=��=�b���X�`Ǝ��\lپMȘB.�J3�Ja�f0�l��ݬ,s�d�خU�����<+�������w�a�&�\�X�ˍe���4D�0$��,�0��0��h����""#5�~�� �,zKLqI��ӤnC�V�;PqTU��f?lq�h:q��a$j"x{�{ؽs+>^�
z��[+W`�{k$S���ȉSX��S���p�0�F�҄��3 +^{�qZ�+�v{�g��+�a���O?�O;��	7��r"�sg	l������/��#=����Hd�R^K�8��	7��5^��o��_���鏣�����	F�Qy��̹Ŧ���H�g�K���X{���}�:{�읐�@�"uֽ�uSW�uq���nPk�ޣ�:ڪmݠ����l����������>}��}�����|�4@��}�}��*��O��P�����a+�/k���y�}wL�ɉ'�ƀ��~�2�����iB3�&�`��M0��0{�1n�TQvl�@Iq�]}5r+�^p���vo���iY��0�T8Ad��m�%�@�!̛@�����z�����o������Ch4��K�q������sf�?������N�0i�f\u�ex����w�����@�4=��x��;G�+W��
9����PV]	�ӡ�����;�fŗ��Kqƙ?�_��6���dBn�D�:� �[��>�'L�6Gu$��9�Ԕ��4,��=�M �'	6ffΘ&z��-*�D�)CSˢ��4��G=��Vd2E��с�ʙ��E��42k�Nă�.cZg�%+�4�������'�#���gj+j& ���l�2��,C�JT:�ѯ�BZږ��,S����օ0�c���r-��E�֛����0����5�t�\wz�B��<������g��'{
k��
�]Λ���>���~��>}:��N|��G8�Cd�Æ���ta�_�\�s��9���2<��kx���`�vQ��]�������'&�N���<�0���kM_]��j�v�v�U>m�t��>x��ź�>��ɁF���
&�ө�r\C�o�&= ��i��Ho��C��0���j����[kbʴ�6���mk���.-Ŝ���DDY��{ 7\w36����>����Ț�<j��Sx~Q�r��ly\}�yh��Aώ.T9�u�7��������_��?��x������fD�>{��m7]��׌��:�;Q�P�#�9�7�̿�V��>��&�(T�}k�N�&�}ɒ{�|�r̛7O���z���.|�|�������"����-[��@F1S.���ǟ�cO8W^u%z�o���BԴT"*WT6�tЖɈ׋�S����j߉�}���vQ���H͕FT�ui�K+��8���j�e���۹m��tk������ƍ��+*Beu�?�p������2,��]5�nZ����)x�y4M���d�F
nd�Y�F[2ID���RS�E��ё��BC�o�������P߄�?�$nY|/�|�����;Mp�S�w�9��ո������o��L;sw��&L�V��z����u�������َ��
�x�|��-��Z��%�t����n���L����@���_�>�d��Gf�1g��b��+�<y
n�ݝؼe�t�4�\��D&���8�p�URT���>�1�ζ�6�_�NA�J��;�Q���<^fH��>5j����>树C�����Y�4�[vN���q	v��t�ta4�@)���8�+ᩪA8C���Y&B�Hs�g�7�Xq�����`����2Q��,�Yn����V���b}U6T�\"��v�*�{��8��y���7�5��oT�V�'@6�i���s����O�W_~�M���՚4�3���O�~|��?�Ǧ�F�[�H�h��9����j�a���S��O:	��"<����c�fr���͂x�����s/�VZ*��%��n��U4�aH8#��L�����(B�Ql޲��aÄK�vt�7�ls�x�&���Z��X$�,G�2o��w��w9���l>�DII������M����F(kA�`5j./S�L���t���r��<y�>_�)�ʫp���������BIY1��38�9tvnä��;2����:�����܄�/8����q��gi�W�X!ݵ)�B��FE�L�;_��}Q�̥�e���$�ث��>��b2a������RS�&t�chtT��g�%��3/�H�③):�Ӑ�"M���_#ܶ�8�|NW���Zqg6� C.��
�6d	cu�,g28m�l���_!������&�搌4��ǚ%Rce,c���f`A��@(gEM�lP3�Y��_��fp,��p����Ƞbi-��u�X�)�i��;�AM!�(�i,��?�f���Q�L!��Vf��e3�};Z�j�/�{o��6�ǁG���x����}��e38<��Ɋ.x�ge�=e�t�t��x�/o�����V�xR�@j%3O>�hdж;���cf�s���oڴI����߈��z����ؼy����p�I'btx��N�''��39�=��s
-�P;����6r
3I�7�~�py�.8N<9͡V��t���T�	6�l.���2�g�]��7�&?��TK8y�^o ?�{?t��wxD\p��b��G���QW]��7ބh(�[n�VG	����P̟!%�0�As�=�MI��9DF��ߒÝ�ߌ��6|���أ�v�o��.��r�M���[M��a�ƛoaG�6e�\q�Uh?�^z�Z�7���[4�"�?�M�#��/���s���DMZ4ef���oV}���J�-h4���cdt~�OM>�}X�vv��L;������/���PA�&	�9�M�)^>��]��D6_�h	N��%�Z���\9�����9gM-b~�1go������i[�ͺÃ�?��7���6oA�l��[�q��"�ͫ,--�u�F6c�u�����a���>�&)���a�5�C�Á��mH�v���/Ǟӛ��G��)��޻�`K[.��R��{���X��j��#�p���?��]���<������	w[z�&~u��]w��Z�bM�x��R��$4��-��ſ�Gu�~�9���������`|s#z{�4��;�>��~*�o)�e���e�r�R`nOJ��t�3&Oj��l������䗦%<��+(.*������M�|Hk��$���ύ��ϑ�@2:0����!j����=�"g��kp�`	ʫ댰s3��C�㝷W��_GU]2
,TI������+�4<��G���bB��C���E��Z���47U����o��߸�fLũ���=��g�y�<�
�g)|�%8�3p���5kq�I����}�:��u�p�`�x���E�&��5I�$�LF�aDʯ�5.�����s���}�����.�m�FF�՗_Lb���5�.���K����������vy��x֞{�#�7_�O?��r���x��=�>o;�v�lm�"�hIi��ј΁t&��"�L���P�)�Z�I�C�"FM[I	~r�AJDeR���;���/����㎇Gy�da���cH�݁T4S:J�9���_��>����a��	��^��y����c�>���[����=�u�p�QG+������3��7_�O���������<\{ݯp͂[�j�7�������g�c��6��Q���8k��x���d@CT�F�v�F�#S�jŞs��������_W�2��k.��f*�Ù���ig��k��߭Y-M.�C���3�k��Msx��p�O��lŖM�y�F�(Cul��{��&�g4Akl�;;K�0u�d��ѹ��100(�Y-4��b��Ͱ:�B��{I���0./f͞�1�M����.^�w>�?�'Ll�&���Y���b����&�T����ￕ���#D_�~�qL�:]r�?��%����!�˖��~v~y�%����{��e~,�a>�O��#�9��Sp������>�ΎNQ�I����_#�W_|�v�n�U�Jꌡa��@��e�.ǖ-mB�{�ad�!\|�||��G�׈{�\���N,^�9f�ʜ�1^���U��?�͒
: ���4�g�zgW�
O��|Lvfr��`s�t&��UC^0�@�DG�C��t
��
�+i�h0�`�`L,�"_)�����o��WOE��0L�]�C��6)Б��;���8��C�յ+��{�5�uUx��AMy%.9�l�vnY����p��������c��MXr��'�pyP^U��]�Ht g�u28২�����>���;d��l����{ｷ��������N�tQ�Y~�+KrX�W}�y�4Ol����nՐs��8���q��ƓO=�7_~��JQn���<��o�:�%CY�#N���e�e2]�ٱ��Bz� y� 0[�(.���F*��l:I��Г&_0\�����5������p���:�|�,ͱ�p��� �������	9���ES��� `ˋ@G�44ԣ��}]�P(��-HeM���жc�L���g�FE��Ca�X�-�utHH�������s�&<��c�0�ݽ�h�҆�� ��#_U�����]��}}r1%%����)�$�ý0�݃��]b���:{O�{�!�a�V�۸	Z&�SN�)��/�	���%H�܇�)}N2l[�-֯3��T&+���G"ExtH1r��E����~k�t؜]}���&�?�%�gTQ�����`@���!ls��<HP3e6��A�¼V�������zW��+M��f�:���mvDp�Y�g�{�A�=D;�m6j�Y��i�k&j�-�N��%7�Q���P�b���v�����o�hg���J�x��W�ҫ��n|�4W��ι�2|�A�i�����8��������ʟ^�#��r��X�e��̩�u�������AmC�6&;yD�2}����z��WѾ�]���n�:y�-�s�v٥���o��6M����i
�g�4.TN����XV��y7'=%z�#C�p�|�='�h�+�ۨ�'�0̰�0Ȭ�4�g�(gȰ���`8���`PF7��$c1m���2,\��h�޶vw�6�n�.
R��hgc.�I��LX�iDc�($c�
z�䷋��Ů�6��<��3x���D�ښ�k���㌳��3N����w�)j��wޥ��I�����:{����P�w8<����g����>�>%'H�~}�bi�؄P�`b�Xy����Ze/��"���e�}���k��C��͛eu~�ͷ`Ӗ�x��G��%pj����c�+�u8�(������ł��¸I�e��tF4#��.�\O<�I��e]RZd����~؜^��8���n�6�i
�-R�<����vT��������k�o����U,W�<7/��ԃ�Q��Gʬ9���nE"�KvW_r6f�T��O>�O��}=#��_��cN�E�]����^|�e$"Q��8|,�8䰃q�����[oǧ＋_^v��6o����'�|���_��Dkva���� ��X�;�#PW;���g�Y��%A̞=|��{�q��F\uՕX��|��w�;�?ފtR�(��p9�Q]]�����]��\{I�1C:���Z�nٺM-��l����I��9z�����h�@wM/�E��ҿ���=��Ն��C�����'�Ｓ�=�j�MF��E��D�B���,r�5΁�AR�s�(�|.,��"��o×��N?I��.�
�{�2���v47���]�'�|Ͻ���y���E���O=W����W����W|��*My6677c�ʕ�a�*&x��0q�������TUW��o���]}��M�Ҋ믽֭����ˎ�9�_y9��n|���c�>:�J�idٱ�n ��8�>vu c|�2"X�XT��r���C���{�hn�����`OO��y���3�hd4����ctx�5u�F"�����v(d�`���Ay�W_� +�]���x5͓`�ya*�10��X�t����Jq���5+��'��s�BKS=^|�)L�8	�8�|��k\3��r9\�x�;�p�u �2�n^|ҭ>�    IDAT�Y��� �>�\yՅ8�܋��m�Z�=}}x��ױa�F�=>�����6a۶�������x՘�S�=Yj`(..����b�׫����~�u�"������#�ğ�1gΛ'��kר �~�N�B�X�0w���Y�7z��L!1\�Iђn�(L	�M(.AMmv�w�ܜ6�#C��d9Єb��d�0C�nU�ƜA��������#lL�>c��W2�A}S�r3�}�S��g0a�LX���V�-v��z���&aɥQ�b����j����;&���a��Y8考��g��ȃ�`WGr�얬�og̜����O�o�Қ
�̊��9���z
&�1A9s4����Oq1�N���s�R��qH�0:;��v:�%J�p�P��LGX�h�礛o.W���q����|�װ��5B�ܽ��Q�f.�p�ό���4��O�r͌<Ai�J��
�x�����#��w?�0���f���O�b�E�|ޠ=�����EM]����8h(-)�p�찢�_����z�;K*�(-C��]�	�>�
�\��(o j���7Ѕ��6��������م��+'Б�!���K�&Mm����PV�E$ÊϾ���nX������~�L.�K/9Wg�������Oz��@�SZQ[S�]}��~�z��V��h����ҵ��CEy�ɰ2z�Uf�O�ك>D��\�D�3x$.��<��x��WPRV��5%=D�=.��C}�������<~/*�+�7 .@ѿ�ձSQb����ن�j�>�1�=f��Hҿ#�l�c6#�����C��� �A���/���Q9���1�*Ϙ�B��ua-��2�`N� ��:�=�C�����[fmYsV��x8����>�rth��81��SƏõW�
�=�p��w��fSF�.sѸ���^�&��P$&*���� <���`5��r*�����h4��Y���de�u�8��cQ5�	o��t����:�{y�%����w�۴Ɉs��@�D� �S^M�xX?Y�d��כA��S3�3Jұfp��`�7m�t͛`u�mi���޿imD�,>�W38F����4Q~��lY",�ѳȚ�H��ȱ�Usrh{�L���������y�z�Ix�������.� ���ǝr�&+����^z��x`�x��g����_�-��`�?`GG��(Muhh�ŲO>1��)���Dw!MB��B��b}�Qj,���Wv��=�ȣ�|�2<���*���kk�pϒ{������T��`|㍸9v��3���zQ][���β�rMF�A#ʔ�m��!�A5,$X:�"���6�Zu{��1k����+���z���a��c2�R()ছ#BS���'X����/�ђπ��v"�
9+��"mKRa�L4�
�~u!6���W,�'���^,��.\q��hl����7LܣS�Ma�P^^��?�T���SNƴ=g��_��&��g���Y���hd+>��O�B�"�i`�Xz�>q����فe˗kB3�K/���S������S� 1���D.3�sX�(�'+���Y�p"����KKf )N�U���	@D����T�P�f7�p׮nW;�V����2Ȧd��fl�ގ�����-����r�*/ío@,��K��S�#��� �l"f�P�7%��f��B:�-�S�=��^,��Vq��8�S��sϢi��Jq���!��e����8��a'�E��M�_�-߯�=w�%��W_;;���$q�!��u�Q�H�$M8�I�θ���/����ٌ�0�����4�����F1��Õޮ^����p�e��;~��+>��c�3��TíV��e3c!�y]��r�p�.vWT�*���vʔ)*H���924���%�iwܗ|��kt�L���ɑÃ�l-Vt��(EeM�zi&���c��?����$X�ȑ�c�@����VS�d�HZ`"�˒ǼS�E��/��#Kp���j�ѧ^Д�7��R� �ܙ!��#�"�'��睆k��g�u�h�W^��]�A.��\>�K�Q���9��㰋��t4��L�����ĺO$U(Θ6�-�VÛ_\p�6����_p�޷_,_fL I��y"3j�R01��bC������2���s����jA"�մ��lnj�ǎ�n彵L��4�/Lf��C�(BqY)��G1)��XgC2�⯤��+����gtH?^�'�q��������ո�'P=n��sYjM�>��u��6a��-BIV}�
55�hn�G*�@��ˡ����&�]���2�s4fL���>��꟱e�7p���rұ�a�e8��_*���N@Ϯ^-"�8�� ��NC]Cvvl�	�4�b$�[Y����Cɭ[�h]����w�t���>*����;Gs<���:�ضՈ�a����{�N��eO�$Ԕ�'K��<Lf�kxN��>�\'����%D�q|<.+����K�KMU���ޞ.�����%e̢+E����Ԍ��H�*��[oƛ�HN��5�3��ΙMs�:��EO"��߻�0��Z�x@Q ���FDCq����Jr��GE���1I�Yr����p���1}F�9�X�G���oܨs���B�9��pvt8�d$�Ӆ<��#7��r�K�z.�|>����%�BũA�=�؆%K�HS��[o�􄍥A37�GB'��Q�1�L�baQL���X��gL�c5�4�Q�a��$���4��A��Ͼ�C�êw�C��;��u�H��|@���q�T��U\oE-�NV}��;6�;Y�:���癘E�D[f�CC6���s�i
V�O��UI�K�S��0sm�p�=��J��x��� �p�gh-�I�K琈�Do�Ylp؝22Jes:#r�U S�f�h����=5��R��l|�n5�n�lv��b��M8�cp���7���/����k#�����~�G�Ν;��E5�b�'�!�S��H:Ё��q?s Z�v�dCie��%v�Tv4�v�:��DF���L&݆�x)����D�偕:lz��ס'��@$��ũ�-w�B�=t�HEFD���KđLdP�	�KCZ�l0;H��!KkH���`w�d������=p�e"�-��P4*ʦ^w*{��e�F�<3w��h����A<�1�|�Z���!Z&���9�t�Y�&44O�^� j��}���0,N�ق�L"	��fmo�V8��a�!1����(��0<4�����n˫*1e��=2hdZs��^&��̘���<L�S�D�����Z��!�o����9Mk�4 +��Z͠����f�Ge�_!���QgMymD]<��J��ɔ|��[H����_\�X4��_|Gs,N<�d��!�������\�4��{^|�i����8��D)�x�r��a�2����`��iF����W�P#!��׺�����X�~�
|Z�Ohi�qǞ�C�)6�/�<�,]�=���H��fЈ*Lb3�M��or�P^Q�E442�ں:�T�֝�N�X��kRA޺��a�y��J� ��t�<e�zJp8�)*Q^Y{�.�T�ו����݁�X��t;��
X�~�E��`!�ΈD�,�����Ia'�;���g.�~�k��{Ϟ�	�x��W��܄_^t���7mقu�����ːO$,
ྥ��V��q��q�I�c����G�#�M�h��.�MEc5r�A�#!M̆{'C���mm2Q(/�@:�U�5�u�2%�X���Y��ׯS3�b3(��q!�e�+��!�U���7Z2Ӂ+���ŏ�<��x(����q M����Р��y���ԡRОHA�D2��e����<��c��V�24�LA8��OMe9�&�M`��;`s�a�y4y���� ���8f^�.��\3Ⱋ☾�x�����[���q���Egg�tn��C�.�d��O�L
.K'��3,\� ���~���ڶ��i�m�8�2���H%����0��h@D��н���Q(��_$<
�Æ�������[C4�����sΙ�ŋa����T۝������DM�Ʋ2D���k���/hT�ԡ�{������뵋��y�^��Et��Ә��z6�];;���p��D����5��h߹N�/?��~�}ܹ�1W6��Y$�̤�p
yc���
G'*?4ЍR�.s;�|/z"��� �:�Q�ج"���m[�`���5�����;��x�;�b���;��زe'����tY�v�Q^Z&��ݻ��o�	�s�6�*O0��r������ ��͍M�|,[������	���L>��C�����j�i�M����N�~v1&�d�2�O+V��!�4)�Xl&��}�C�|`��f�rH׻k�QQY�;�&WQ]�AG갱��3p��a��~���^5�U�RL׌�5~��Zp���ȏQ�Q�;Б��iB�g�"��%A��I:	Ӡ��E>���5�G!M���K�QZ�T�:y!�t�Ό��N���W��,_���!��MF�'�uY.3�]=��'FC�0����4-�Q�@\?<��G�s��1�P����1::�ۃ�>���DKݶu+r�(@�И��)�ޛ�����4[�[�]�����U���,(F*�=�@���0�=���PR�G<Qd���M:�I�N&�pY[_�݁H"��]}ң��so��=��5s~���x��w�h�BX|E@ަR'��.R3�~���2C�0��dP�#ðҰ����	�ʛ-���2��9�YT^V�)�t~���v&Mn�駝$d���j2���)V��n*��R��䬙�$`���ͮ���w�N2��^:�F�1��@4 �AIY%n��.Dba\��=oR߉HP{��$2��U��rDn��s:U`MoS1�2PE+��1,r#$M�����k�Ɣ�A����S��߃��},f@U��:���� �%��":�)oEC�p�V�WY�8������S��[�DV��K��5|nCk�C�b��Sc�2io��P��w����jw�asI�\�T�������_��by�^�����ÍD<�F��,��]]�������_-'J��Ř?2�>��J+�$��.�͚��>���
^�55>��=�a��G�}Bڶt4"��$(�[f3B����թ�?�r���gs���Z҅ݴ���1�`�Ƿ�_�X��t��F�2R�2D��.ؼ�Vy*��ͣ/�DF��n3�l0�2ʟ�A.#�&;�Y!t)� �M"k�˜��F��h �QV�+6��D\�����3��?��B���gL�T����9��h�t!.�u�������fi���\�l�T�fo�qp�i�=Nd�9�ǌ�5޲
��օ�/[�0ז��O@9�h���ц|d�TV��IF���+'�z��/��A5��W�A�Ly���hᐍ�ƌɂ�Ճ�4P7}/4N���2H}5�+�ߚA�X'�!��j<�=��O�A����2����h����)��t�д�L�����7�JV�(*&G9	�Չ��rlX��|���4a�_��6��0�n-���X��+/<��}3����`æ���n2���^�r�y	i�B��&�7^�X�f'E�9!v'��d׾�PV^�yg������}GBF1�4V;�	��P�0��Mk_�I<D�q���= ����Q�P6�<hC�AU��n}�=*d�1���� ��I��f�K���V��3g���I�hj��U�Wc�ƍ����������H�^� fg &��>�)�����;�A�MȘj�\Fs.EY�'��]ʲ++.F$������UF#�������yՈN�8A�l�'L��m;�0��,�a� s:���EUp��&�yJ>����=�B��۰i�k�p$�Ғ�r���z쑇�N�ǚA��fֱ���ppaP��h��bQC�"�7y�0?���A����
�`0���Z���h��/��d�Z�������@Cc��݃��W��e*�G#X��+��T���/��9�^(cf�Ȃ:o4A�MJ������	��i����l�4b�aX�7�E7�]�QP�b34�t���3N������|��^{4G:�Ҿ�vq�	ˍ�U>Me8ͤ��A!#�jRIG����8J'㢇ќ��.l#�̙��/���w/֬�ZkL��&R+>��f8���4נ����6��IqI�4a�祻�m����a�<�I�1'��~�A"�k�D�jwa�=�&z�Q\U���qذ�{x6���x�/�`����D&g� ͛aѬ^h�F����aC���t�	�D&sn'�p�*6�l�^=��P&��S���z���睄�.?�]r�X���\�_i	£�'�j���[�b��Rq�s��PWRY�[��hF:�s�"��e5/\��L��:m�,}��s�]r`�Џ�ǢX{(�ۦgf�QK��B6����b��b$3y��41�h|�G"a�q4�*)�C_ÃCړt}&Ϳ��SE���T�s"
4����פ�Y\�����.��`&5M�o.�|�	��� P��i���pqK~�O��g
���F�$�{�,��*T�T`"8ɔ�&�_l��(h�v�����%^�%w݅?��'�%�6�5��fq[崽��\,t&�v�T� �x12�/��QD�AJ7l68ٸ���tz�8���p<�*���6n2�f�|D 9]W3(�P�*�XX{��:Z�<5�p0c���{3�LB	-l
��1�!�v��e������؈�	�j,.ҟ�98<�t<_Y%��NWlA,Ş�f�w�-�Kz7^{�� �Lgg��Ca�c��S,���td��.����`>��¦��3�T9��3q!��b��Ӈ:��S���>���#aQ��i	ŒY�wP3�����DJ�b��)�:e��T��9UcU^���a���`�j�;q���ᛵ��x�B�&3��7�U�{214h��3"�L#����CM:��ʉA"�r�E�-6�N7�4y�<C9������F�2@Z��chxX����6���@t$���a�0�e2l�RX9�X��'��=��,b���0L5���vIQV�r�5�YC�.�'�R�����T@�K,v>�bm�,N$��?��+̞U����Fw]����A��{7 �Ɇh"�O>����=�r�PYS�3�8S'M���5I��O}&���2VoX�2�y���{�i+46e��4Ң;5s9�a-�	�Æq�ԭG�y�դԿ�+�D��#����n�P3���F�A�h���Ysp��H�M,d ������^���K&"Rpb�9���T�M��a5�}dF�y��7�Fx�w��{	�$�L���砓�]�kŊ���ɠ�$�C����"�!Mp�O�14��[JWL&�˫��pWo_��;vvK���Q0��~{3Ӛ�+�'^Y�n��Bv���E����lh������ݭ����8l�B]����=�#����J�(-	��$����N���?j�o�A)������]E.�t:�4,�Z\Θ�0c�����2t���s3HF���!���8v7��.�TqҢB<�Ȃbx��,ʜ�%$�0�`���À�P�ݨ�~�%7$"�f$y��݆NJ9X�F3'C�<�r	�S�0^����Ʋ��Ia"b����`�N�2馱�L^w%^���x����*$�F��!ϬI�7%0M���c�Ư&}?9�<u�p
j�!ou�	q"D�����Y�桮���wFF�����[֠��ҺhY��^0:���8H-���L�w^��a⦠u5]�Vq�����((�)���T<�I)�!7Ѿ�Q]�~$�͞����.���Q1�O�2���s��ܹ��e�a|�,\iNB�)]��f5��X��,pr�GB��eqȬ�L�T��N
4�������͋�u�d�u���U�r<�M*z�٬,+Mѩc��y`�͆���P/    IDAT-iO98�.$�Q���M�e��� �)�6[�8�W]�l�L���(��s|Yl��`��@X�NL=KQb�5>_�~|���x�t�z�R�H'���o5|��p{�%�0,����!Ѝ�͚���YW�a¤���|���:<��cB�O8��H��Ϝ�32&t���l�JDu9����"E���pGe鲨Qt؉��Eaw�����ub�Fq�)��[�W6���7�>����!�J���i��]ohd6,0�;�C�� n�h�G�H����!�@���������9�1,_�⩸qX�0�j���,l�g�GIK��Ϙ�c($����p/�fH*8��d�y�	�~�� *�Yb:����_'�v� �Ӄ��h��BYm�9_�Z�ۅ�^{o��6���6X�劕��*d"�������"�*�s�pH᱊�(6���8ݢX���di���̸��)
���c�=W_y^x�Y�]��YR����	���]a��3�&��3,��^�տTD-��8�ǘ��9�B��~!<׹�2������p���a�}���?I�6��I#����,�9hɳ4ju;���!��L�b�� }9�A���U�N#!)N�(���Ee�`���Zs���ܛ���0g�}���Kk���-��q�%W��㪫�ZZ	��N�yR��]�ŵ֘��{ �^Ln�4���˔��K�	"%	�qȖ�c5'�n�}~%����g��k��m�z�q�:�\<'Mj��  "M��?uk�4����G���hfAj<��܃�Rg��'�8sO����=Q�qM��_v�AB�>� y���CzN|��>qy*d��:�IњESSLf�n��k��|E�%h�8A�,)���^�۷m�����@�.*k���04<���X�N�U֢i�D�x�M�<�.����O�v�(��C�Jc+B1��4r��`q���/�pl�8�ʥ2*��A!�KF(v��f��l��4ӡ�a��fB&矉3O�7t�ﵫ,��[���R�Q��v �zSX�|%�~�yx�Je$�yp�1G���@�ͨ���B��a$��7S�U��`TM�;�����ge&�,���{Lڐ�$�^���&(H����J�K���� i���d ���I$҈�2ɤ(��axxXkHA�V��e��t�d�fIY��>��D8��f�~|l�<>x+���z>�B��~�P}mH1x$	�ߑ� Oڬ�@�X��x�\�Z^�6"%ia�=S�3Ɍ�f�1������hi)5��x|����I�m>�4�]�$S,���X�i��H�翹��=1���X��7s�3yn2�1�$�&�f,�C&���o�픍������M������ф�����}�ع��6뮠���,-��U5�3�p!��n�W3�5�����2��'w�
�m� 7ͻ|�sb<Qm��`�c��90���[�*X�Ό�js�3�N�+ݽ-f��ry3��E\6�� �ۮC�Xs�y��������)�x��p���3����@��'���Y@���09<�ͅ�P�t�`�8 6!���bf��x�R�(���mfD�X�������R��Ț8x`��M����a>g>�������U0�cr	.�{Q^l�<ww�)ގ�ļP�OC3�_i�+���[bw3ȜAƳ�dL7so4���f��Ԑ���r8�f��'<G@� ��A�	&S��ps!���!U��9��`���N�"�s;(r���1Q�ط�{�u0}#톗���i�ʩ�A��͍i��0�@��C:��"#O9N��ۮ��M� ���17\s���s|��k��E�EE2E1�r9]��UTV*G/^��f�!E��n�4I:�H(����#��!N�j�USS>$B�z���=��:��'Qp&~�%16I�	QC� vM\�qIWe��&�\lJ6�tL�HL�FN�1�'mT(��3fElL�<}C��50�?��;s��o��&>�}эZ&N���C��w�/P`aJ�?ቺq��fP����x�0�f74���Q|N����� �?�湂�H
4��7��Bv�p����3��cOcx` U����1:��뒑�@���i��`�m۷㫯Vi!�)����	
���%5�Q����*X2Y�|����8��c��W+�ܳO#�"
B�)�v�<3*���9]c������BD.���E���`!����(j
�y����z���D�e>�Ŋ��&Lh�C��h2�ʺ&!��]�X��K�6��'A>�ıǜ
�2�H��EhD^��{u�P�3+L�,L.�6��9EZ�g�&�=9.�$,v��>Ài{-��B�|��S�u�����U�و��EEd�v�ZL�H�꯿Q�Jo�
��Պ��*�;�L����P��ѡ"0��!�q	��;��M�%K�ƪ��ݮ�&M�칍4V�r��3�ƆQ���F��A�幢"�.qV��:N��2��Z����P�K��x�����B#�;��f`y�9:��Q\͂�k�Y��ۍ7^{��߱��%�3�\�#��ذ�tP6D|�&XhR�gME�A��y��œ)�C�a��h�8�q�kJ��*-A>C.:�Ï8 ��z��r�d�H&
b^q�/X��u.��PTd���\�"|�z5����O�|\�`>����a�p���N��&|&E�$�Y�8xrcGgz�|��F�DY�K|nF��KNN�Dyg�H�=hX��L�Ϥ^Ǭ3��jt&M�$������;~\��+m���+��fD�8��?�?�A2��e������U�V,AS�8\~�X�������/QN���i8&�b�꘮����.n�J;�b��⺗��r�hhG�&��ҧź�i��Ȑc�|
���\��T�`1��h��ScKJ!�T���)�l���O>���,6���_p�/0i�x���f�G8�h,�Ǣ\8���vt�m�N|��J�1l�YxS@j/#A"�lN�����ep�^�9�r�9f�Ds- h4����QZV������ؼ�{447�i\֭[���*��kV�en��#�rP�Fð�r%��4_�?���F�p�5x��O���G�VX�~�H�4[��GA�6^ndlm���;T45��i�-�1��T�.��%r�Wq�
VF�@Ui{L�B{�V�T� 	���Q��d�x�=�Y��'�$6���S\����\�k+��E��d�WT� vKK�K���4 �<�g*��Y#���:ǍIC�DLwq���B%�E���@��h۰n���?�A��tJO�s0����DUU%>��6��E�~9/s@kw9ѹ�[�k��<;�dZ�R(+�@��)�U!Nӓ�qq�w*gP�-i���5�5�G1�)o�٭[��Q3��5\ �K$��B�tQ��Ye����� 2�gϵ;
��X30����&Q�A�T������Y?tS�S7��l�9�`����(����|V<�X�����ϟ��3"�^G-1�,l�L9�j'�a��Q$FFD�,.�.:�f>2��-5�3�>95��f,NT��)�Ofw��vجvCGO}3�:��?g�>K������)ލ�n��ơ~�L��%H0c��a�~�k ���a1k ��6�Fv��Sx
f ٕ1�������Dx����J�g�#E>B6��H�F�!� <ЇB"�ΰ\E���P�0�@	Lf���p 2:�/]<LdM�O)_�ƁO6��E��X*#�|o�.o1<+8,���{ל���Dw����~|�0w.*\tmoCg�N�KA��oCD�5�Dow3Hɖ�:�ݚX�>\#c`�7�:1�!����
��l�dބ�Ɂ���lg�Q8%+��k�!�np�p-�e����Z�f6��C9��&a*;�V�x�[ŋ�_� abq�)*gqeP�w\����������=J;�E������k̪�}���r���_�ȥ�B3���a�����qXpŅ�Fh)=�)��وy$�I�t.�_:N�E^l�څ��"�c~3�	��8�g?C0�q�쀉�D(R��J[d��2ʴ�;�X�a^~�iT�р3��e�͑I'�F&����c��Aĕ�>/E� �;�2��ډpH�p�� �l�"�e��Q�x%�hni��h�C�p�}h�6�x��C�Z��@�����Oep�eW�j#��%cɋi�:�`��u��B�׀�e�2��*SQBk.��OC̦fXt�BN���a�Y���}�"�aAeA��B&EZ�4�}2�Li���y8Ɗ/��+/�,)j�� N>�D|��ZرXD�j@w����ʟwx4�dƄ�~��.3�Y:R|�OÔ��Jj�X�D���Q�a4�,����xcs �'7z	�&�hTA#��7�Sм��a�ԻR7�Lº����%Z�8�7n��m���~ǭ�۬����`s�z΂A����N=7��"�:%���U��IWcC�z�0��y�X,��z���J=8�ģ�����cI��T�Mm*Y��G-��\@4μ1�F�����P���XY���58��3PLײDZ�'��@�✚&|M����^��D����k� �ͯ�H�45�:8�EdD��GD�#j�!�D�
K�*0�f457����hmm���v��V�Ԡ��C���!�o�QD�]� &Ϙ!����'N�a��`��<�w��	�z�/�����B'v���Rk��tR���Z� ��ޠKS��3Ak�a�66���Pr�3+�Uԛx$�b�3['�b�t%�"!%}}�GF1��AcOo�%�2h��Ǫ�W���]n��G4��9}��<�fdy�����[{�8�� )СTTW)�l][�&켼�L�� *4�'-5Q�ё�����cxW�ܖ��H�v�}k&�d�]�X�c���\)�'�y}�<y��ܹ�����FS���[U�I3f!��a��Smu-~�뫰a�6<�ĳ��o��[����6����g�Q����)
��7�F�I�*JUг�il����o�	�]&&S�Tݝ[Q�ƴ�s�BѤ��+��԰����YQY�0�M!�.�GY����|��څd"�۩���Hg�z\jV��v�Ii�3��]��1�<����r��*cTTosC���Z�(s�1�������5lٽv�/�f�����lUQD�nE�0֮]��e�D�1eH�N[��J5|�ã��/��Ӳ�T������꾼�7�t#���<�g4M�
�ݭ�6Ἒ,�s�aP"�EAdqK:��Գ���2h����wS����c�p�����!��	Q��d\��3k�˦Z��N9�����$*ʫ�p�eԑH�eO/1�DH\�&i���`�5@�=2�Z>�9P%#H]�h6���Y$4���g����(Axp��w`�ڵj46�)�.i�U0��n�hԊ�����j����N�<��H��c``�`*E�:߽~��O�P�V�/E�D�DK��8Q�Ԍ�hfG)hh�*R���R��Z��H��k��MZ�B������hL�a6sX�g��� �=XlŎ�z�� 2U��xJ /�ѡa1.Ȑia�YFWU�]JMhzFgt��dX�fQ\�Q��%Zf��������.��pЌ����Y��B�h!��'W[�=gN�@O��%46
��Y稻�@�ETF�wKx�9�z��$kG�FC`|�!ͅ8�s�i�����P��͠�5Mp�V�?�G�W��)�(�bԓR�n�)m>5���t6��.�X�Y��NLV�HS�ߓ7	)U-��La����Bn�5��p���t�#6�7�Dq6��G����2^�$��#�q�"��.��
�İ�=�e6�a��+)���B��i8���50�솒صuz֯Ayu9N<� �t�������QW-��˽���ck�݊Վ��
�N�.�L��gR�e�F4���H ZAώw�Qey�l܉βL0��3�
d3!�b'���~��Rn�O���B���A#g��cf*�,j�=�\X��{K!c�� 28���C1��0�PDTژ��W>��MTM�񂕯1��4�j�X0�)�y4<��;̈g���q�n=��/!�)M�xP�4�m㱓F"ɠjq�	�uQ��ǽ}�X��k�s���#����y�6���<j���۟�����eQHh
C����F�� \��IG�P�F/�͑�G0:ЇD����vS؄��L��Q;��26�<p�5���t2�Bh4��s{�8�K�Y��Yv�����?��x�e�.|�޳Jz/$$�Ы�����"(�qە�wEFu,�Q�6�e,3�`A�"�J� �u����ϻ�8���s�?^�@�Z�����<�s� �����aک�a�֝ع{�L��L�yϽB=x��E�d����3�ʼ/�N�h縰�X	V�)i"��3~!m�"ş҂O���f�IE&]
n��Y�5*���zB7�������F�F��D����)m)�j����0�U�ȩ� �<��5�r�=!.�e]�|~�dq�F-��&c����r�S�0M|8
Q�N�2eȢ�VG6�|-�� �:d�P)�	�Q�ъ��F~^��m�&�gӵ��0�*�PQ]���ls�������Б�h<��ۉ;�Z ��O� �%&�:�U�<���@aN�e��SV+����2�� *E�e�F�������V�)rSq�}ԣza3$��8�GTv75ȼ�4d�;3�̃�_l4x/�fƢ̪�Iɰp�42����ϐ��Ă��8R91�}��񚊯!�TmN�x�2?������+�`H�J!E�4.��-����ܹK��$P�I�hMMv��.�;/7Ot��h��s�� 
��eJ����;�5���Ά1���	����}��DK�a�@ln�< 8EWY��YRC40�3mN�H�Qe� ]6	$5l<�s)C�Ն��6���b�L1=)S&1�s����"Ԁ�0���WX(v�|y��T����Шh���) �ϵ�x�hH�}l���\,�M���$��u�O�{D�H�b��dg�P7�
��n��M��KAņ�S�:�I*�}�S+J�e�c�:i�4�*��'f��z��k �} c����l���C���f0M�l��f��[nǮ_����#��F[���ؠ#�� )4��h4L�@��>�Z
�B͖����X��t�%퐦<)�4��"Hć;�T������yQ�P��h��0���Eg�.H҄��HDNU��(�M�&0���4� *��ÈLJl���|}�47�QN��&L�c(�����>�0e�e�P7�mm�e�Nlظ^>��XpˡV�j�� ��lT)�J(��_�H��3�z�'�^�d������a���^��)5B~I�8��I8��$s�G���;�����kĐ���aBfI�ɻ��P�쐚:iL��M4�A\֏hv��l3h�nH9��2N��{�_��[#���ӂx"��FR	�PCh��/.�@�>t�$=�{>��#��я�(�l|���y�)r�`�#Å��N���k�0��b\�X,t:��3��)��'S�̀sg�D�ۏ�?���cG�'?�4�aJ$H�Wz6�l�9�bÂ��
)�����#e9�H��ڎƵP��M���@_w���v�%�j`���N��ض��L����}>YS�Ԫf�g���	^:I%�>��%E �
�j;Ԋ��#�j����	�Q\/��IЖ����Lё2Ó�|_M���{��%�$���Wi���R�d�I&X������Vj0I�'˅N��}�T�S���FO����RA��O���qc1f�|����t`"�4�2c4�c�D�L�f+.�	�`�X�ٌ��N��l�f؈4��7�����)e9\�"۰�`��G��Fso �!ꄭjr��/���)�Ti'SxNQ9�d�kH1;���I�h,.��Ⱥ�$�C�5���� �&��C#7�N�IaB9s����ޢ�1��Z��p������9�z�奥Ũ�.�uFa���_X�E<n�f�T��`�����|5&�@�v    IDATqr��"�D$ #�h?�GwmC^�gO=[V-Ǧ�+E;�I}yI1�[[�v�r�(+�u���0R�Ȕ �@�H�隝��O<dJ.ս�'����D#�HR�64f�4�Ai�h4Fx���G��tu�T�c��DP(�Աs�T,�Va�P���s�#���[���d0S� �Y�[��Y�����bqcN�2hU�2`���T5��s3UFD[c0���Sw%g-��0�������4i`L�a������逗�p�$)���7���Ŧ��N�Z�4V��P戸q��F3\tDc)�� T._0 :	)�&��Y�r���ƅ���lG��S��l���>��F�y�Ԝ��f�̍��&�~���DS�Ny�H���4��:�f���E �Hi�c��Ӱ���J'����N1�Y���WP�َ��g�1T�B�����A�A�~�A+�),�LM߫�.����J�$�������R��:�э�C��2E�"��DHoR�oY�B���l"F��	`��f�H�8JI���vF�y���6��ش�$΍G�,�ba�}�� &T��+�Bݥ#%?��k7~�ҟ�R��Ӊ����gC��C�ݡx��x���dP9>�ف��������mhl:g����v#),z�e���0�=��)Sz9�)��\i�����C��G� Ij��-(�6n
�uG;rR�R��D�!�-3��1��Z���&3i��Dg3h��*�4�|v�IT��s�fa!� D@��:�Ŕ-wu����@��ZQ�R�Î>�W�1%�����Rv{z�`sI�a2!�5�x�3��膟VCfr��[J�&�J1s���J
�];w
�����x!�q�FYWԂ����t��!䚔F���ĵ���[V>�j�p���42���|�����o�g���$��с�`M9�*�?��*�]�L�v��5:�t��M Ѳj�R�E�N���iC[��,�0X���J�M��!D��G�l�IJ�~N�LP���fS��ֆ��>�6eޟ؟s`ҋF�{��Y�Z�<�it�J�����C��=b~��	Y��O�1a�hL�8K���V/G2�|;~B�tҘt�[�R\WS+�A0�#i��?���=��$ϛ�㑽�h9]��g�a�8��C�c��\����7ނ�����?�wN�Щ#4��a���|�9���oC��7�!Ƈ��2ˡ���(��i�,X\K<|0��G�%#���8�H�>?�F:���+����H��c0;킌��%�o���r���	ӑ�	�U�_���=vK)�,�_lV�v��1��&���"'�O8��:�Z�>=y�x�:_��K���WS��/��g��S2���eg� 7� �N&&�`?z��Q^Z*밧�WL���zD��}ғ�%t?�tB�\#���>?�7�U��G��_���xI���1�2#��vR�h�x��-@K�ފ�ܬ(�ZI�V,{q�gޞEY��٣T�f?�o���4%3Â��
A��}���χ�j�)ꇨ���d
���'Q:B�g��H�S\ �l�ń��61મ��}���k�Ty�a2�$������loUu�Yt�1�@�SdЀ*�(�=�vm�O�~GR�QI�aЊ.\�s��JD�@�4�R�I(����A&��i��ή���'��vf�z���7#����س����ò��$xz���d0E�R��0�wQN���׫1�$cF��9�	�#B�g�DFYJ�4R1��Y0���Fň�A0Y,��	�$8�}��噬��1����X�v#~Z�!���d3y�T�i6��ClH0�����ZX��T���Վ�?X����Bg�!AJi��Ԧi�F�C%��'O����J���?K�A ��=j�c����(�aɠ3Ù�����4+�f?ʈK(�"�W��f�0��$j�����]�*���� �^��6X<��;s�ꍢ/L��Yj'Ҩ��V�2���Bf��$�WEO،4,���e0�A��P̤hP��SzN��1N!���iР�4W\<ե����Xk��Բ�����;�D0ž��رc��z���V���*�U#R�D�Tu�g�5��g��YX�Ƿ��X��с����x�f@"�Ă~�RQ�7�Ñ=��,'g�:�V.Æ�?ʶg�[QZT(z箶v��L�(���/DC�p���-YwL �N�*)4o��-�s�`d�P��I&u��5�faF�4��Ԛ���l� �����)��]'�A���?6�����:3,�3$�_��k��_4�'��j28P�ȡ�.z�H��@Y֊�0M-尚�8{��7��a���6�}=���>�L,����nG��"���z'q< �Hc�-,�q\H�]]RpE|~�H��(.tQ�͇�)-�&��g�ƂNcd2A���>)
v� ��ӡ��Zі�@[��
6�<I��f��Z|�Đ�
��`F�ǃ¢)��K�����ԩ���Ԍ]���C����B,����=�'_6f�Z^k�Ɉ-<��� r��G���JO�T�� ����xI6��H�m�P�������!��;,D}~|^�ڰy�F�ȷ�@�<�<l����z��C5T��H�_�q���Q><��V�~���I��D�AM,�,�p�/ᰢ�ku�G��y:��$��^kk�L�x����>�j<xP4�xψw��"�g��D^i�P#���I�YQ� T�ԋ�gמ������'ʤ��[�����!Sa����6�u�Lى���O���&��7�'�<4%�It�YTHq�oR����%��A�	#��䨴�\���H)R:��d�D��,��qjJPEO0GD�tQ���5�LҜ������f���i�N����RF3���\K~O�FA"�W/�oN�h�2��6��f�4��M���u��Z�&��'
N�WW�31 ��Γ�E�?�2~�.��}�B�3Z�� �cG/uҳ�`��ݰ�Lx�ݷ������s��N-��^cB��bu N��6=��_�:G9,y�)�8s*l����dãEϛ�"���Z'�F�(�&S�G��-,�����v�E����.E"hil���P�9���:�y��=*�[��\`���,F8lVx�z��y%ԗLG;c��0�4�@�LާDX�Y�V�͘�Q������b��'
p�A��s�ͩ�3�v������:��E;ŉ � ן����Á���'�9��|�a���#�	Cb�z�pÍX�jn���\�,�E�
�Q��ŉ�+��U�P�T<�4^����e3(�O�S�aiI7e�����i'!ӓ���JhMV��J�:�����wl�޲�*mi�Ok�a����P��v�贸d�\��r�I"�T6)�Y�x�{䚱�kkkǡC��r�J�:;#i����F�WD?���N?m����o�o�nid��{怙��X���6�Cѳ���40ڌ�|�p8"����|^x]ss�"-���z�	�p�i�E*�Ő�Z<��>|���x���	[�b�!h��q���#?U3��[\��Q5�K��v�(�ެ����A*�C	F�"8#˃�W]�s���,�c ��nVf/�(B�8�N��¤�����X��ט0�dُ��5b�p�)��36�m\��-�}"e��K���_d3����/�嗟����3���{�_\���:��n��5��E����y^sV�b��$��S�4b��Fv�Ƴ��%kaJ�}I�/7�8��(H��2BCcDk
g�E咝���oB��֗(�Cz-%U���Sl$)'����蠴G��&��d+���^/�ۏ��<<~��__�C�����tx��\.�4��|��/	s )d8\رk�4�4z�9C�Ԩ1�Q3��]��:� ��CGZ�����H��Lz���5����/��O?�_�.����2HÈ�����0a<��w�x�o��<������T�XH�Ý�����cU��D^�g��_�P;��'���DnO�1��V͠O̙�hD��Cwڙ�$Q����6=�I���s-�3
�aUr��V�`4�PB�V�&���_Ǹ1N)���ZQ��g��S_.�^��@��H�Y������_4�>�_MAib#����RKK.t2��?$�奥�Df���!�Æ�c�I�Lxk�G�w�vw��n҉�� ������q?��Jq��gbŪ��
��bFa~.�	fQ�eVS}���[\����
�sD��1o�3��]�C��8��/�'���������-�È�z:ҙ�%@h"L��Qډ��i�'&�����`���Rzl
5$%���)�OEШ8�"��o>X���l���r�T���������(T�_tD�'J{Ƨ�h8 /�QK|&�`w2)8�)h#a8�4h���c65yhS�j萙���V�ǰ��~ed�+�;/�յB�1H�����(�h�Q���P����)���f(n�l�d���M�`H�q�O�����a͇�ׂ��l"r,Z��;��W��Y��dgKs���%Sj���e������^x}t�����H3x�`֭^+����<���$p�on�VkE�BM�S�˦����?�˕��ҙ��1��ג�Q�m�U�%�1��������䡾a���fx�"�fHo�@AV�8�v��I��[4�];v`��}�o��σ��������'�T,3)��e������ۏ`4!cg{�L��wh�C��]|�*�<.�x6,�8e#=��(��&)�x�بpzˆ��1�����MMR��� ��Z-�YD��FZP^i�8vv�B��J38����އ�7���/���Ξ1z�)c#T�8�'��F�+�fPx[4(!�&2�Uj}U�J3��䍣6�D#!�
�2i��sb��(.�Gum-�ۻ������I/F7�HpBD�6��B1����<|D
L1bɰcĔ�\S�Ն��V1�/�&e�����*F
��%_���`c�.M������v%��=9r$\N,�Ǘ��J�o:�~���ӓ)4P,l*h8�	3AN���r��&��CjKvn�4�=]����R�x����՛���ՙ��*�ܺ��N,��/��������� �+3�~���
oLZ<�k�6NQh�D"��6��%v����g�>#�E��S'��+/FŠ2���b���F*�B���.7v#z���Cp�ضm'>x���s����>�9
7�prr�q�p3LV�dw������5��<t���Ɔ����c�Ɵ��q�UM�V��f�@}}��/h=�,�D��$-�����Q�����M������h��>�f}�����?g#ȯ1p��˘��PC��@8����ڡ�񆛱z�:�t�̀;WED�tk�n�?\S�@r���Vi0T���
ŗu$n*�N,�#�&̆�н���sg���4��&��������qH�K��e����43��ǎ�c�����~��.'O���.�/�i:�r%%u��Of�N�LRI_�T�����m[�� Qb��fApʠ�3�g�v��r_~�%E����֫�i�!�+����s�J=�p*h�CJ�� .���M�S*9/(���J秪}�`6I���Q�H
Æţ��G/��<X����F���4�K1@���� )z��f�u��,E� �d�3F�왾9�X��=�z�`���b�ٷťe���I0��,O&�z�l܀�c��(�p�1?zN�5�! SiI<z�z�s:�x� ��~�2\z�h;ކL���%�2�$��e;�}�Y1�ⴕ�?i�l��N#�����<s&vn݂�7J�L�� �)�ezM2�g�'yf4ţ�K��%�A��Ԩ�u�l�2���7�#�?�Y <�>4�3議9��0:`�)�ɓ��k�"E1m�g�l�sl��6* �F(�ԯ��f�Ns�����3�ZNfJD�����gl�ZR����~�X��A�oԏ���l�m�ک � ��yB'�u�@�ăQ��s��ۉQ�F����]�ؽ�1h"��jwbPE��R|����1v�d,������W_��1��ۘ�_�$�$���x��Ga����[s=@#-��'c��t��	�O'����Ț�}�=C+�uI3(b3yn�ǘ�/�+pQj��@�ם�3�A��kV!\���!>[t��V��	`���X�A����瞹��X6q\����hG J�f
�D�_(j�F*l"ԏ�<7.?�t�z���'���L�̿�c�h�l:�f=*ʊQ_� ��'��2x!�O?�+���.C��z�c�X��7�JT�7�~�׮�c0g�<�N����p�H;,6��#��  ��v5@um.��b����X�byZΡCvN�D�� �C6�tަ���C����e}L�>kt��l��ǐ�s��p�x>���@U*NJaEљ�K�%t��a�z�4��y�i��_6�b��u���gܗ�mJ3�����+�o>���̿kO;G)�?ӆ�BUŪ�w��/,Z)P�f��I��6"��X����sZ��%a3I�$�=�����6u	�s�޻���6n�֘������UW̗����a7�G��^��ďҰ�B�W���ö����������A�P�1(��^�c��Ӓ�)��4��΂f�f:pU����&v�u5n�S���^)^U��9�E�\���Nt�z�]����4N��o��oPU��e��1\6g>�$��L��S�|��K��J'��r��(�=��YY僘6��Fc�1V
�t��L��q��y���+.t�y5"s�aπYg��\$��/ ��*A�?���?x�x!�W
�/��L��\��1���Z�1ď��@]=�"��n�w���dR��� '1zA��%7�W1j��4V���vG�h7�K뻈���H#�{����/�k��=)�t�6��#�̑��/Cu�p��l[����x��/�h���F́%g8���VP��'+M)T���XŒY-1���Ab�/�E��:̜q2�N�\:vd���s:�0Y�+����.*δޞ >���طg����f���k��.����������1����>��v�=wa���i�)����R��bMŇP8b�i��jI:[M��\��F#���J�?&f1��L֟�ϙzfx/I���L5�^ѫ
m:�.�.��ǻ�`vdK3�g�.d��X��;���e�e��А�#�*Ê��t(�)��А|RA�e4C�^uOӢ}e9&�p�����Bے!\s�|<|��ؿ�	6m�q�Dy��,���О�.o>�����.y��PԸ���G��I'OVN���PI;{{�a��lD�`\�˅��<1.�0�_���
-��ZUq�"R���[20u�i�%����p��0"���Zv���y =R��J|��'3�G����^�C��LS{G�$���}���83$�uPU5���}�vyPQ17�|+6l؊���jMj���.\(U���/u���쏤�QcG�	T��\OʥN&N\4	�i`g����p�m������g�}�$Cd���a�<��S'�����쳿�nSl:z����0�,�������]]hn>"`��	�n>
�Ն�s���)�`��[�k�Vu��%�����������N��Ae�x�O/+�3��C����rߵ#�nWZ�hR�����>x9�t;%7@gaF�ʽwI�&%� 0��8;'G2��L	�¨R�G{ �}�=]�4��@k�It,�I�FCe:�r�e����*�Vi4�L�>�T�M?AAe�������,��[�Gmu!���Z<�_3�����FSN��������j�����n?����Q]]��b�jhi9~¬nܘ�8m�i�j������������၇��%:mR���,��P���*�Å^��[�`��5�e@�nJ��b�1"��b����P��4 )).ێ�.59���;O�{��L�X��PX��y��ꉛD�Y���*͘'O�Dwl�%M`� 5t�����x[���TUѮU�D�t��    IDATGa� D���i�L:�������\�i�Cl�������7W^��aC������Ϗ�}�7�Z���,�6c:F5���~��bDGʹҌ�`��l���,1�[��ZlڰU·駞�9s.űcX��hoi��I�h�"|����/
��Z>Ƹh�N(1B-�)�ĈQ#0n�p����B��oi8��p�uE�DY9�2���d�5�Z��xm���~�yT�ꔇ�)� V�K��L5���И3��_���um�i��bn���j�dX��su�+�nN���^Y�0�X��ĸК��� M�0���T��玴g�N����fϚ��#�x��{p��ٰ���p�G8v�0���g��ΐ�F��f>|D�|�{tM�d�ǥHL&�TW���/�b���7n*�aɷ˰e�V�;��]):�?��>:�B0����ar�6�>ő=�жw���e�]��-���˔�GC'n��=�<	Pr�K�!o����V_�<�fi��Œ��ڐM3c�xF� ҠS\ue�Rة�H��j�i�&�(6
#�"l��ǿC�)O4���z�6�I��<K��ɠ��{SZ�V�%��p3T��'�R�����50'�~�=W���B����~4=�L;J�l�� D"A8lhb~��mZQ���.@��;6lFW�q�|�v\��$���·ǝ��c����%}��UX��B��FTQQ�)�OE��%�(��0�%����+�y,�y�8��(���^@gk�2���(�T�ԅ��|1zsscs�v{�be���\�/�Uχ����@�4��y�"V�n*M�!�������r=֊>o 6���\L�2���o��]EU%��Oe0��~C�lTb@F�]OCXI6����Ղ�*�I�L�C�m�L�ғ�Xȏ��L<���8��������H�!DI���PVR���.��87G����V��� v��/ׁ�<��*//U7����B�6"��r��)�Y�Ζ��'-��A�J�]E7�s������4��f���b]�1�Zc�H�̩�R�y�rRɍ���j���C��"���*������Ⰹ���Nw.�6����e�v����������/W��,P��U�+�z��IL��6��VQ���(�Uj�K�BFԹK�=6o�i�����3������g�ϼ�"ʫ*���H��i�Q=z���X�\�j���@Y���7[QXQ!EawG�4���>9��A���J������c�����SN�ٳf᱅�q�:f�YK�y��ڟ�����Ē%Kd�q"h2h�ㄅfJ��ڝ.���E��>'����&�	?���.���?)�y��]��!fKWL������M�%����������§`�:���T^�39�S2��Vψ��lu�H�}P�s*�z$��E	�Y�
C��e���k朏��Otpg�y.�;:ő��v �z�`XMf�Y�Z_�8ҥx(�v�떓�S���H0�Ζ6�~�ˉ#��ށm��`�bx}=�z�),\��/[*�F��RoN)��p*Æ����SNÔ�O��o����%j�M@�3�_��&ٗ	f,����� �n�f�,Iy�I?f���Dç�͑!�r�E%`T�͞���b�z�o�ko#n]p/\9E�[ܒ��{Ţ��đд���@W�b|�)�'�@Waǂ��	& E ��-�#jb����	�p��w���xx��4[�ɗ��Ν;D73���QUZ����c���ضe��'L"��sQQ1F�-�H4$S+��3�̾��3�L,~�<��ga10{�<���kq�m7c��?��.�saIP
A:#�2��SQ];/��'��qۧ暑SԯS���#�C�>2=Hs����r�T�� wր?$�J�3N7�x6j��A�%A*4u�U�������e���Ko ��
:�M�XI�	M��2�R���US)��4�lIh����f+�,�(5�6�>I��`�g��07�x-�����ߊo��^�����0�)�sх0poN[͓RH:hkG'��YF���AAa>��;��ҥؼyJKJp�E���.���{���dgf�'�GǛn�I�c��)w�7Fi�B!?2��$�u׶mX��7J�Kc8JV�	���q#q"�!TUU�Ý���gef�b�	e�� �`9u���4�� �(�?�ćTE�E#}�`r�������h��#�v��.���#�1��=�I��y����K}�����`�a037"���<�	�o��q����o�U��Ƅq�q�uף��>��oذ~�s�1��98����>lڰY�w�'��Q:l���=Ê�c�t�W�b��ݨ����9�=^<����2?~<~����_��/���/X5�6�4`�P��Ə���ax��g����W��|>��K�Pj��+����g�<�O���Tւ<��qL:4�͠P�Q�ļ
���&��-��u�����y8i��J��X��A�I8,&��Qt�i_���hARk@8Io�lF=J�Vq������jk�$Q�m�EgNF�����k1��Y9�h>����Q��,��_5C���>���?���\��|�l����f�����3fLŲ����߀���)�t3���K.E0�Ǜ��m=�MV1*3u��s$G���hݽ%��1���j�R���P )l/yX{��=6C��Ύn���~�1�!�'�*x�z��0']E��M�ө 2L*~��2(�B�~iG�b�XD��I��`C�� ��on�� ]zb�I��r�"��7��� ��N�b�*�D����&�R(���!��Z'�,�O|��'R������҅��9��|�����[(!Rhj��H��!%͠����*��������+�JAɼ��(����;�L6mٌM[�H���� :�tR�ݪ�����%���=}�|(-���Ξ.�߷O��ο�R�>��"kjN�i�FDx�i�^^Aǉ��
%<ﴂ�W6����P�͖�ѐ��R�E$?dl0 3'EE%8�F������a�I����~��q��}��<��"�޶��t6�6���2&�Z�8R@yp�� CW5B �K(A��1���hǀ1	c��mA_<.��N���������cž��*�=]�����'�����b�*i!���d�F�#f��'d�A�X�7'�'�c�ڵ8�xHУ�{=�t�zb��i- z|j�$'�K��V�2�VѬ2SH�nn$�G��� ���G�h�t�S�7m�+"��*,d�a�ֱ�1��@Xnm�+k��ޅ�M�(,.��E�!��⚫o��h�h�q($5��z�q�U�+'|\S�Q��I�ÇQ'���H�e�D� �fО<�߃�O�n��?��nބ�Ν%M޺u����1v�X�8uz�{�i�F�����xb���� �����An~�P.�oߊΎ6*/ìs�D]}6����i�'�'L;��sϿ��V�RF��F�P-H�� ��Vjh��������5�x�}2�S�`�HQJ���4��E$�`���&iͨ���e�٠ɒ1Í�a��ب����T�����׃���V�^��^~y�� �p�R�h�=��@s�dJ3(@�]�)uH�ս�@�
�����l�XQ��?Ԙh����iÙS�c�3p���G�W^Ǫ���G���B\�y����g�)��3��
N
8���D�Pˠ�	H�����c�D�~�s��x�'�{�Q̽|.ڛ�q��x�������!)��$f��Z�L�'&N���'���^~��j0����R��92<��y"��=��4�iok�QQ2��`i�W�ҙ�ŵ����xVO2s�]�K����<�~��8r�ϼ�\9�0�3�H�sj�8͒����r�Pb� *QDC�H�3<�|�5p���t��lҊ�U$�miW�a�W������w?��۶b�G���Gq�C��p�q�)'㲋Η�6z��N��̽���B{G�䙶�����bŊ�p�3p�-7�+�᧕�1�����>��p�ͷ��o��k֊�߫�1�)1a�E��)Ӧc�����/�F����m�����gW6xt[�	
]i�Aw~A�'Z�ۄ�O:"'�,"@2�Z4�
%-�E�٢�StFW��G������ŕC�7;��Ha�D*�t3��#��u1F��4��h BggmJb���H��F�ŏ �����-��U��Aq�	�7fp�e�aǮ]؛��O?W͝#g��͛�T �\����a��iS�*�l�����i;k�LL�2U���{k��Dm]|�a�8q����DV2�c���Y�2|�&2x�sq�Wb���X���R��^"�OŤ�#���P�t:mkoW�h���+ϔ;3�9��a����Ly_4��Y�Â$�:B�8�v7��h�n��5cfƕ�3����/��U4F�v,�J�P\�-@RSs�?&y��ٲ�c�Kȼ�n'�F=< ZT֕��W]t|�1��0i��:�llټ	�DOw'�;�ͽSN:?,�o���4���r:�:�Jn��F���~�7,^���)Æ5��܁�q��1�;��s/>��x���%k��1����3D���� L�&O�(4��~
6��Oԙ�����,P��LȪ�!�ī�H�������(P�N2��I&�l9��>��@��F;��|�ՏE��/³��EN]IWL ���m3��"C+��2�G���������*Csk?���l1���sa�i�����~��wD^�ͨCq��6v������s��z\�\��l̩(jj*�_\�EO�?._�sϽ ��
;�MaWW�Ej:��SO�ܹ�b��}x��wE��u8z�8�=t�|�8�4�2s����O�,Sq$�~XZ�6D�/��[\���:�}��˾���<���2r�I&A���1�>|��cd���ƒ�����e�6.ʄ��E�E��@lc��H�j�l���c5��͠�U�������is�}<Nh`�E#GZD�"p�I6/p��$�a gn���_�P�H�@~/����Ks[�Y[����cD�ɴ=e6_"F8ć�[N���ҩ��Oj�S�~�z�a��!x��������W_Ü9�è7���B+��b���QX��CG�����#BB��!o$;w"�DC��k�N��)+-Ɲ��99����O��믉���s�Ą�'����C�F��KC�G�l��rbt/��
�f�LZ��;���q�kĞ;����_}��gf碨�=�>(����_�1��aߡ&lزv��ٸ���B����'� �=&S����HA6��*�8�rd-:dNMT�h��G�C�O)ٸH��D_o����F��DE�n!�z��(�v��/Fqq!�̽kV�ƆD�UW[��sfK��c-��'��������粴�T&��!d�z�̙x�ߡ���_3֮Z���\����bC�� ������'�b����f�U��E��	�I��/BGMOMx�d��;M F�b_,�9)�I�`s6]z�j��F���b�[P���rt�zq��18\v,����o���'��ff�M��|R8k�D�Ԕ�kL��z�MG`��K�9�9�jv�wư]�h�l!���#"N�,tB]�__��n����Z�}q�m����_|��}}B��y�7f���G�HS�g�ׄK���x}(*ʗ�����9�t,Xp� ����[\�7�D�vh~��Sx��������U�ƼBg�n=�Պ1�Ơ����.Lz�(*!����F Ac@X&�zAPI��v��7�}�§�t�~@��Zc�ɕ���Jq��PƑ��*�3;���K�?�u����?/F��zq��@?�kP&L���g��
�d2ꅅN�Y�cn7��^83�J�� +3GփP~���RW�$��a�đ�5}��.�ܼ�߲ �Pk֯F���d;q�%������'�����aGoO��f�W,؝7��è1#q��������?�-ӟa�uVW����x��w��%q�̙x��q����|�\��*ګ�K�GF���O��	c&�7�@K�����$l���P4�4衫n����d��+� u�D��5��6;l�8f�aq5�h��������!�lΕس�(�|�dT���B,EݔA(R��1�
��d��`3�6�`_2���&tw�@�ţ����6�,V��ֺ���@%���k9��q���{�ϫWaҔSLj��󡣳K@ȹ���o��|�֮^�É�>��QE}L��_$#F6��;o�߿��=�Y��%E�t{`5��n�O��S�6�ƛpѥ�q��w����s���*[S����Uo��3����x��'����v
X��0�ʡ���V� N�XX����m������1?ܫ8��Z�*ͅ��ٜ���o�11�Ō�V���xx��X�f7^x�]dV"��"���l���h��F�h=]�1ib-�Ֆ�(ۅ����ۥh>ւQc����������B4@��?E�hm�a���gO��`OEq��i�����:[�c��D��Z���Ǎ����6o�#��/��v�8��x\`��{1{���[{��}�N�~X=U��={���D���/�Hk�y�!-	��8M�ď���0�8�K
q֙3Ѵw/���g���X��6��j�
�7�PSS�p�N��V�d �@���[��\��p��*>ɶ�e޲r�U�&tgnTo�������m��?L}�E�%�5��A���D<Ћ��]|2r3�����vc�O۰u�>�w�H�x��/M�0l��:e��ѷ��Djw��e��撙�<҄k/�cƌĘѣ�<b���E�p�磡�o��&V�\���N�����.�6���@��O.z�F��ͷ?�o�-S���C0i�d��|烏���;�����}
�'[09`WWq����A2���D�7��W^Fg��0uE��S~�{Ԗ�����i�ɓ�<�3&q��Ȑ:� ����,�I"�-����8���92;�w�|�DL�E9�ML�q�_<�E��g�G����ϰ;�(��ƞ}ML_��ێa�w+�����Qu�4���jCvn1�7V�ٍ֖61�)δ��3�a߶]���x*)�@u�`L�8%�Y�Ldf�`�d��O?�u�6`�e��"�Dp�����\�S�L��ٗʀ�o����[䙼��ߠ���k~�'�U\���,EO gv��2�K��MD�~�(��	�ӍsgLÖ�a�eiݥ��`�ْ�I��w!+/�u#`u؅:/?d�����|^��t��*����6�Oh�|f(Y�/�ހHJ��h
�C�Q5z<��8DK'����f�1�@T��j��MU\�5t�׈S��`�8-�`R㯚�H�S,�Ɖv
�N�������)��>05<��5����_�f�� �-�l�>($�d"�&3��FHב<R̄�ĤQ����yx������.���[�Js�����'��~�A�d��kk�èU�g"�����\�]�w�O?�ċ/:O?���^����xo�bq�w�U���ó�#V��}�P�t@�"�����P�x ҝ(�J�NlYP��������Wp�@3C��H�˝�2�� !J�ܙ9h9��î��b����­�j��E��j͂ќ!ŭu�$=M�h�&��J1�%�@�&�V&���q^A'$�!���MqD�D�bB���^{%�*�U�]	�Q�s�9;w�B��&���'L���b��X��k���L!+�#�n��~�4����C�x�'e�q�������҂k�����DEM5�|�q�Z��B�+�~U���U�.qi��ɓ�K�(!�VE�-�J�+N�7�������aG��%6K����tCkR͠�`AnQ9J˫����Б#b�t���`�yp�}�����B(�$#1�>��I�    IDAT��jR�B�zH$�����v:��ʐ��������PRR���|#AjjZ����^4*��w�O��y����1��3�,���ro]�,Lo��F:�/]*=�
R�$�M���"(����ysq�����hmk�%�\��W����/�����P8�����{x=�V.�Z�Y���7�o7��H�j���(+)ħ}(�����#A8�VN9�e�+�4���Lj/ztvt�)����ᦍB�N�!/SK��&��%%�}�86JU	jΩɟ��~ڸϼ�&
ˇe��nt�U�>T�(�(�$�1\���ф�U���(��Č�(��a���df#��Z�#�����.Ӂ���1W^<ޱ+�]��΃���E��2�:m��;��)�"�3y�����Š�Jlg��$|���O��W�ƻ＇!�Ce?[�l�����h<Ԅ����{����Ǫ~�����4�P�m��
�l�c���pҸ�x�ͷp�*63��8���e��{Cp���U�Ϝ�2�Α���;^~�#ut`]�1gORk���M'^���b|O.�|>���|Y����r@p� u��$Й��/I�aJFp��8��Qp;���~޴E4�d0\s�|�U��.�5���w>D�D�Q�I��0g�,��Z4�ۋ�ӦCCj��`N\rǦL�K/>�<�$�����1��f���	�t������7��a���?����Ïޗ�,5iԈ�w�r&.[�#��>�_<�=��n�)@�x���e���=e�D����+/�,Q�E\|	H0 0@Ͽ҃k4����p��P��F�P5�Ur�pbs$�x��E�V:�5N��$�s�f"���
+�p��������k���z�1擆�eh��Y4Џ[7�0��zt?�L����_��3f������7lڴ�����+d
�|�(r�D����Kqh���s�9(-����V���A�#9���R\p�9ش�g�饗q�g"��H藼^\�[6oĲ�Ü�/��~�8�z���+�`����T^>s�]���b���w�|�J,z����$�񧞁��V��[�Bd���˨�� k�'�CK�!,��eA:sA�\v����1�΄�!�&2@�Y� )�<�y}r�)a�|8ĆT|�e�+��j*X`�s3�H�j��NT�Sf]��V���ވ
��K&s3u��s���`�ʲp���b�ڟ�f�J�>�d��O?��f!����O��@(������a����·����;1�9ڄ뮼ÆVu��TNv�3��r�h<����/���+�_)�ԭ69,��W__7^~�i������@gO?�+�qݍ7���-z�D7/�-֮߀%�|�������YB�Y4�����;1tp%F��o�oW��l���A�������VM]�	�HňR4q>�ݽ���׸~�������V9����	�I���2T�:	>���r#e�J���l�#���0����DM�`̽j.v�=����9眆u;�b銟`ue��+��"�ӦO�;;K�߂���mv�d;0{�8��y;��(��EIQ)�UbXM�f���?��+Ƈ�o¹�\�ѣǉ�]�m$��X��;̚5g�u�w~���n��݁�g���[w`�ڟ0q�8J��g_�?���b��8�z�P����ơ}��9p��b���n��QN�pT,	Y t��:�>;�"��Ճkau�Q�$@&:���v#B#B�m��K�9{�R�����x2��5�%x�+CV�P?�]�tb�TQ������8�O�y��	MJ����.�9b�d��0����A'4R�~�&i3K6�j��&�_����fPK���()!�z��xQ����)�`20B!,!��-[-��q�'�h��O�-G�=���G����/X���1r��ԏ� ,,�ǥ矋�~Z�w�~z�p��C:�p��ps�j�|t���iS$����b�e#�i�3�=�e?��/Ƶ�����~�,�ۺU���@��S��(ĺ]Y⒏�����|&��<b��(�!�?�y�jZ��ޘ��X���t#��D���T��b�R?|$��wa��&�2�x�q��"�5�E��b��`!=ؐ��P�ziӀ>'��x�b���J�q�)�1��
�hV��ތo����1}�8�.i�(��q�J����3Z��EYn�_2W���N=��F<a��1�����׏>�[o������dGD���G�ݻ~�"䩧���/�(�t��{ec����a�����ܸ�G��م��IgS�FIq��I ����2�I�8���Ã�\}���^D�^��D�{%��f����w�s�h WR�A��[l2����)N�|�\��(.�B�׏��G��q�λ�h��]�<���iy��|� �}3�[�D��&�C2�Ù3�`�g��X���PP�~����|Ӎ��˄?؋}�]���o��t�	jq�W��������F�D6�h:��ܸs�o����{�G�֘��(	R8T����*T΅��a��o��������#F���!���S��|2n��.<������zX��2�5�j�?�!:��Q>�97�^��'���X�N��$E�Nz�dlI�NDp��� f@�; ڰ@���;$��t��s�Ť@�Y�(���v6�?o؅EO����t�Ii��z(��ʃT�cp�J�ý�Y����K0bX6��:,�f�n�~�5lټUU5�2�d�z�$|��R|��[�!h;҈sϘ��矆G�˾��c&ؐ������`�g`��	���{%s�0q�4�Ǝ��M��U���?˳��'�k��\�NXD@W�X!��S�㛥K�����=����"�o؈7uz�lr���F=eH��:L�0	'���w�|M���d�̳�(/�N,�~f4�Ԩ�i?���z��~4��>��^`8���:���n�ߓ_����MG��~eUCk�F�}5Q,��c�gc���D�X �`?2���M�{�GY���k&�'S�LzB*%��{�ޭ�t�bł]��(��(��T��
����!	IH2�����w�ާ\����k�}�[���>�]��-�8��d����߈��O�nظ�;��:0`@W<����#��=�����w�mF�=݊1g�X,~n~�v�@x\� F3����ӡSI;���{�n�W]uڶ/�\��={a߾�=��8�f�o��:v��K��S�Q�Ѥ�v(*0�K�^E��=q����[��ęs�-g��m���d�\-}"��ؾ-�t��k?A��b��7�=�PW�#I��l2�g#+9q܌�)EOvf���R~�f_@%���P��"��ty��H��ym�`�O������7?Bf���3%��B	� ��
�u6�}�7����~��ￋ!��ډW�ݥ�2��x��O�k�v2 �gL��Mߊ,z���f�D�Y��ܵ��	�5�Z�;�q���������Fv��%��d�$����97�P�^�����|�zfϚ�_x
g�Ta���s�.\��i��B�NExg��X�b5�=�8LI��ʫp$�J���G}���E�<���h��_A�M/�|��_wɆ�C�;#�aQrx	�bp�WSލ���$�W�t`�����D��"���Z\>����v����#�b��
��8��Q��A�)���7�iD�6��u�X�l���͹	�'\��o,An�"�9o,�g.�!99W���v�x�饲)MKIC�ÎW�A��3�e��(.ꀼ�B�^��ʒ����S�ӻ7�w�u���&i��Q]W���T\���sh���q�������JK���?ɐ���RG�|�mh�{�p�b�l6�1w.~�e6l�,��/�gR���O��P��]J�У�k>��U��O����	J��HLBa���3���Wr����V��bɭ<��p�$�$����BH����_c�)�9]��E� �.�H�:ŉ��}�j��G#�Ħ�Ѷ� �����_˅�0y�$���_��Q�	.gF�o�.hۮ�?�}�!.�mT��Ӯ썃;�Λf��C{�blV��#~7R-�ܵ�r��܂�{���ݻ�(D�0�6���gΜ��ٳpՕ�p��I�TQQT�܀��݄�qդ)HmS���~����%O'CSU$ ��.�<)�����[�˖��B2���4�{<��wB%H8E��<��A��
 �[��EN|k��L0$?�4����� Ɇ��{�@d���-F���&��HY�
�9�k�J�)��&܄���	m�� v�c��рx\N2�~_L&JJ�A��[s�b�������4J#���f\y�:%��:���zu¬��q��Q��!t(j�U�~���a���S�t��b�\�o������w_~�eK�@ANR�S�CP�uHON��q��/��'��s��ҭ���fO!v6�ܹs&y����f�7���+*+���cp�hv����|�k&N���_�Z�"\Y�̕0Y;�-O�%�]�Js�n�T��dqM�	62�{��IT�߭2Q�US>O���dĳ��FC�[b4z3�	�(-�ڦ&T�<-�cJ����?�
��D�Z�B�`3��5�f��J3H: �uG�	��:��a��}�rӐ�����6


1�__��c�###�V���w#'+��9�vn�2U������
-�W�n�5cV�X!�����g��"�����B�c�ZSS�^xA�/���O����Ƭ�31f��V�_�{�܇�~M-n����B�ĉ�y��4���G)�@D�a�a�6�A�Ɉp�+�J���HFP/nSȯ,<9�ܾ�c�7�
�O-�kz ��,�f3�Ԍ��JdLA{��u�4�IV<�����xp��0���1��fQ���fPǠk����G4�E��Mԋ97NA�)X�x)r�1l�(���;��߇Ç���cb���9ؽ�+�/���^]pی�����톍(�P*��|�����y��q���EVv6���#~A�6(7���/�DaA!{�Q���`��oq��\�d��t¨1�Чo/��Wc��3����{�+�|�#G�)YX�l�����g�M�ǫĊ���b�a�/?��&��HD��0d�Kt�l��Q��!}q���Rp���Q������a����lBRF*|� �� �vr
�	����ͷ���
,|e��J�#�W+�~��I���K����h��D�݀'�u�'p�-�С�<�]���w�Ô�7`�u���b������ϑ��'�Hc�Ę���ؼ���ǟѡ{7�d�e�Gi�<�a�F����{�����1y�4��.T�CQ{���Lf6m�,:.�g+/b��%�b�GaA�|�������Pڥ3n�}�y�C�<$~#n�)!tv8$  >;_ �:uB������p��QX)�%)��f�G�F���Kp6�e�
��ŋ�˓��F�V��ll�����"L�P!�ဏ��h	�Ih_R�Y7���O��EK���:K*Z���F�H�|�2�H8�@F3u�lv����p׭3q���A��X���8|�����g_XO$�G�~;��ҥ +=�;�b�5�������O<
�������B���e��[�.xv���v�&L�4���jtii)��a��u�QE�j�J8��~�)2�2dj�ՙ0v���`�y�\�m_�;��}�H&��x=�Z�}�� l��#����mѿgW�Y��4��=��#a���ERb��.�գ��I<}�F�A@^T&�ӕ���9��ȳL�J(ͽ2"{��R��i�1��70���?����#�}7�5f�����E����ӌ�6��>e~�����}\5��r�,,\��y�^|���bS�ӯ&O�����ۈ��b���z��8z� 
3R0q�t�O���o@��>f4�����%M%�ݺv8�˖I������D�d�TT�����	���k��¹:lٲY�{ƅ��:L��J��X�.v�ދǞ~ѿ��O=� ��$�т���/I!�/��ZR�f�>UgN���ݭ��?���Dj�^�T��@��/���d�Zbؠ��a����<h�c¬���4�� 3ҁ�O?y��D�������_�`�ORە�sa�]��Ψ���P��T�wN:��[�2
-��R���	�&O�[�Z���j`6�0�A�ҹ�.zG���i�IM��kƢ��	̞|-:��aʔ�r�P�t��y�*9b�(֮]����t�|�{�v����?����:��pzu/�w�����x
:������7�7�c���oރ�t�W�A�����D�o���9�����>ݻ�U+p�X�"��R�C�NJ]HxLBj:���I�́�D�p`M�YHY0P�b`qo4șEH� �X��C�tl&���}�f�g�.� �e�Ь1#g�!�A#cS���]H4�a�C��\<ۈ�4�d~���w�L��G����ߡ�ؐ`1�8ρn�p�Tv�.Gcs�ə��Ȱ�1��A8y�n�5�;���h��,qba�yYi4�
�w(Ŋ�k���}��X�D:�%>^{�Y��~�m7v$���BSS���@؇�_|��W�D^an��Xl�x��p�|-Lf�oZ����Ⱥ��K8��

q�ͳPqd7~��'x[Z�=;�+֝��z��9@ao��PN^�(ǘq���5>��ۡ�Kb���M�&7s�&�4���8�W��%k��EJ��h׳<j�@e�)�ґ5����>���?�A��u3H@^ �ıO��� ��U�}���d�������o�7Ϡ"TL��mj�l	V!$�Ouċ���Fİ�]����v9qۼ��������g����Pˇ[ �..��rq�������x{���A~n�t�l��ap�^���/E>u�t� %%;�h��y���=زy3:v�{�K�a��rpZL(���]?I�)����{�C��C�o�`,Z�&t�xY�r�F e��9]�z�pU���٨d�QN��?��gS�B��&6�<�Y�*R ���l�k(٬��hd������/���l�(%���ىS�/@�g�s$8ƀ��]$͠�hE��a~G2J��H3����,����p$q��7���=����ؽ3/z+Wm���b�<�� ��x#F��W�ů�~G�ň��m�p���49ѯO?��^_$/��%E�a�L|���x�r�t�oH-�Oz<,f�����[oJ���_�K�d��~�����{�e{�O�_e� !���@_X��c��/L�f0(��f��Z�E�c�7C��� � ���у�I�󁶂e$�>M�y(����:K�F�E�AFK$�d���������f�#�=,����>[R&�a�D�1�=%�
�_� �K��Q��j�Ι�$�
�r�X��뒩��K/�d��lF��#q��ⷭ{���aѪ0�G'̹a
��
>�t�lZ��s��F!ב�ņ�gϞ(*.y7GD_3S��W^C���ԓ�Ez������vJ1ٵ{'�7R��C�+0e��i����b�'8y�,�Y�ӿ�o奼�E$�EE�a��a5�A?�f��b􁻥�uu���I�d{o�B�L�$��ͻx� �]� 0�>g���$�B>4�'&	q��������{Y�~�����(�m��;%�IT";�QA�6��C�7��f�/���w�Aa�������w�(����s��A�S���:|�bN�8-۵��ń�e�w�|lۼ}��kVf:����Ç������ȣ��H�!9ee�r����
t��������CQb�=[%���������n�v���(*툹>��������be'�|^����C�!/В�"���e��6�,�1�"�GRJ��Y4:��V�(Q�rDǘ�<�΄�ˉ��t[��M�?�X����1���x3I"����8\q���2�ˠ�����/���s��f��Bj�����n��P�    IDAT7πI§+?@n�4̘6Y۶ᆙ3ѧ_/D��1���xg��0�ֿ'fM�G�~��=F�#[�Ң�Rԝ<~�}��Ɠ�?�-?�$��A�f�9|MMn����c�����������A��#���|~��z>�h��Y�M���^^���@fg��٭�Q�n)@����"�o���(nW�7�\�&���'�Ii��Jϖ0ƶ��tU��+�h�s9�jF�Xd���%�@�i� �e���s,f�H���YZF-��2�Ԃ���xu��-���&P �:��1�5���\s�v-�x�fD�MpV� ;+��_�˯��̬6�X��;��cz�o�kV�ǧk֠�С����X��'�-w���5c��gi&�O��F��ӞA���3�`�Yнkgɭ[��{h������Qˬ��F44��m�W୷^e��r�;5��b����O���aKH�K����Q���	�%��K�D
�E�1��&�&���Gaê���%w!
@�%�A�?�1*h�N�p1�B�wM���(o�U�p�A���
�5`4��K���A`���b�Uc����%��dh�QQ�Q�2F��=��e�)xp�X4�	4�n�cӖ-����0x�p�7o�k9N��AJJ:F�)�ܕ+V���I��)�u�5h�<%��n�;��ٷ���(/? C]�Y��(�����"���j�kh����-��йS)>Z�'N�����1t�@�5:q���p��!���*<�ģ��{+��w��$�C�� ]k6U��� ��W�C�����C�Xw9p���T��]�8�J�@zflV�>�H�	P1[�@+Ec�(-�\��>��L�Jo6�0Q��͠�I4�6��s�Q��q&T$L��Q%:Ag3����rD_T.T_�A^N��j|�i+�&M������mp�"���)��8��ğO���NkB�@^�S��Fͩsx��w����l{����Ξ�I�Cnf:F�����:sgϝK���!5H$Jr;����������@K�3fLGNA
V}�K?x�:w��o�Ng����EMm�P�	J��/�&!�Ϟĩ}{��~���`���ױ�B��p�*Ϟ��Z�0t�u��L:)p����ǡ5k=yBl�%)���!	��&[w*3	�j%!��`�����L�Q�AVY���^��6<��o9�
;B�a1�(�N���F�A��D�GϠm�ѐJ'>��A?�����Q!`��V�?���:����{@&���	��p@6�3��=C�u�[�^���Č[n��lüG���w߃��\<��"Y�3(�C�,<p����Z��`>�w@ۂ�hnrA�1�sI)��/֯��oǔiSE�AZ#��̻#La�G�ѩ[w�v�-�+?w��\�9yHNKCA�|��o���g6j4z���/��P����+�t��$�`3<u��5;�S�� 0 ��T#�NI�J�=�N�L�b ��9�~��[�Ն�vEpzh��&j�ٖ �U}S�_�(�PN�������4$�`�	�[	��[7�a�����T�Q��h3��;o���bÚ�(��w�z֬Y�6I��y����N���S�����ɹs�0���� o�6)M;�,2�Rp�������j�J���8j��,
d��7�l�^|�Ei�N�8��)<(ϲY�عk7֮]��������}ɻK����r~����p�d��Lf8�49E*�F��'a	�N��r�Ή�D0[�@�X�G�̐�4��[É7��:�ȅ#�&&!���e�Ֆ��ŝ���p����=1�1����0�'Bo�����0	D��	dޣ�A�M��x�jp��ףKQ&6|��x7��c�{���dDi�.�4e*�3��p����ͷH��ѯ[)�3o��.֬Z���H6���&yƯ��`Єς�����Di$8haq���7ѩSw���U!�>r �zvB~~�|_�8_U��V��g�D��q�w`��Wp��Q8�RI�g�SQ>���ps�����|��x��ra��6��j�;�6,^������3ʅ� �]ŧ��?�Vl:6zX̫�	NO�7@��*sJ*���䙳0��h�"��}P<Mm�j�
���f�"�qb���R����Az��Xy�{#���Ł�G�氊��k`�$`ؐa��.���o,�
�u
���HF���������0k���f˥Y~��������b<���8z�&�C��M���3���!#=�Ϝ��A��Wq����)q�\75Ł�����˰��!�<w=� ��~ٺ]������>�E���pq^\j�[��5r(>]�G��!��h�!�Z��ht1&��6�S����8,c�B�����3+^3e��ȉ�n&3Zx�j�$GGJ�N��G,�_�&2r;�`π'�?¹9m�2S#b�a5CԽҼ�Uax�.��[�ǰ>Y���"+À�Ǫ��c����th��5Qܩ��q.\j�[ﾏx�	zu��k�����/?��w܁��Jd�|���:y]�J0�ʱ�w��᧟��H��Krm�שg�uH��=zt��Kބ�Ռ�5U��m#Y�f�7n������ō��݆)S��C�Z�%%Uh��r"��pU-��O�0mr2���P]u:��YE1����d���K��Py���]�i�1�� ����sQ|�,Rc$g�Q���2�9V؆�qp"���"<���qk^_�	�3;�lK��pԇ@��x���kk��i�c�L��)���*����u�����7` f�06���B��p�ܛ�������1d�0\;q$V�����6�^3�J��ߎDK<|�~=~۶m����%Ř0~4�._ƢE/�TϞ�,u
0RS��<��� ���%�R�TVV�aW�
,|�u����+-�{�(g��M������BE~BB���k"H����I�B�V�辽p75��铸XU%C4Y��k�7 ��@(���P!�mKk�#=�1S
iB/�5�R�HK(�!��Bb�f!�r3Xֿ?V}��^�l`��Xe�C�;-RZuo��a�2صA_#쁆�:��d�|'�{�a�'[�}�df���)�����5[$����6�v�3{2�q۬�ұ��_l���x�J9���ҹ��d�;�Do�9��S��%��[�0
�#���_o���G0z�X���=������ޅC��1n�ux�'��ݏ��+��$�'��W��%�*VWm��L����cF����47I4α�q�|\�&�	�p�x�dQEx=^�$�����5��AG���V٢B�f��G���������H|2Lm�Цk85��p@�B�� $:G��v֪S�s���jq��Id��I�HUe���ѽ_?n;���F��V���D~I��_g�Pq���`�ơ0=	c�����Y�|	:�Y�ϿlEcc3�����Y�ee���G�T�B@`�$��H�HE��,N�9}�s>y�H�'M��]��m�>���Ϣ�n�D�vy��u8~�
zS�(Q�|�Q����<�3��e�^�/�n����3�p>�674*lQ�P�k�57�P>Ɣ���rx�Ƅ��PQ�q�b��΋�qp���zB��i�3Xј��s ����O�س*1^�P���i) E�)'o�]e�	���3�b��eģѰ�a�l�(W� 3�H�
ȔA�������lm���T�MZȭ�!'B�	B�#.�&�Ơ^e�a�XԜ?	�*�1	_m��l���O��˯/�)>��鉘�����X8�1!dg��rl�I�ڱ��tú�>�/����&MB��Q�r�/\�Is}]=��b=�
���;�D��e�aBIbr2���_��V�Ben�uJ:u��������l��5�𿛠�׉��-���f�/���)�)����$_K/Ŏ�A����B"�����?]��6�j�f+
�K�����Ńx{�xy����rc���y��@���cP�̘��"�	0���َ,p�#�*�1��b����4!ѪǼ�o���ǉc�MV/��޿���މ^��cĨ1��<�-���s5�0������� ł��¬�ᦛn�SS��+`��W���}�/֭��/P�$Yi��/߾}<��<�s��w%=E�p�l��2�&�������F����a�t�����ڂц�b(#���b5K��xc�Or���������Ge�D�؊�I�^���H\�A$�TY����&��9��mK�Eq��	$�$�Go�C?#��)��m�@� ���韣܀��0�o�������>�Z\9�#N�U��E98s��}�e8]N��"��s���~�]��` C{u�}�NĂ�^Ʀ_c��E|��	TVUɅ��Fʤ��ߥJ���,��*++�����ѩ�3.X �#Юm>��S���&����:}�`�G���|�=��n�.���(�`�X�<��4�e�{�kY)��	�j/>l��y�-��|��2A崗��k��H ���4�t�Ђ�\4eS���F9_�A��p�p��4�m�ʋU�Z�x��y�y۟X��k��!a��U�)�����͠U��9�*���Q��=z������J��N���
<����f��=w�l��z{�@���~�0�ʞ����'�?��w~�����K2-������n�z�>}Z
27�f����h(�	���	W����u���?�QÇ`���P�~�p�py=>~<�]��?�"6|�`�9�����=^��WF��o�@L�:��Y��|/�:�JvdzF&,6;�4�2c� �-��S� MɛU�����*ަ�M<�䘝��J"[��Z������خ�zbܕq��	O>��sJ����E�(���y�PE��u�T1����FMW=fL�����#������H�zv뉏>Z��vmp˜����;�l�Jded�_�Θq�,^�;~ق���h4?��� -�q�c1v�h,~m1�TT��7Iqh����������[n����ŗ_}!�s�G��5W_��{�1s�,يϾ�F�1g6��1��q#�<S��M�
Ȍ��F��9w���Cصs'��������,!�&��A��E*�&��aąC���@�s��G$*[��R3p8�&W���R<��!w���س'��p~��V}�=4���v�[��i	�
��GPT��+��Ş�P�kfL��-n����ڭ�M���j���
��.�{�m�-HBum�F?Q��_lK�^��׎E�v)�e��HKJ��qc���_���}0%%���S'OBVF:v��#�WBΌ�	�)�n��b�����C��w�nJ�c�u�Ѯ����1R�3���o�����6G�-������	Ŕ8��������کL̕�������2��Ua*���*�+n����0$�G!'.�7�=��@Kr�D��kG�GlԖD�������u��� ��.�7K�q1�Hϰ��9����8���Կ���9.Ǭ�L������/�ϣxK~ߺ��jd�l���_-��F��+BYql��{T:$��v���b�`$��8{��jke��w�W<�����ӄ�]]S)�F�*48�P\\��&]'���V���#��3���g_a�kK��O��$40�*���]� gc��~��B�f���3'���_B�Ԟ�&6>�HBec�H�o�5
�:n���Iv&%�!e�MY���$�(�o�ө����Ҙ���!�����ה$9��Vp�ǅ�gh�[%<^�h�%sQg��`M����:�/�[mc3Z�!�;l��p5�#!1��/]�A�ń�dF�)���y��כ�7ė}�\%|>�Щ���͕g����ΜE�%%'��f�/��)HI�Bc6
ą��AO+��)i0�P�Ԉ��i']��b�ڭ���qF;\>��*%-�GK}�Ϝ��Rta�jT!�4Q�H�^$,@�I��nHKM�0��^o@6��NWL���GJF0%���K#O�5}��P5��hqCe� g4&������ jN�W�F�w� 8[w�J��?�`,��T��j�{�4
@FG+X ��1�G*� �--A��b<U�S
g1�?%�rL�C��ߏ������K���(�4A�j��h���:�n�:�CF�	�x<9�u	��s��H��������F���$����f�Z����>r2��q�\��!3=}zu���~���nH(G�����!�H��_P�iS���}�*/�ԩS�{�ٯ�s��ݷ��瞃-ނ{y��:��'���c�tC*l'�F��	��!D�	�Vɴ���B�I���R�^'�%8|�9�&x^0����5������iWq�l�]�oMDǲ�rh���I0sbz:�];�j�xe�;r$$�Fb��l���LHq(������j��n�so�V݂���ѻ{9to���u��S��?l��!+� ��>?��(�q:
�l�5y
�2q��������7TV�GA^F��?v������c$�j��_�Dy��1r�\HĮ79�����7̂���/b�gk�W�O?���Mx�{bN)/)�1,sy�1��WX|��	�6�'HNId�w%S��"�
��kJq�\i.��	�(A�f����'\R�E�����DG�ȃ��.xal*�	� �=�� �XzH ��p��:�:���GQv"6~�	�'��?�sϿ���"�?k׭��h��w��]���50 ������)����pp�A<��������/p��R$�#F�@����Ï?Y���Yh�����^���Ǉܬ\̞9S$m����2��_y�8�y�`�G)���1c��������o�J +��_�1����nE�]�v��OQW]�������$S�L�=4�K���F3�*��[x�*�UN���b�|D�>���� �b��p��AE�iTkj:����Ҏ�Է��R�V}�Ĵ<x�E�	~,VB�آ�Q��r3J9����I&��;t _�[�Y3���S��ـ���P���fΐL�ի�Ñ���ַ3&��'�>�X��8}�^{�-��f�-)F�~��h�3g���G��N��jj�,�u�#(mۺu+W��Q#p��{Pu� dX�O�>����k׮|�hQ�9�%"��rLq:zn�i֭]���O�K
���=I�6��C/-���4]n��H.�X^�������ļ:Ҧ���&Wȇ��ě`OIL��B�~�1}�dgرn����s$g�&�(� bM\���݄i%Z�`f��C��-7�
4�^���bȄј5�jl��gT�� ���N	��b���X��+)��j5J�f���`���ġr,x�\�m�˖���3�бC�o�6V["��E�Ę	�o,�㫩�BB����;c>j�(̘1KfΘ!g��c����{�O�}C��!�b�L������vh�k����\�߿�W��%��/p���#Ji�A�P��=N���f���,L�DĶ���ISKO��O��@o0�l�@o�Ñ���vХ� <Z����59���� ;t˹`�����D�T�>'����Qrz
j�j^�_�>_���q��Ydf��}Q���5z��؋��&�d�#��5��G�̽�~�W�P|�i��ִz�оm!RS�e�H LeM-� ´$ؑ��!ߍ��(�4�O���Eu(Bi�RT���?����/��K�p���`Kd��^k�l|^�������p$��������g�ʹK?�x�Y[�<�{ǂ����
��C�`4V�)A�̙����fP��3M�ۤ[�T���'�]����`J���Z'��d��s`NUL����,�b,�PIN�:'�լ����x=qj��
	Z��:n�C�PK��elJM��룘3�J�[�[�MCzr2	�8{�.U׈�ޠ��5AWN��F���ؘ�=㰖T<��Vbo��f}l0�ğf6������K��x��װu�n����s��    IDAT���1W8�ߍx�O*P�/���=��OE�Ō�˗�쬗���6�lL��-�r.����$�c���r��&��7B<#cQ-�*H%�H�;����nFmC#�!5T�X:tE�Q�"��)�6
��/�gֵ��$��n�Nq��@�<A��Ò���Ghq:��zą}�,Vp��&$^�L����A�Y��^x'O���N��J"�4{��K�'�rZ�Y~�F������J��-:�m6�\�������h�����g 1͂�mEU�{*��'�Ƶ8�s6 �v���i4�u ƨڿ�0
T8��O�C���*Ų��"7/_ȵl�n=�Uk�\�y������E���y��i����r�q[~��{���b�%������z�۠���l�3P2��g3�����QJ]�e��(�:�d�R�=�S#l���Wβ���fxHNE����?��VH��'�B�4�����J%���E����޻!�aǸ�#��Gp��)�p�Tj����Oy�J��m��؜i���u��}��HJ���?���"_~`��A��=�X]#�z�HYР+�~
I�4D"����c�����!d�`��W�T��^)�<�n�{��'�CJ�����l��)�[Kz(iE|��+^�`s:��J����Nc�*L?%h9���Vhl4�r��A|R2s� �rH��
������@��=��pFXm������vǪO�@8��#9>/W�J���������ɖި���	�5W��sgO����񣑕���?߀�}{��1�P{������ӯ����ը��'�S�DL�f: @���q�-�
Րp�%�(-.����@��ih��BB���8A�J8��d�y��(.76ȁ5x�p\{��عc'��L@�[�P.�[o�I6!,����*�4
�9�a�F.�����"Q^%�a�D�Ɛr^6�D �E������T(�������V#�`$���.M;'��D��6t����!���"���΃��������ق-?���{��Q6g�?�'�|U=n'Ba?�2S�>/jo6}�-��;��k��`�Q�8�9�̈́ݮ�l�C��凟q��
Fx1�wG�s�D,~a!~�a;n�qZZ�Y�ϳ����J`�Z������2eVb/�F#|n��$Ǯ��q��]��|�͆��_1k׮�͐#��K���ӯ`����@H�,D��`%S�)Ivt(,���?%���^-�>1}-�� ��|?yօd���S9	�����=7��Ŧ>��53̶Dd�C���x;z�QcF#���_Uغc�W7!g4f��2`�-��U���Q����<�*.ȅ�ی��nAZj&\5g�7`��r)�-v+l���_�X-E��y	�w��+{a���v�1R�c{DP�Gaq�)1���hgN��_'O��r���g{Fj*�w�"[���p�B�����-�ҵ
�,�y�F������S�>�g������dٶR��9�R�ssc�"+;y��h��F��r�=n��j$�^l��စY�l(��IV)a1GP�I,,9���\6�а�T˻É9�1u���48R3�pd�Ciwd�u���=s�a���Q�䰼�j�;Y4E���ݼ�(���"���������y������d5�}��������+Ͽ�_؈1#����W�<��E0��j�M!�;�?g��yҌHIM�����GH���"�j��d����%\���q�'��[o�������*DTm�����/�Q�q�;�vB�n@�A'����Y���Dx�킯g�� yR�X{iQ]]%Sz�/ E�WJ�)4b����&�yGD�V��",*ȅ1tv;rKJaNɀʘ���0t�4]p�j�Y��:cyu���\�3��L���py\R##�[EI�'�$S�8�����6ƛ��m4�`���U}7\?�ڥ�����٣������K�d�	����g�:�ۧҊ�+JD-=���Ա�iAD2Q��(�*\0�w#���Є��m��+��{� �|4!*
�H��m$!�x%}.��#a� ������0]lh�f��s��x~3o���S��iY@���8��w��  J��/*;Lf+�.\��,?�119�{�5�,lH�,'9\#�F�Ne +w%�M~�i�m#U( }�MZ@�;�%��� BN(��?�C6�V}�'\��O�� N���&u-�p�A�����Y�ɞ$�P%��f�?Cq��cK|���n�҄Riz;}A?����[Э� �������]X���HL�@��D幒����
�`�/T���-5�S�������%uS @0�;H�wڕ���@��H,ҡ�0���K�6��!?N��,C�{
��s������W����R�n��ئ-�FN�93�pL����0k��Bæ��*�_��;�"�Ml����p�@�&�I��ϐ۽p�~�(�� r�~L?��\����8u�l�Bb�����R��K_���*�>_��U^̌�-������v �dJ��������Ż�p*J���=)={�FU����5-��������*��*��i�����cpD����Rd��o�q��]AZ8?�!C�@�¶���x���g9��c/�NR�U2����)#=�����w�u���L��?ƑSg���8p�$4�T�s�3!!3���*�X��t+@F8"��C����=�_��TQ�&�:�9�-�4�Zh6�'$�?D����J"������j�'�E-(�%1)ul3�l�6%�Ë�ms��hy�I�EYǮPÀښj���I�_[�Du�%��*��C7O¶���%�c�+�jP�����`[Y�V�l@�s��B����� �O��A���^��q��ii�$�1A���Ĝ�����b�ٹkw<��BT^���T����S/�L~�Ф��i)� �U)H��FJC���
)���W����.�[�!���#f�h��o�ʤ�fbR*�z3��z�Mv�P��qZx������j�硣��{��+t��*���洒&񈚲).И��K��ˇ������2RHIN�ub��&��ރ��<z�M�v�p�I0��ćv��Ξ=/�B�#	��D����f�����)��fR�M�)�`�oUu�@A�����G�Ҏp9]�s�>X����Bk6��ɢ"#���Ai�5q*X@�=�4)'���F8p�,!lNd�DRT�45����&)&�V�Q�r�-F,	I"��Ho�%9��r�\njFN���''#j�"D$~�Z�ldv�:���� 
����0\]��|FX���k�S!�n�%���Λ\��Fjr�lB}����<ȭ&-ܗ/��<u�l,{�]���uF0��ʋR�[��&���@��fl�uz��@>�0,���U��p�O��S�R�U�󬭩BS�}�CO/�+o�-?���
����^�$�R
�]�}�����$I��)��E��*�~�-$����"[0�<������������B���;� n8D=��Zg�KԞ���v�����Y�s�
��
�-��Dx��k������c�D*�Z���4�� � !�"g"/��r=��4���v�0�Z�1��ô�a��x�g����DL�^��+�����<�<�����)Í6��TS��)3��ae�U���Fi������Da0�K>�����c��SO��w?��~�#-3�0�J�(/�a��G�S���$N�����S>Li1�+^�&�I� p���E��)5�����t%2\dD��@j�H���3�M$ݢ���MkMEA�N(��W�+N_D�hABf.|q:I�Sk��`�,{F��(��3�T�q^���&�>���l��ɤl�O�B��K\�OJ3x˔����%X��k�X�r�����1G8쓌W���wG��&��@��l�=Pi��j�Ƭȉ�>X&���vn�c�{�_8}�����̸T��!!]�Ce�૿ߙ
��-���$"?��*XLf)lx��"���M4���S!���ReKH�Z�CQ�)�ge�Э�r̔w��������^�LhIMGR�|����5�`O���;D`�7�����7�@��
E�y,����@n[���ƀ��Qdz���DO����
z`6㺱Q����y{v��d B�ņP(���z�X,&��!�0"����.~HiP�Z$ۉ��y%�~�lH�/��ܖ�*�rvnn��hlIx�����`�������nA$������_�e��1'6l��j�|M�E��X��9���BAA�4q`��H��͛7Ŕ1�H,{�>�X�Z��Ά��g��&h4&���C�`�61����{��g�"I]R^J�����F�(bL^�w�dY�1u��j$�U�����c���D��돒L5��y/N)��n�s�V�X	�"`��L��o��߷����K����b1cܘ��Z�W�[j���.�l��^��h�%�+!%m
�j����NX������p�݊8$�.��Y��N�DͩcP�]��NCVz\-��k������\=v
��K��v�ETk��>��^�эp���!-+[T$��a�ȑ"���Rf[~؆�뿂֞[NT���,�
�#.z���2+�&7L�:�|��T�+���?Mdl���ϣX�y�{���hfu�V��[��841�!�X�36�B���lIF=��E�K9_��O;v�������SI����PLe���@1�(��)���<ӄ�����b���ZG�M8~�U򡥡��Z$�|0}�EC��En�:��2����c��"+3S�]�'��;w���`��=R#�CL�;���6�X��2T�?��/-D^N�(�B.4�`ï?��?��ƫBJ���wd�=�e�*����&@�F�A�uT	���1(�FE��F�[~�&�γ�L�v6��^��aW���c�E)z����7x�?��7�X\�?��?��/��7)�8�t5��d���Q����mFxC~DHQ$��y��g♹3�ㆵX��HHJD ���h�@F�Q��,8ҿ÷������r���?��2���|��iZ�Ղ�J�0m��~�_���e'��Fy�m���J�`��wm5®�5qS`��'�Q�~�B���p��4�*E]1�a���Iu��	*�P��a0[`�LԒ���.p��ˏ�gw�˟�&��`�(��V/bl�����%�o�B��ɠnP)}���Xn��>��Zd�HI�.�����՘?�.$["�1q
j+�"19Y��8-��
�?�gaHM<'�!��S���%�7C�L���p:�C�h�)�d��f� ���6x�g�{[��/�`�@��	^��N����
���k����*���~~��(fm�2�0[9�ŭ�΋�FM>[ԕ+�V���!<��M�t0��,�_N���Ѿ�յ8t�8l��&%#��CH��;�M�	6{� ��Q�Ӱ���Z�R��Qep6��xa�R�Ʃl���쒳��6K��n"��D�@�ٯ��8�.^��o��5Q�����Z)
:�a�gVn��	%X',c�yh�������d2�# ��a��]�<�����O;H�:Pt�S�zb�n�Mp^�FKc�"u`�%Pl�#!)v(ѥG�Ŗl��aN���KJ��I3$�Nǀ�8-���ٔ��دe{�	E`�&�]�2=uV"	�9�9���Z�3�"*����ô�|A��#�IYV��U&�hYx�G���ln�����tڈ����fTo\5�>|�|��'tz�P�P�T���Ms�dS�F�`����e՗���fTG©I/�\Km��Q�vM��MR qHֵG,z���l#���w��"yfө�!?���,^VuЍ�s'ᬽ ���QP&�lY��O�' 5-M�2G$MY�ѣG廠o��w���|��<nI���Ȁ����P���h�0��S-�Y�1|�d��48YYKJ6|qz�����QJ:�
:ʯ8 e�#E�R�(�N��(�~�ىy0�$r�!��` ����^'��Έ������Û/�(&�lU���K+'�.o3�ڈL�[�;z
�&���s�3�!//��̹=e�n��/LF�L��@��ĩ�нoo,xi9�:U����!M0e�����Ol�0h����:k��iE:G�5�t	v�(i�?��N��:�j������}_���͋l�0��C @���LB�d���LH2L�$@���+`c��elK��$˒%kW����־Wݪ�5|�Vc�7�������d�]]]���?�|����C(�?  K����/_���d�Ĕ���	�1�f�7�G3��F9��p��a��E��ju��G�o:�7�bqC5��g��+����Mn�F顯�� H}]�Ii�9�3�C�<ku�����N���Y�ɲF}����=�l��7�`jf��]�n0��_�Δaw���q9��/����,t\v���ߎ[nޅ���F*�FJF43�|�$k<��*�i͑&���5|�;�@gtJ�P����Y�2tJQ���:���\�X!��&�Qj��"����׉��83�����+��]}.���~��|測�=y��7a���⩠�4[`�����^Ŀ>�8��VXmhZWs*F'T�*}	�4�P��:�p'�<J5e���n��!��s�H�5&=�M�萩�1ZC��:��A������k�[P.)��ٜ� ����B4�����G4zU�����m{vA��HJ�Wdf������e8��TU$x1����gpm&�َRR��D������7�a,�p��.��E�c��MX;:��gN����<��y�s�|��>�ps3�M^�����va~n_���177'R.�u&�,�"-mp9ݸ���p���P.�p�`�:��#O�K_�<m��ۼ��^T��`FYo�����2Ih5����<�'�&wMn N��4s����:J՚�1<۬��cP0��C�� g��nD��&���aV��Ku��k@�V�l,�����"V]�Á��&�a�)�e.��FXo՚d�tSz���(�X�+HV�0�|(�yU�W`60��R>-��j2�R�.���b��L�BV<@��X^�۷m�o~�3��J�>V�<��><��G%f�l5��;��W���F�W���c����=���b9�B��́�B/>�C'�K�0F�He��6pQ�B��薚�芃	�e��2J�%!\.3g��j��a�hq���"�T�5K47���I�ݚ���@ȭ���w��r�����Pk����M"�u��I�B�C��hE��s��;�(�L�����~�^~���/"[Ƞ�#�.7m�X�Á�*�ʹ:�He2(gs0;�o���']�ͪI�Wn7\./
��XHӉ���6��}��00�_�οa>���΂���6DT�@%Ei~�L
f����h1��ch&��zw:x�A,,/���+o�rI4X:��R����r{awz�+hB}�F��.��Me���`��o��r'�xzO�`|�]0y��2>�dGM������+�:U̍e�M����Ps�{���.K6��ޙ��Kj)+N�tv�&�`�)������<���~	c�NI+��R(J@6Gr���C��Up��4L��T��*Bᐘ�(JQ\I��he��
"ඹP���=���;�_qab	��I>���њt�	�\V��4����N�"�X@::�Z)/('��ߏ&f�5"A�vtu᭓'K�5N�hYTh�@�u]��_h?H��Ϡ�i4D����m)W��Ӌ���!�U05��ۇ`K�8>��BJ��rU:nc5c%��g��I�P�y��,�J����fRp�}��%��Z�F^�"4���].fQ�.����w>�_x	?|��p{}�I�A�X��-(���E��y�p��������I���	��t���A�� L�LH�!E�������}�-�a�{��y
�N^D�9��.�'    IDATR %�i�9D-/A_-ʵ��OJ�-�;u1�����FKSX�Yj�XLI�{���%��*���U57=�'����E[un�"�
�:�:yZr�B-m�v�{?�	��
B�nX�MHfj�譀�)��Om���Ȼѿ
����}�D�ݶ ��j��7r�x�u�kͪ�d�D��qˍ���߇��$&��e N��0���xm�$��5�b�_�O�}^�Z�$lO7޷�z�t�¤�#�L�V�"i�3��KF&͓
%������z?~း�Ic�;!k����W�
��
�yT�qy�ܴ'z[.Kx��{�����D9.�lV�Z����ǅ3g��D��Jt�~lj��q�&D�â�d�(sj�}�y��4��!�2e,L/�ix½���̰�è��\����0Hv"���>{u+��k�B��%�����#�2r�eǩ��臘Q��P)��k�����^��������DU�\WyPE ���K��$~�{x��	�t&��55�����p�He��lE29�����oҤ�Y�6jj.��~�L�d����M�jj
��IsTJ����喐�|�̒П|>�PF[�Bhj
��q�={��Co2����Bww/b���O�G��+��r��i@SK�p6lي;�S�W�5��R����9�2%
�8r:_���ێ�Ï�jF��Q.z:1��Fd���{R�[صjg�� t��/�n��&��6�(��:Y#E�Il^݅����5�t`"rt�f>��rN(���9�g^����T9�vl\3����Q��Q���ٴ yi`��a�l���	Mo��<L��/,.~6��a�sK�竘A�n���%̏��^W��nD/s ��3�z��8��>�|�MB��򀌉ݻ��駟��?���1�5:Y��u�}
��������fSt�T�,����=�?�ӿ�-�Ws��#p6�!�V��������.���bQ�twV���Z"��L�#��l� `�b���d��>�gZ]�f��N6��*�6��t!6-��)�v5���u��3�)V*�vZ��h-*?+��E���@�B8�N#W*��;c�jzj\.q��'@@��R ~��b��b��9����G?�ÄG~ �.��'n�6m�G����g.]�b��]�Ƣ��7�!���k�������b&�PS����aÆ��Ɨ�pXܲH~�����3?E��(�6oG��HЇ�RG���&+ʬ���@D]P�w���Pvd���$O+H/QzD��:iR�W�ۢ�X�i��I����f�#z���T�F�9EE�h����~�Y|(�S(%�022�Aae\�v͑��������׶�Q����[��\r����R� V����	��Q\���l��f�Eyn����u��2���͞�9�^_f�3x�'ψ��g��w�C��O�����mC$Ҋx2#���vl�s����z��h_�M��2�h�t��k:�ג�����x��������R(��5��ݪ-����!+Ƞ���I��9�����K�ڍ�����ڦG3%Y!�
Q����
��C8	[W)�����f��X5�]2�E	|��9�q	�{C����4Μ~e"5jE@��hͰ����0�뭨x�W��BT�`�@?n�s#��B�t�"�m�Z��V�A)��KO���d�:����B"���aPo-Q?�b���s@&uy:�ѥ���c����M� �����[#B���ګ87vQ�IJE����BH�
5N&��������f���+�nO��	A&��g��0Hj��Ǚ�Ǡ�8aij����@3����:چ�i�GL�r���o���#.��&�%:'tRne��Fkf�D&����R>�������ع�/"�8/���u�H�U��a�(���&�/O��~JU�[t�<��}7�=�������E1y�H�R(�p�\R��`�ZZ1�y^>t���PA#j��i����<i6�k�KI��`T+"foooŪ�!��D���3�����{�����U���T�}T���܂=7� ��-�`�\AW?HG|�G?����h�,&��8w�*
�
��Z:{�k�D���)[Q��e��L~��� �r��c�uPkX���
Be �B(����a�(<'M�׺R�^�`�`���;��6SN)�\�P�R�&>��>�n'Lŉ�W��<�ӧN����:�;�W���8��#7��)�.�*�!���NW���������9�t��2��:Nj0�.(y�+Y��s�M_�N���~��	�P�_��#���Mki��'.��bQ=�4��0Jd�`6���7�|�:�E�R/W1�? �ۋ}?{[��D�������<�BE�H�(<�dꃼb|�{�"���hy�ӡE�����/��`��'�0�@�s�o"M�{p:2���޺�¦�|��=9�P��!��,h�2<1��~U'�ՙI|��bl�
�[܎���7>�a4��(Tx�zTK�����(*5X�l|5C+����oN`߁#8z�� ��|�D��3��y%�z>�|l��4*�E8�f��
#��κu�Q�x�8w�H�;Z1�a����{LiԲFs���z]L���݋�o��@ �LV�{\|�����t	��(U=����7���������Fh�,�9j�>�X]�kD��5j���@�B�%�vX
Ä�{�^�5����DȫE4�����}{g[X���y�-C~�+�s���e���EW�� �ʣ)�����v��x�\>Ԑ��9y�E+E��h	7IF��r����Ұ�"0Z�H�i�A}3�^4�@��X�E�Ͽ�c���
���#C��u�c�m��*��J�>��:�<�����[\PI�6u!M�����o����o��,�EA�9`U�58=A�?x<�T���v���;�"^.W�2�> sA�@��7�1��_���_���r�׈��\,p�A\3�1���G�EEA%��߮G�k@���e�D;��,I��uD�3����]���ְ8rY��Z�!�I	M�.�ٷXlf�?�xZ�#�s����o�zW����ʒO�ײ�ey�6=b�c�?�������G1�7,�Ձ��z߽®�;��'f��h��}�w_���5�j�����7o�����?�#�Z�
�3S�h��yÆM�py��_d�g� �Vo�7҃l ��q0�F�(���#qFhI�Z�]��P��i��k���M�C%��p�I�è�TI��d�6p�YGE�i�	4P�*UWoD��J=s����rjgY{�R�xT��x�I�%��*(�2�����"�́Q5��:ԡ�M"��:�*
̪� 5��<�Ͼ����Xq���H��q��ttF��J��Ãk��\�"�ˈF��ꉩ)YD��V\�zU���{o���8y���0�1�D����f6�m��j����"Zz��@���HW�(��3���k�g��̨���;���7��_V>�o�g��$�@�,L>^�j9����%1���dQ��m�¨7��Y��
���t���t�8��٠�ҨVQN%�K�tՌZp(����U�2Z���GP1X$��lv�t�f�Q�M]��P�y��(ԅI�f��V��k5�XS�jh ]2D��	��a�}3+��RR��F�M�P��������z�Z���]!�\����m�M�����m}h��,R�k�)�2���Ҙ�Is�'үE�㍶D�@Of�_cdOFw�_f'|����1K�1�Eef��5>���^P�@>�+��ނv-�Mc0��K�3_���"4TR��G�*� �Մ"���C���g���m��B*dS�,66��<"-�-H�#^��b1!���ş����gN�(wdd7��]t,�^%�)J�?�4�UՈ�Rǹ�	<���4�`�<!m�j�� �t����"��z!'�E$���]��pXrnҹ,GF�f�F<����_-^��"�R#��V*����cx�j9�(AO�響&��墵��>o�����g��h�퇳�U��
�t`k�]rs!M�\g͐>GD���q)�1H�m%u.��(��� �zT׫��T��0�սx��zPGĭ$�F|}�hp+M��nQt!�`jz���TK:�ـ�5��e�:�\ZCLĕ��V�f=ʢ4s����e\[����	�>wQ~^n)��JsNT���bV�AR(&QNGaթh�q�m�������SBɠ)ώ]��䏞£�>*�!5��tF�IY8i1<Џ�?�a��:��ڻ{���k?G[j[#���"x�琈a�"��_{'2,�t/�s�^��`��
�$SF�29�,��Y�*�x�q.k��4��]�$�YE��%�HE�ʣ�'
X�ӂH�G<���Rh�S���b;Nǿt��1����1�Q�JaV�E���R-$��w#V8|��s��N��Kc>��t"�|݌Q�JE޳����9)q�$2�I9PH��L�hmA��	�]�ر}�h�ƯL�k���<U��%������B�.Ui�z���������x
Ãð;]���7���d��o��Èe�^��p�U3�T�UK�1��.Q\�}��H[�hϚ85y�y�����:�h�p��}΢i+�٢�R(�eXuit�Е�(f��f:�n��MEKuʓҙ���Pw�RU4�"z�e�N�`3�آlF��_�����Φ%���ўP3Ju3���#\�&����I����h�N��Bzq����%8-:�u�崉>���M{��j�czzZ���� �[�����œO<]�Խ�!��H۷��Ν;��gs�0�"����"��8�[��j������0�"o@��en��`�!�6��I�L���o8E�k�I2�ؤ�{���n��ED^��fQ.&d��vrc^DQ��X�&��UjE��.،vD��7w�a��g��g��
��l�+n�\N��V��Tv�
�߃LQ�b<�r�
��:k Jŀ�uR���U�)*Ȳ(B�]D��a �$��KK��Hţ�ǻ������Y�v�y.,.㡇�����ͩU��^�۲E��R������4*�5��(
0��X�aN������/� ,�6�m�
{�U�%�:uU��f�����S7ؠ�I�=Z��;�Ⴆ�'��&٘�����Ia3��2����G9j3N�ǹ?�����-F�w3�������zU�FB��H%e���,�W�]Q�ř̈ƒb�B��<[?l�*�EL4ʪ�]C�+XT:7��5Ր�����'�ӕa5T�e��Y���Y����+eKK����0������o?.�P4����P.h>�����G����q�}����[d84�X\Xƚ5kq������(���>X��ݹ��>�j:�$�@��w&���h�"�c��D��l�47F4�(�+�B,=z�8#����rr���2<�WМ:�9�q0���F�]��#������0#�V��I	�@�$�v1dG-��8Zm�6���-ny��fT�Y��4�M�O+��U490)%L�}�N�E-�+D!E_'n��=��4>����@Oo �^�_b=҅��O%���"y��;�l�ųgp��7q��6][s�\v/��c�X��������s��>���A�B6�u�U�1�@����n�VDe�cr^�y�0nߋ�1�h��5Ԫ�$�u���]W��P��TA16��ܤ��V�<�ƺ�]h�Y��3L^��2f055)K�ǅ��w�kH��I�V�|e@`�w^�%(e�xM/g��+�bu#K)���!�ղ,�l�jP���a�,���`{G�Q�&�02�an��Z4Ξ���g���8��h����B@�ܠ`dt��=ȥ�q��1�=��g����;�����8u-��Ƒ����vZۤ��B��<�H��4Id(����zȤ��+�12���� L�a0��0ȍ���������&*���ͅ�K���ސ�����z�`SDw?�alxE[D�P]�i�@�7��]�������d`1h���
��x�tBE"����H�����nm�"�k7�Y�bS�N�h6 ���&@�+@.�"�d1wAo������Z%��z�j��J�e(�j�>/>t���n���f������c�����F��/d��	=�EKE3�8o�]�!������q�9������|dUU�����#���!�F����v������.?��� �f������h����e"�F���k��B�3iA����J�
5d5�ݱ��*�6ȡ��k%o���a�Sll�\8j�hJ�F���#��
��"-��U�A�%�$�q�*<v�Rq���ʶ�J#S�����d�E�N,oDZ�g��!�JȧP�-@IDa�+hm	�����):���i�M!����؉�x��Qi���e�%��EoBo>��қ*���lw��0��k����G��7��=�,�s��_s���P����[6M���(:"�Rt�(`�p�I�ױ8r�V��)�3�x�Ă�TV���"�hR]��ě;
]f	�Bz��B	N�W�!�l܌r�a�ԕY,�M��.r(P��,R��.��ܬ��MpX�kj+)96M��0�F;J�@��B� 2��V���Bf��s���k1�0�׃�N.A��B�RѲ�
�#?��������عsR��"�Y𠳿���6��A�R��,�MX��q��A�7n��Ǐ�>�T`���Axt#|��(֭P�$��XW馪�j�ejȠ֜�bcA4�K\.P��'tq�UJ�r)��˃SW��^G�0�Zf�R
6��R��q�uir��~�\�Uu&�\^��m��a�׈F#�dL�1k� l���y�X�y���b���,���h�l�L��RE])�u���sא_��Q�5t��`��K8�x[ZZ����`3�-dQP
8�,��_j�(D���sZ�a�PW�ay��,/-cptru�|A�ȷ��0��:�� Z�7!��/�N��4�V�4�Z#�|D��䁫m��Kt�J���A��7�p�-vV�ֈ��9�1rq�q1FbG�\��]:�s���%3l6�M�ڜ����A�W2��Rt�Ϥ�-bn���%��Tp��u���.�J4�`S�!U��OE�Z֌��%�QDǏ�fPkw�K�K{kr�$�f5D��F��e���s���_�{������d�Rc�֩s�]�3�TȠV,�n��;ޏm;w��C'����A3>K���6�hA��:�;^q��Y�K$���1��44d����3��4i46m�o�=~�*��l
���Z@1:�噋H�f�D����L�#��J�.�D�km4�\�`��ā��\/���B
�R�#��0�cv��7����h���B	6�^�l^*д͊��Ҳ�k�-L�ʉ�CoP�s��fx�[�Rq�6�066&K���5�&�}ffZ�a9����70�O}�S8|�:zT�D�$��RA>���]׋��~�2���߄��C����ҍ,q��V W8�g^�Ct�_"�"Qш�ڒ���Nݼ^t&�a��OS�ȯ�g�!hS���ebp9̒H�|��s=d�Hِ���C��|��z��3R���C����A�B�@�T�YY65U�;�Kv�]����_�G4_��F�l$��(�;��t஖p��[?qv�1:܋B&&@Qw��*T����P���у�w���q�_�&(Y"�FGW�䁒2���47��ܜ�^�K�鼶��B[k�<���Ú��DS� ����Q��ZȞ��
�� ���U:� �f
���hESc��6�(�B�񊡔Cg���l_��U3���ނB��A4�ݲ�I���r�bR19�ġ�o�ț4%L�j2`��|��CBR��-���ҜL�����(Ø�e������By�#�󌽑���\��� �<����j	�\�������a��^~�%;~LrkI���������bH    IDAT����h��~�X(�j��)���V|��b����Y���p��9q���D�\���)���:,�f�����뗞��*�e�v[(��� �ӫ_i�B%:��D)��.i���B��i��h	�[��w�De�ll\t�w����QL3ޕ3�￈7�-�q�c�J
 9��lY�4���O{q��U65+�NA��l�7z��"\��Y��8��˨�c88 JBᰘ��7��$�-V�Lq�׸�ԏs�i��zp�VNg�A7.�y�n@�"'�� l�*UK�ԃ���qR@�������]D)������p޻�F����r0]�%7c��8�z���͸x�(����]kg��	m�����>�;��CtiA���Lz3WBX�v^�w S��Йlp����k z���f����1� � nXi� .^�5�SR I��\��kL�,)b4�Q>�T��Z�i���0�0��Q4I�K�<Y>4�$�(��	���;(bo����U6���jI���7cv����v�a�O�x�m�˃�� sr�2R96�f��L�k(Ѧr�l��9(�%��G���=7�EJ�V�n�K�(f�Q�����7�IvQ,B���7����5�S��1���6o��)���Mp{Bxn�k��MB�;�i@k�0l����u��ʦ�(1	܊�=���{q�&���rmX�}6Q�C*XI�����*��'��������@��C�V�S�--�iiM7--�͉jUGY�d+���"������֐���$���Ѵ�d��[�rM���A��@��F�dd�f;6�US=�<��<��>>���y��U 8@ǿW��!�w� �ɢ)��Q��
�S-d�9����̙��X�!@Uq���HaS{��p=�m�`�Y�\N`��hkk�Չitv�"���O?#�;�ى��:��Q3�P�r`a=b�ƻ�� .+O�Nh��v�����A��X�mb&�͆�B��.�!���YtK���Z��i��0��?�Jz6��dFLd�C�k�*.M�S��s{aq��3R#m՞5��D�LȑMM%�*N�d�iH��Hc��	ws;l��7�F�la9<�A�k�聮�D0��X�z�Ԓ�t�ctd@��\>�k׮ai9��+�3��G�eIw���B��y�8�1���*Aq�����p�i,�g?�۸�����4>���W�r^��Ad��auB����-�fL"͍��sj�į��iKM^�w����/��u>sԻ�<A)$`@J1�dl���&،A3y��l�,F�0�F��Z��PH3>��U�*ibv��́���]X�G������ز,2��t�A�d��AU���G�X�J�1?�L	��BKW�c��PⳢ�wua�P?�>�7��;��Q��[73�f�\n�?�d}
$����͊�oڋP�/��P,)��gS�%n���?�o>z
?��
5,�.t����j�#_aD�A��D;C�C#��0!��@�E#�*�������=�3��d i��ܝɂ��U
:f��E�m>��{t���$�Og$Ӭ�=�+����X�L���$�typ��E<���b��3���݋�?p;n�~=je���d�Q�`��X��au9`��3�qeE�3W�8���%��d�4P���AX-(���QX�����?���@W*C�B�:1��O�D0���P��/�i/��".�;/׏�*.]�D��p���d���SB��ڭ�r�\bl2<4*�G�����8{עmd�M(�:�_�V���R�nC�C�{j��*R]x�ZX� �+QPBfL�9hj��s���z�ݶ
������C�/I��M�j���t�K��7Z��ſ>� �������]���g�N�X?9�Qg6�"������ĳiq"�����g�ґS�x�`v�Q���D��Var:%��±70��x�&lݴF�Ў;,���Un�I��p�֝���~��O���"�X�CK[+ZZ�Q�d0vꔘ��JE��8e�U�6o��U��ơ8z5�����ټ��,g�����uHr��8D�{s��eҿ����@�G��Z����\����d��ZfX�@9�`��v��k��S��3y������T���O2�1D�~�:��/�ʵI��ܕu���z��+(s��_�brrNg n7]�k�y��N<����0�����#Y"�L���R�Z\L�P\���ܰe>��#�$E��x"�����V������^���|oF�]6�'�JNc]��سs+�l[/26���� �&��܁cx��S(\r���}h:2�x>Q+-�-?[}��0���:jC9����]n��w~g���.x�j�6��U9�Ȭ�Z^��r���K	�&U��o�v��Bgq�7�p�-/�;)MZs�Y�a��^�����%����0h�,�����`!W@]g��O��Sgf�i\o6��dL�ډ5���J47]|O|�UE�~n\H��dr#q�g���a0i�@gpCg�����*�,jET�,t�,�r�9��ÍSW'����L�E�m_����p�u���G��>�|���-X�v���#kA�%��{�B 藨���8P7���_��7���`u�30�@{/���bN!L����:7t]32��A�@PK�-,�64��1��=&�bz�td}H����uV�
�N
I$�P.�$�߇C �4���s��P���R�ѷ���j�p�\��BZ���J&�Y�6�E�LGS3�nb���:��J�F;P��}�
+�r�L��9�a6 �}����1q� x��$��H��z���y���K�E���z�ViB���+��D�x0�ڼ��_��W8�ⵟ�.Ԝ��&�������k0:�hZ_3f̨6���$r!SC�"j%n����� e��
JP�l��8� �A11����}GdШS�6*@~�|���\S]:sa�3VDtID��efRy��E��q�#r�����m�A��53֩!�	������ں�����UM ��Fd�Z ��ٍjzfvV�0Բ�c�?�:1T�e�F���T�UD��B�d	����rᦛ�H��#�<$1)Z�7,ؤ��Y=�9Y�j0T�X�_��޻����ġçD�������A�ŷ6w �= gs'�&;��~����.��Nq�f�a}%�A��v�2���Ύ�@�m�C%?yRT��jY�D�ft�������V/��L"M���Ut�5%�B1���׃X<%ל����8�+��ar�P���ݷݎ�&?��(R�%ɂ��eP1T��.Yj�G�p�H��ӗf���!�1�D��݉Z��7���"��\���4q���A��� ����;��������.�t-��a���h
���Je���2�?��Z�ipp�����+W��q��D��(Ώ]��Nbf>�z�s��6��F����"q"=�\b��󲘯U����F\�.���k.�|�����0��?+܎�-b1�zi�[��k�!�>�ɻ��aif	�M!At��
�N�Ui����V���f��'���j���֮]���?��!�X�Dx�"�"B]��TG��G�b�R*�ǟ<�����9��D��IZ�S묱<�
ir�r� ��SR�06�]�{��CC�z�2�&&Dc8?7/���7݌�/��ſ�e5�H�Q���o�	��c)v�?�z�\
���0azv	W����b$�eͤ]��PMV	q�������,�p�Q�c���0i��3���_@E����^���D�)I�"-cxt�����x������(kpڍ(��<v�R	6�[�t≨d:�̉4c��G��S?��!��9҆�oy�lX%�Q���׃��E�C�2.�dB2�E�%�ǅޡ~�}a_���0��8�H*Bw�R�K�j!-v�N����gq��a��jU/�߱�J7^��h�8ⱸ<G<���&��O�6�''dY�3�*��HG:(a!�LH���χ��N����!^=�x� ����ztm �^�9�����Zj�A��E�K-��x~k=��'P���'�Vn4w{#L��FEP?>�
�l:;�j���ݸiSf�L������"f��073���/����T%�*(���L��፣o`ffV��I�]�r!�ttY4g�O[�Z�`@|&��˓�X"%�od���O���1|���n��߄4f-wZL ���	�<�N��˧O�%��G>x�d;���<�Ɗg)̰���?����<��G���/�	���l.'Z#�b�2vZ��[�4
����"�A1�$Nͬ�����,,�nt��*ъ�*��?�͊*����ҩ�Z���p1h�˙Ʌ?q�:��6���	A�)�������E�׊ݲ.�����!���b�~~'��IK+8~t�E��*�	��f����r8�
at��|���X\��:�����-�L�GN�9�����?����߉�>�$�������)l9�9п�R�����CWE{ȅu#�p[(k�bɠ��f� &3�Z+x�g�puf	M�.��PTFZ�eqgԫ�.̡���G��6���ΉSg������צ �[rU�&|��G:�����~e��I�r�3���� ����� ��lV�~9�%Z��'���)�-~c�)`��|��M���"����4~`��L��d��I�ɦ��OCť��х��	%e�(I�����,�n�J7��EO��LBf�����af�+R�&R�(��!�/����8y�-$�q�]^��]w�.�Vd3e��F�� �k�j�y�ɬ:��,ep��1kF�.Е�J[x,P)ga��a-g���@faV8���l�`W�^���r�.{����,����z֬�W��L]�*�1R8B�f�}A�\��&��ͥ����$֯_�+W&055�|�"(���~�lY�,��~xZ�D(��ަ��B�ef���TE�{�9e��
�QUn|� ���pǭQT���с��0nIYbcD�Z��R�7�`��A��Q)e�;����n6�?CZE�hQ-C�����tj�O����A!��ZB���

���̢�]0��.dTN���3�/�bw�6���&&�[+�h&j�)��NN]'ё�^ܲ�F��LI�Y2�D,����&lܼI��yT�WB�<Hy�s�a�W�� B�f�)���������E�ޟ����0����B�g�Zߛ��a0�B�!UF�<��!���В�ȯ�h�bP�B�����p����|f$�JJc!��6/��l8�z<�b��s�v{���łHZ_�J�M?|�Gx��O��N�a۶-�ϟ��.��;�$��Ú^P��R�B2���9N\�&��ÕNg�G6?�G%}5�j>���d�d����Po��
�\>������+���Z��+F@�D�>�8�R�D���;�OЇ���SЮ*z�L̈NhǶ��l����8r��+���:~�[P�3�M#�-|.�*�n��\.+H�� �a�;r6�H�r9$�9ak�K#RjMV#L6:�2<�&Zy+)��Ѝ?��{�2T��t�Fs��2���W���n�B6���'��1{�{��[l���w����0�>Z�7�h�۔�*�`s:1%S#��as[�����_��^{n�Ͱ�⢅�����I���4�.�A96�߅�����q �Nc�����35�.^�k��7�����o�&ϟY�	���2�����b�/4�#�V��ǋ���KqO_?��GD;x����
��������􂇭�J�v�V�AR�M4��AڠA�r�x���D�9���	���ԒAPಋ%:�A��R�J�=~��>$�:պ�X����HƘ�����e%C��`��+������K��]%ν\V��{#%��ϵkW�y��Mgv`h�:��v��G^����ӿe�
��k�m7����ZV�M��ء�O���tbh��ݝX�f5����3�g4������(�c1�����4�N�M�]e:�9]���ds���H'���͡%BkK;fg�1vi
ٲ����W�0���d��Jz�\�T�b����)���ZY��b�,C �:�^�zP���5��"F�MD�Fmf��������7��G?������rI�=Ԛ�:qJ�NR��e���}�N�[|��?��<�g�L\��'��p{�r�����{�W�^�����18:����߁������`��`u�PP���"*�u�V)KX9�άz�㘽zVC�wmƝ��&��9�/G�"�aA>���m�?��?��,9؋&�R�zϜFaS�����u�E:==���9$S9\�6�u́VD����֋�j��QBf�h&YI��0h�mPQ�Q�ҹ��_ѥ2
�nu�\�����X��L��T���2��O`��vX�>z��ع:�W����� �E����o�8���E���3��Ӈ`S^?����|�6�ϣ��O��L:%~M�&x>�S9�˷���+p��شy������>���׿�;�
�ۇL�&�4;bV-i�*�ԛ֪H,�"9?�pȋ~�1�9��a��aF�7�;��v߈Hk���3pX�ơ����cnz
�R��&\�uX�~-B-~9�~�ӟ":��,59�m�Ee�=BŤL�n.M�f>��er���X���\I#�(�|�ȶ����K��U�8�&rx'�F�� 6Ya��� �2���[�֗q���65���8z{{e9{�ʘ�hk2�n����q�;sNL�H�رy=z�[5}7�����
��Sx�ٗ�M�Y����_�?�×��޺xMXH�ŕ��3f����gϾ�C3J%�Z>%L�:�Btt.7ʽM@�=;�H7����#�5�!��AI����X)�ҫbU_�P�<��1\�vu�@���8��o�3���AM�Q�1�54�+��;��
"�@���Ls��T��(��0HUA9R3�h	���Txe$L^���_���`�h��m^��E4���$� ���[��C���"6�:�Y����i���؁���O`�͍"�+�~�lE��Z,#��a�(�5Jg
��U>|D�3��ۍ�n�n'iZ�J�gR�(�u4��R��P����ލ��8����a)]��@�Ș�W-�+��V�1���ed�aR�X52���C~.�@鼶�!W(�o`]=݈�E�=���#MG+�F�������ذ~�U�N����HkD�U�Չt����8f�ydk��w���h�	�#px���f��+����7��*k���Z��J4�MB1���3j�h� r�ːId"6�O�w~�c�Ct.��׆ٙ9�x��X�
Ճ����a���p��E<��Ҽ��b�D�#C}0�
��t�s��"��z<��C���X7!�Ջ�cW��w�(�?�2br��A0Ll�e˚��ՋX�|A�׬�a0���m3�ߓ�bi��?�!|����>LOL��E4n<Lzlq�h��m�����\���l6%־�>,.�09��x��v�Ýv��Ԃ2Mo�P�t?ͩU~$DX84�����b3�X��(�ᴐN���&�i�r��R�P��;�ЩE�^n[݅��/���X_)Mfߋ�d�����}�}dH��yC8x��8,����)�^;��[��I+c#��taS%�)_*�uz�)�@.�����<�����+����yER����-�[T����c;���p�=ؽczۻ�j�����'0~i\��6���imO��b�D4�||�i��yډ��nx�>Y�6LML�kv�w�f�#�W0~m%���_g?�m=09���ڶT�H��˰l�ifA���U��9�7�	)t�JҨ�_Ë�a��:�)����%��g�2�t�G[�'��0��9������Ï!�a���j]^�H������y����p8=�fr0*�޼���:���,�L��D:{$f��#GD��҂]�߀���_�w?���{m]ð��R��`��PJA�`5�X�����s(�����y�Z
�i���rˡͅ�Sgp��i�4�&�    IDAT�k�D{<���ݧռP�%��(��ۃ�գ��)E::װc�NY0y����4AFB�p���E/��k�q&�|���(K��Z.�.�f^/M�I�43�h~��Ɯ��H9i��k�"[V��H���k1��WP�ObUO ��/�}�	l\Տ�_��}矿U�afr�/_����X�~�,j騚O��50�M�6bhhSSS���&f2\�������� �f���o~C�}�����}��I|�;?ľ��``h*DĄiČ_��Y�℗�Fq��1(��N;���ᡣ_U�x�P0�t"�d*%�;:��t��XXX�7��M1�ѱ`i�8;��b�N_ ��ع};��z0u�"��~˳�H���d��{p|���[���Z�����e>/bZE͹�gAܼ�E'�(�����Э���l�i\���e��!L�?3ǓԾj>].�O�s3������"������FW���s	aP"�\�������vϼ�V�Cѵ�k�y�8�&LOMK�3F7�Ao���Ǟ��?xZ����|��_��g~����`v���m�8�.�H��0%���p!��¨����[6mD6�C2��|.�4b��������<m���Y��q$�\����݉�n���p�4��<�,��y�P�R��0�Bb���(�z�61_��à��o�D5T�*�L�*�J^| h�V)U�a[��D��91�rY��}���5S˅�Y,�d��E|������=�6�Y�s��a� �w�@1��lc>�Ի3�ҕ�8��!\�:!�$����^lݼA�=i���$��('���s����O8?vY�M����gx�g��s��\~��1�P�.s��*Ԍ���5S�y�"��#p�tB�e�5Y��Ќ��h�H=!�G��u��3�4R�e�;�;�c�D"aT�%����C��.���OS+"�p�v�fu��-�m �r8I��~�.�՜H3�z���I�d���&�,Q�.�\')q��>���
��QX�<�O�0]Pʡ�o��w�M)`��%aa=��O�m��{? �K�t� ��f�e�/�q��Yėc"/��t���]hn
���Ch�4ʲ8�]ZƷ|�΍��t#�㾏}�H _��x{lV_�<�u�>�yu��G���C�������,��3�8�ZxU�z�3���7J�0M�#��I�-M��m��hC��kWawؠ0��\���FkW/���OJ�4�@M��0�k��f+2-cU�p�2��f���m8�If���a�H^�nyl��'U��>�8��[s=d��/n�y�{_D��عe'��A��4��b-N���*��^����N<���1um�rA�W��Ɂ�躻�W(Yo?���yq��{bCB'���i�\v��)p����/E���eplj��]�(Z:��?��/�XH��ʀ�4��(S�,{5����$����:�[���,��;d��|j�mmR�'�&$h���#b�Aڝ����0���c�ƍD&��
/<?��brr���PV����~9�z�s"�  ( ���0kk��6��l��0KR1 �$#�*�r~�r�����f�kf��bAQE�{������g?ь@ʂ��Sf6�y��92�)bV�Fc-?N���I@�S=8I�}ԱQ��<$�ɨ8��Lg3(F,2�e�����LZ5"]m��[��+gc�����Uد7v�څ�˖	:�����g�j1#';G\I�kjDN^>�h0��I�Jc#NT}���Y8` �n/~�u3j���W�ۃ{{�?Lcy�Y��	8=9�&��H?%�JQ�pW�j����1if��/�-?��]AS�n�#'/O6CZ<�3�k�T?.n�&-A�=2�iLE�J�����H4Q���@`�s�{���pw��epf�Cms"�6 �5ȵ唞�0���"Ҧ�	B�lKRj��dCH�����c4�d(�gx,�BR��JZh�?���`�"<rǵ���Z��5J^�GK>FAA�L�i�bc�J��+##n�k����k�t;`��1j�(9�؇��:y����!;'�p-��pL�D�]<=� >����x)�J���$��CD$Ȧ@,Ԏ�G����b�٣QYV��{��>f&�z<�A��ԕ��8y���O���&ׄ��O-�=#L,�h9��J�)
���>}a�wt�f��FCF2
���.�8M	H�$@ a޴�����Rp]0N����% ؝i<N��I�h7ۤ�%ՓtA�pD	`NF�գo�w�t)V,[��Z�r�_��ǌ��-����^�?��,��p�$4�t�W_��=��,+��ų/@��2�ھ�-�eE9���%=�`��pǿ�m��jØ�c��^���Va��K���QE�PB\eu-Ba� (��q/no��f����@�W4{Q���b6�C�76H�,֬\)L6�"c D`2Ao0 ����#H5��E�2h(�9�5_�B[���
[��V ��zg&"*�,��o�`r
��;w���	kK�H����2���H��P'�H�>Lxx�p�B�a0r2�@[NޅQC���=W��7߇�a���å�3�bi�y^�����O�L'���λ�HF�nYY�>|�=w"<��<+X�1/�f?����e�\.�����]w-�y�mx깅�x�g�T"澡PC����H�h\�YBLe�B!e�G��ζ��0���A��)9S;;|�=~\��Y#8�� �I]�f�z���W�E~Vv�����Շ������f���CN�AH�\*#�b�L2(_HO�8}�٥c��� �kF�fpF���Km��DSS3��]p�J�gR��.`"�-��/�0�.��5�����c@��>p?�
�1d`?��B���`�: ����t}���\���tr��x1f��8w�Y�K�=��L�È�M��+����#��������m��ֿ�d]TF�6��NJZ�^V���@��M@��hJ9��t:e��X�C�2� �#� H%��Rѓ�HX�
rQRR$��d�)��w��ѭ�|1����`veAe�"�i;A�_�4=��B	Є\#�jU�Q��G�h(�ښz�_�3�V������w_=�;�^0�H�N���رc���â������+����<］�e%���K���F�8Z�d
E�H��hhl�uJ#$���^�2�(,̇��kl6�c^?��^{��Bq�54aԨ�x��G���?��[�����pG:�@xئ3-���,̸��A����d��e�k���n� �l#�A�h�Ǭl�Y4E��:&'�����Ro�h�$֞<%��*{�YP��ь0����@�Z%��#p �ܘ�P3*�rP^��A'Y�m]8v���0z��	O�V�N�M���~4r�@$I���P�؉��N�a�U�AI��N�8��Lu�/_���l�p�հ�u8r��Y��\\!z1Ó�'�'�B�N�D.@�p�ך�6�7�a�W��ہ#�K'��Dni��h-6��V���d2H# ��ՒL�����ө��I0��̩���nR��-�J�4zfw)r2�	�x\b��̋y����pJ
rr��q����6+8u�����UP$S� c��V��:���씦O��ӆg"�MG),���͠Vo;M'�}*RP������Nw,=y��l�jy�����b�a������8Ƕ�3ń��MS��lC�Ǆg���o��][1f�h<�����gi9�s2�m�����B��ik�cɲ�رs��r<����bA�)�'��a�!77�9Y�Ծ����iqzp�?nÄ)3��/`�����<v��*nj,��qL�@�v���HR����L����t��6m=9ǡ ��������GMM��b`��@ۊ` ,��Ǜ�^��`��!&U����8��A4Ե"�4@eɔ�g�ʑI����J��h�D(��lI��;$5e@8�D6	��8�Hh��D���5'Z&��ǌ�ɢeg���p�q�%�'�?�<.�9M�l�ׯǈQ�� '�TY^�4��lԝ��WII�DB�z���FWg'�O��&�(?�F�@vn��!��DLr2�x��վ�[��
���
M�tbN H��]4���!"�v�T�%�q�P1�{&u��Pf\uv����Y����f��P\�N�p $���`��\9y�>��9��j�e���k�dF�k�n�rK��+���!�x0e@���"���҄k(�\$!]��r�)1(����H+T�lRH�洝Z.�p��:i��mq_�����]�e�,F,��a#�f���1c��&��FcA333Q�_(b�|X��"����/�9�'���V(�|M̂�k�7U5�p������C��M��/=��o/��O>sVbj'b	>,xX��&BG����$��*�3Í��456�s��H"���4wR�y5��ځ��D��F�M��R31XZ�Y�(��jG���XZ��b��ZO6%=`�ʃՙ�cK����wF�HB��"�
�@3��`����!���nr:I� w����.�<�3Gz�᤽%b,P4���0�g6�q:�[�v��%e�f�Z���=(,�
P�jT)��mںO?�:*SB3�M��\���"q�$��hԋ�	1��ۏ�_�> ��'��W�2|�t!�Y�
O=�L�C�Y�R��b��lE��{GJ3w"�����#��ÌbS���.$F�	�F�?�5'��V1�i6��SK�tˤ���L�F�}?�kČBmu�^X&���\��V��lԩɣ�Y/��8c�h$�B4�G����2-!Ŏ�jII�P��jO���I8���I�L�Xm��0��덒+K�u[S=ꫫ0z� <���p�B����?���ǟzJ���ښp���=���R�,&�!d�X]sB����@_%JB�����#
��6�{��֎V���K����}��� �;T�(��d(N�J1!�LUW������4݄0;M�ol�Q��=�0d�{P�����B,�wj�f���,d��&�&RG?�S�k�@��]���^0� �5 B�&�@ҳ*-��<G��`�S��)�d�M���\a@=zD=N�x��y�z:&G�r8e���
���R"0EiT��3`�����y��;1l� 1��ۅ�1�3d����:ڐ���re��p�d���`N5����͒xLQ휆�ؽ�^z�X��Vqu�����7��D8���_��f���]�I�S�@��Ӡ$��VJg���_>'�X~-�~�@��yg���8�v���Ya���)2i2QP���
���'�\K��`�
��S���lX�^$4:��;�i��ZN�R�2u��1"�h��(f_0��g����Q�eeb�/�JTa����6�)�	�o���,����^��>�;w�F�ێ�.���l+��b%�<��� ̗]z1rs2q��@/;��2�����h&N�eo���{k�/�Ep8lb
�q�|��z4v����2d�lܼ�?�P��z��8�\b��%�c���@ˉ6���&KG%M�Dq�1�X�)p�;1
!��@���)��Ez`�#/��9٢=^u��N�nk�1+����(ݪI��:�D�3�q��_�M�1ڌ�gG�^�hih�(ݺ��J�~��=p�hԚl�FQa*+��`�6�N~�z{���`@�ێ��A�1�ݿl��̪����ρ�aƁ�w�����z-�� � _`*�N�#!���׳J�k�,i����'N��=�q��)�ǟ{r�3�巻���)hmn�լ}�B�J/�0�� ���P��	i��_�gH�1zb��"P�x6P*&k���6��g��l�
u��O��֖&��!��r �������$x��ә��Կ�5eX&�2�6����PrU��4�t�6���[3���ڧ+��>i^������<�h7O�5���D�u��-0�{�Gt�Fm�
_��҂9N<w��q�صu#�M��G{Ŝ�M��A�{!�4i_l���ǟ|"9���ѣC��n1�}r��#�9�ȟ6l���އ��N�د��F̺�"̻�q��~Tf'R4� ��,���f�'$�}��l��3�RX�i!��&�����)���qfR�k�{#Uc���jF�>��֩�6�dU5:|h�V�M.����=0x2�����3XT�r�P\a��x6,b��1Fd�D�Fĉ04E�a�(���"��Z����O�D�M�؍Q���/��;v`���b�<x02�N%׆j �P���k��a�Z�Q�gG�0x� 	��@�4�Y/��֎���B���h6x<^<�䓂�Ͼ�2DCQ�xH��͏�彧�Ai.�d;y�['�S�E���X��d�f��BCKm?愕��`���G1�Q�q:�I�]��0��ԡ��$)4f�Y�pd�A�pC���7#ļ=�M�@1�JC�<�*>S�,Kp(�Y��jM�-�-7���F�WP� �"v��HF���-`0[���tԣG��6�ߚ���>=���7`����g���i���	��s,D���MM�R�̜1#����B)ب��&��/[�b�]�ʴ��׎sƝ��{,ƳO<�;ḙQ)V�1�w6����oA�y�	%=�ϡV�tLZE�!�̀0-�Yqc'E6��/
rG}V"����%".O��͵��u@�3)�$����3��:Ģ���"$�I�x\'�\8L�m��:a2��vY�vɚ�N���	��eZE��pD�;C����&	�5�m��R�uh�?��Kp�M�㣷#/#yY�x��'p�5Wc��)����ho���	���Ĭ%/�X� ���e@��6x0z��ɳF�a,�B][���Ͽ��<ל�2�=�>��S<���GIi-�J�@5���R�J�����>(�xN9h�MM�С���[(�GJ�I95�6>��5IKdG�t������:��'nm�Fh,V�
K�QP"�Τ֌(�!z����H��A꣍D��HE|��ZPQ����|����^���w��lǰ�C1�ap8�nX���x��WJvf*�Y�ƶM��fշ�:|�xSfN��ݎϖ�O�ͻ�]w�~��=U���Dwl�ZЧW�Q�֚��#��r��"%,��F��(����'��ƛ�,C(�@(��f�w܎W_��*�Br�$�+�Y6��H��V-�Fi�\���i����Q9�t�e�����!�T1%��6��6�l���G^Q�V:�Z�p��a��d1�2QX����F��Q7�f�!�s$���Z��0fYMjL�0
}zzh��.�M���W+W���W_s�IE���܂O�����3��Y�I��_��cǎ����#�`δ!��Gp��^������[o�Æa��طo��#Y^�hf3��ࠞ�A+FZ�YWC�o�X]�,vt=���ي����h������?*��o����i^&#tE�A�ou��Q̵c��j�uѨ7Ia�5�X�����'Ź[%��b�'�8��'S�Ќ���lD$ԅ���hj�G#�bI��n��Wv!�4&�Li�A���kH9�V�,�v�Q��L�Q�������̛��/*Y����������\n�P��]�6���� �_1���l�:Ԟj��a��3'�oI&���+��Q��׬��+.Cv�����n���gkJ��)� jr%#5�ha�-�N+��qæ�<�L�5��oGN����q��1������������]�0{ħB-�PN����P�ɾ"�V�B~NaDP�D�9N�4z%c��9��(k��$�Dj�UW�l�ٜ��=U���F��:�#����=QַRf#�#D�4*R�{@��J>3s�W6�0�[0}�h�^��'�B!L�2	f�--(*�`��Ps�%���8@r ��a��9�3x 6�¯������!�3i��Zl�i�d
~��Z8mV̾h
s��>�7���S��� ��&�&*��C��&�m�)�Bܳw    IDAT/�́0~�s�w��m��I�������8x�VJ�h�(W@y���K%J����IN_)��gCJ%g"�K,��0�y�[�]I���E�,���0�R�e�A�q���.ҷp�]�-*DF._�A�0>Ϥ��N��0�N���t?؍�)�b�0n�l���f�4���d�h�On��͓�����4���v-�dA��#�xPE�f-�r���K�m��'o�ߏ��|���Ϻ�D��e:F
�V�M�p0#�@�Q�����۰e�:̾�"�}�(�+�E3f`��>hh����+S�WW�(�rRz$[P�BnN6�ˊ�!�@T�����+V�Ľw�#ֻ��{�՘u��t�#���6��iSD�D��ȸ��܄y�'�5Ґ",v�jp�C�q�8Nm8���rA�HIR:n�ic�y��vA0�RDs���&�ԏ��P�Й�Л���.����jC�q�T�2b��+d6lR@��&[0Fn��{�A� |>�8Y����bPЧO/de9d�<x����[e�
��e�ӹ9
��U4�KgMĄѽ���゙S��'c����?o��A�$'��=��nj���v����ڊ@4WF&�+�QQZ;i�86��<�����/��_��Ɂ���Ͻ �׊��__��Ji>�H�R���-�K>&�-��x�rz�LN��gTnl|Y��:\/\�:>
I�9e����mm�r��&tv���Ǥ��*(�՛�8�1)�����5II�l�b⤊DN�#����fs����ؾm�����CF�����&��q�P��: ��(�lͩlڶ�pFf��P�5�{nƒ�`V��g�}��M���g��v�Rt�(da ,@ӿFE[A�
�gO�T���I4F�k��f���I�A��u�X��z��У�(K�Ř�F�駞�����^�ə�`��?;+��bC��)mO��$�VR�d�b�)���2ĝ�t�A�*f<z�>�a'��k��>�a������b�KxkC#~DX�PA�΂��YE���鹦H�V�<^h�MgPEh1��$3����p��0S�Sز�.|[���W]���rtt��g��ر9��������o��N�`G#��7_5.x�n/ʋK��Oc���8g��28Q}]�6��䡤�P�N�߰Q-,(F0��!�.���	NE�`s�������'�)���?���x��;����x���a"]cB4E�#-كP�Ђ��E�U6��š�SK�d�u��S'Ip'�
Ag�!��J� i�� �}3�<B�aoV��rD;T�5U��kkS
�d��BT��ٝ���@�
�M B2#O��m	���I�
A����1�p��3�ЙR�~U�.����p����3�9z}���x7�0U�P}�(�N���o��Ѫ��h���̙S��}7�O���d��o����zc��sq���h9?d(4	5�N7"MZ1� 8!��d
���()-VHss�D�x<Ntt����ؼ�0��܍p"�q�åW^�w?��|��y���Xh2W,mr@��mB�R�YtҶ����t�i��[xO������yI�#X�B:��x�xVPw�����*y��O�3��2���Փ%&$t&E��5��_��x:�,�V�/uJb��n�qo��EK1bpo�<c���%1��x����;q��Iغyv��-����&J�7k��#'���)K.�1c����ǞEv�^�;�m��W^�aÆ��=�q������r(�{v�&$�)> �H3�TJƹy�[����8ZS��V���C�%ri"+ÄG�yS���,Dji��H�H_F80��n��2��x"*�29�����a��}�&G�3A[����
՗����-�8q�0��j#�YeV�Yȭ��Ņ@R��F-T�(30����5�A5*�4��F̾��V5a\w����x�'�Yp�]����ǖ_7c�1��8R}�����BEyL�q�s<���
��o�J��I�����bX���x5z���ۯ��'��.�޵.�={��+�=,�>�R"�!0�����!ΡF���6x]���bJj��h-���Q����o�;w���.GvY_�]���Ԉ2���$csn4*TG1ɹ&t�TR��I?�T�Sl�A�-�a �@&6�ZD�Vh0CJ#Y�|Q Bֶ�6:|��u�b���W?�8��&D�.J�4�j	Lg�ˈ�L5��It��b͘9i4r2���O%_������l�ƺ�� �p���q-P�<j�P�crP`qg`Ն-�����1V.<�ld[�طu����K�i1~���8�Z�	=+z�l4	+L�2U`��l��3��3z��D��.R0�_w���c�E�w��ː�����`ӮC0�3�U�A��a��D� �Y�Ѡr��6@��QN�,2n�Cj`�Fa�6W׏��N�Bۤ�*�?6��B���&��JL	MIs���8~��!��2	TX�J�uz2�n�ҩbJ�QzB(�4>#���k�SH�ԙ��e�ЕA��8���Q1�-?�<Ii��_:ƿN.�kEB�JT�0b�v�*�Õ�M�IǼ2?�
�e�ƍ��PVY�P4��N6l�+���.���v�Y�\�<�pn�
/?r7n߂�~�3�M�#=����K�[p���1K��p�`6)7D�D�)��禐��ayC]=�5�

���ª������G}k�&+.��rL�6	7��q��{ ")�H��A}15r����h�(׊����ʖ�t\�\d$AB�V*�S+�;|��$r���ŧ�V���s|N�IcS�hg�TtN/��,8����Dr9�4:�Mm	��#h*:8U>:]0c2ƌ*{yRqN�j����i�9s�6tyljc�ҏ������ ��X<�__~�5�;�݆Kg��у���˯��a��Uغ}�y˭�߿�=���S���DQc�f�.r��a���1$��ό�HH�,0�Z;�����W�I���3��?����{����$�^pJ�'}�ӭ��)��R�%�Gʯb�ÆB�5N���v�H3Ph0�f�\��c2����)�*�G��7����ͨ+����'�P���s�����/_i�jNY\G����I�0zD\u���j�7�X�շ8Y[����L6;��o�)A��'���L:�[�����7����
�"nC�7���&|��|�յ`��q��ֻ��6d(��e�h4�PRV, C|�.W��&!�y�V�fex���X'���yhF����r�7س�0�[;D��Ѓ��OW�w�N}�ڄub�uHc�􁈪8n����4=P����תD�N-�y s�#�Y'�'�&�q�E1�� �x�G��ب�?@1 ��f��0���J�#>�@*�*3���K-��w���ʭ7_��R>��g��,��!%X�n;FF���W�FGG;��?k܁e�>CIQ���
\��V���|�L���0�on�t
���*�+��/a��)���d�Rw�Z�ɋ�rŰ���|�i������Qt�v�C��\wZ��$a��Ջ��N��i6l܄�;wc��~x��y�j��X����vDIe��a6��� JP5i��IMY"�K]ZR��8��r<�P�K�<�F/�6�Z����3j�	#��ĉ8|� ���a,�� Gi	<���#WI~�x�"��a��EYl1���A��e��c��"�w߿�<����6��۶c���x�އq`�v�9R(��9��K^,�C֭���� ������ &O����k֬��E�5`ŗ+PYQ���ACm5J
�Q^\"�.��O�Y����Nق��ǃ������F�JJ�����Y�ƖF:��O��OVa��j��7�I��lLX�H�,)Ӣ�T�3d��g3ĞՎ���	���?\Sk�S{�HT'�W���-����ǏF]�1�a��r������Ȑ�=H�u���cwIm�Iq2��6��a/�P��n�k/��������_�2<���"� ˧g�X�hZ�ڐ�&p��!1��c� ���?��ن��R�L�8g��}�zn�}{�DuU5�N�"�}��=z�2=4�.z�6:`G��4A��p8$� ��f�C�MOMaԈ��ƶ���s��k��p�E3��o�cO/�����I-�V��NS;f73_9�1���JH�1��æ� �tJ�f�����ڂ綒ġ��mS*t��������Y��6���彐���N e���+t=���J3��N�/u���Π��A��7̆�����=�A�G�@\h_{�-�e#�ԃ�^��Y��J�<ق��8]6���+�9p6�G�U�p.�y�������`P�>���Uhkn�i��f���;��5d�@�.fd8���]��d����vR+�F��zX-Fq���NG4��;Ǘ?l�������ǰ�}��ݷ`ۖ}x��נ1{c./��R�l�̓���E���iD'�8I�d�ts�1|��N�Zb�5��ʔ��!����)��ZXLq�eV��hCye?x��⤑t$&�QO��g� ��{Ļ�I#}C���@���?�E9X��gtv���_�D<�o�Y#Y�.��H��֭[�����"a�fg���_��~ݱ.o&�v&�>.�
'��`�ҏ�	��O�2h�h�A��b@��}��a6Ԝp� ��t����-l9ݥ,��l�Ӂ�� -]�7m]��i�W^������UX�e�0�B1�+)�
���4�^�G��GGf?�/b,����PΣ�I~ݾ9.T&+I��p�O�]�a��b)���Fv��,�s�����/��k��mw7������Νn�9�6�Q����A��dQ��1�%�;�ʜ����2&�4M�cw�|:+��$��8%�����n�)��a�d�n6JW��0M*D�:��^9�����a��s�jC7�	����͛�g��U�@B�	�m7]�֎v<���PkM�X�u���o�o�a��͘v�yBWг�^%�����_X cXTt"��l�]>q�"u�t��f�H��!��Dm�n߃O���-�8�Er�?��p����%H�8Y�{dSG��VnN��`(�������1��D�%��4/Xɭ"rGz�����l��A'ϟ&
�,���'�W�Bq�ZZ�f����@M{~�^i.���9��m%�Ux�tgb�mѓ��En����[�x�݅(--�y�'���#����v���4���P2�J
�ΰ��o�Gvi	����Z�>Z�2�N\��i8{h9�z�5L~ۺ�ހ����L�]۶���C�GIQ��s����Ԇ����g6W�`P��p��p;�����_�^+O7��_w����;���D�3�a��Z+A�D��\��Y;�oN$Ԗo�H�4ybp�^�|-|� �[�_��i�(�'��}*���fԝ��KR��VL�y�f狞3�1"�Р3J�G��?��^�7�y
#��!n�y�c�ax��$��ko�73;v��c������(����S[*���g�Ft��M�n8�x����!�aԠ���YX��=��*�7�?�*ƍ���G�Egk+�OV��4����
_@1i�ke&[4�	�����@(ЅN'2r2���F�y�5�j�ҫq��	��(���n��?b����-큘���J1����BF<q�P(�tdQφ@��D�Ƚ�_�Oڦ��-�7-�Q	0DD�ͣ 퐉@өSh�������b�'���	+2v�6�v�)˫R&�B5�����L�4� .�h*��f�����pZq�=w� ?'yMK�����ĉjx
��N ##7_5��U�V��M{���%2��H�J��Ϲ�`��-V���ᱧ���)�0g�L��}��{�큞�+ez��0�QѢ��jQS+�N�T.���x��ѧ\q��c8x�o-X"y����?o�k؎��,C�C��Sc���>E�J�+��Z�L')Re=)��^Ξ��$�i��j9a ���P#�I=�+a7&��w��DN�G���&�6�`��CQ�~H�Mbh�:g�'zU��*�ty�D�ΌN��$:������_�l������gଳ�������F[c#��Va��mX��W�0a,^|�a�����A:��|����<3f���^����g�E{XZX�7__���8y���$�pZЪc6l �n��s��k�`���P����69���F��qj�	g�vư~�~|�r�0u�DL�9.���WF�D$ټ�'4��p�Є����4���^�Ma�ȹ�\��?���YG�/���6Voߺ]�#�57 A����Eȯ�3��:�L���Jb��&���3�6�� s�ɑ��b�$p�����lƫ/?��/���Vq�]�r.�s1zTV�#����ĸb�ԩ�1c�����	@��ߢ��nw��Ĝ#���O`��-�ۧ��;�_8�Dn���ԟ<���L�0^ΫC���C퐾ˆ�ZN^a��9��0�l�G"�l��x���hl�D�~�q��۠�Fp�5�J�%̜�i%
D�x�>\j�pǡ��4.�(�R*v���XK( �r�)y���|�tT�I��#Ǩ�`@���-�tT7:\�����]�!3.I��7�s�hH�0_�h;��$����a��0�����r��n@sS߬���v��>}{��ٗ`Ӷ�0��(�,�G���_vÝ��D��4�Y�0�_V}�������_����ǎEW{��n�:=�K����d����h�(gX$�h?f�֊)i�[E�OV~�W.FB�G ��g��߁o�ق�*����y�� R�h�ťY���~��!J����b�'� �F�ic3NY�Л���(o�Z`F2��#�Kd�Q�c�XQX��}$�L�脺��wB�'�?�Oe �T/R��ﵒBM�c�DEa~��ɫ�~�$9Ov��.��.��D���6�:��Erd�_wUa�ϛ%��9{�Ɯ��9pf��~򅸍�����Qx]zL�p��˥�!P@p")���sm�.�J{3�r�>R���݆�����[D�a3�$�;'ύ��]�M{���ʆ/ʦ���"J�2�S�F�/��\K�z��(M!�}��CWy�O�z�����s�Z8i�ܗ������9��f�Hm�������&爆�.�����]c���*�ӔͿ�7��8�?H!�2�K�J̘�z�d���r�&*&i�q���I�w%gI�������1�������ǻ(Hy"��$B�v�a`�R\3w��6��.�3_4~ވ��Ґ��q�i�̼<�W]{����ߗ�nTe�Y���b禟�ۦ_p�̙x��gP���9���}oS}3���˔���F�NB�}�465�����F��ܜ䉎�[D2ܸ.]���̜}!Ɵw�yq>���EFnr��Y�D�F8���n�N7�ܜ����3m�&���+���^���}�'�ˢ��4~?�BJ.���'6�*�Q��t��)N�d_�Ak)�צR��t�@�N���C*�ǣ͓��#=,��8���t��ho��d}���tؤ!��sf������w�`���"����0nx%^~�y�5j��݃m;v��/BYi)�: ���a�~���u��zd�b�i��Ѫo���dB�޽ž����nim��oĲ�@��H����i��?cT\��ԧ��ypt�����D<�\K5�fj2��4~rX*��n0D�X.RA��{7PB�8�uhc�ֆ�z:|�J��Z�sy�,*��遆�*�<�	U��S)h�$��V(v�x:Mɸ�@=fN��c�{@gK+.��t>�r�Ϛ,T�_�o�o�W���/��*�M���.���F�m{���w4im>��yxb����ޔƱg��g�|�G��3���Φ&4����eŔ��";?�-�1�Vo�R8@ͱ�(),��zZ�����G`ԣ3�ĩ�v��eV��͍-�գ���,]�+�Z���C���Z	���3�0t,K��5    IDATt&6�l(��鯥k*M H��f5��i�=���l�J�	��	Z[����)8�8�6�%pf�1�q�N�)-����@r}�c��l��H%��f$Њ��w�z=2	<���b�u�u� ��o���7߀�7�`�o���c`��w�u�u�`2���[��� ̃z���[����������I�0�w_y/�H0��ُ�hl�]���j/��,"L�R e2���Dv^�L-�A�\���vjj�"C��v=�Z�^�ϛ2-�
'�PE�E$��]�T:��M��O��D�#���n�	�Nf�1J����F�&�_Gz1��d�v���j��,x�
`��ARg���Y���I�����_я*�;"��
���}���|*�Vd��^#�k��E���ͷ�gE	�q�u��f�iu`��_��7k��q��HO����Fqi\y�y�d���Y��.���/FyY���c/`���p[]h�������ۻ6�^�K,X��{'ib4� ��(�=��uͨ���4X�݃7|��U���̹ϙ�����.�\r�I�� ��Q�2��+f2��	N��u��)��i�H��:�J7��MŠJ�'�����Cf�B�fi�p����,�U��Y�$i� E���t���M����0̼o�L��f.��|����ԓ��� �>��=��.��bAs�I�;W]}����%�2���%���y���U���/e�4��	�0�O<�,L:5z���cƎ��g��l�T����A���XV�����<:��hli�Fo�	�#��)���|���f�WX�_|�h'�\|�8��q�7EQ��\J�.�r��-g2E0,mt�0K�!M���7��w�J�K�8@Z7���Bd��h���V�?�KD�AFSi=)?Q)�P"��	�J%��X��H&�3��*GS�I�hbr૯��~~��hh�V�Ǖ�;��Wρhm���V �6����V��"n���Ő�^|�|�",�TB������!d�l�h�tx=�50p�df.#�t���b?�Y��f�us8A��3F�ơ��x��W%�����G����ʕ��=�A�ɄJG�7Ru��R��e��0�(9�Hd���{�V��""�L���[Y?�Ř�&S)j�ilBGJ
ݜ�9(��_�Յi$�1
c�k[Ʉ�K�-�*��Y*�J��6K�� ��.ǐ�e�5���^cw}�G�!Fhf�
��lBϾ=�i�:�p4��{�p��N���3&��QÞ������~�'kN�b֢��(.�ܹ�h��@�A6���3U@%�5杁 "!�@�
����_��УOlޱ��Z#TU�Q�KH��b�����`���I� �Q�i��r�+:B��"z�:Di���K�G� [Nq� xGREC�fd��lX-6�������y
�#Jz[�Ai�fl�#�t�?�>��v�����?I ؤ�ª����AݓAΛt8<2�a���R�4��sB��g�������^#h�c��#�B9y
�Zѳ,���B���R���L=o��_0_��'N��Q�V_;�o܃_~�ӦMŨ�c��[����&o2�i���ގ�������<i"�z�)�����3����� F�y&F�y���:����,)zXD��Gs��`P� �����RB�M�ؽo��m�?|X��K/�؉���/���`r{�ԅ�5]�⡨r�ؑw�x���4*.ib�񧋛��@�٧���J1�V,|I-�;�di�08�pd�������Z�H��DH�b�T���v�7M�;TI�䶚t���N�����ʳ�>�-,ܿ�3gN��ӃcǏ��7���C2��=�b����6`�ʯa�z�p�E�1ad_���⦺c�N��i=�\z9�&���Z��cF����N���8��z�rXS(L:/�疶V�������`2��+�ϿZ��?�u�-��x�ɧa��p͵�#��lu�'�J�h�;(��*��4%]�t�zZ�B���@{��J�J�w��L*c,�P&�)�Y�dfÜ�sVb:�L�h��ޔ�)-��pI��4�DR#�#�i�⃿���3W��g�|	U�c��K1b����##Ӎ�.�V���
l��;�.����������~8p�Ͽ�@z_kz���c�c����T#���'�|�M�������g��
]*�sƎAYy�O�J����FQI	�6+ڛ���ꄯ����0٭�3i4���~�wރ��v���9�?� ��)^�8J� P��qR6��Hk��:�-�ݏ�	M�F�(�{�W�tgyZ+��A�(AjG(�'5�t`��WV�X>�NA©�R�b���H��0!�L���������ab�V�}��p٢���;�L��Gk[��6q��d�1���8{�x�ӵغ�7T�"�ڎ�.�9n<�������}J���m�cٻH~Qqi1^~�5L<w2\�	ug����AQT\��G���Nl����a�`�LU�W��@,��V�=�p��8�"��ڛ�cJ���Q���+Oa��5x��`�̅/H�:RfĲ�PbqN�7u_� ��w͟�wEx��-�1} ůB��� ���2qTf���+(�;� ]��S�EM�H���s])�<�CŌ%�����j�ڠN�cάQܿ���(��x�٧��4��y��~�痟Pܻ^y�%1�Y���&�%,F�Ãg��
{���<WN6#<.3n��B,[�n�	.���� �fp�D�Ӈ�sfcH��H$��\�e��KWg@\�iŨ�sp�9RuG�j�w� d����u�p�=���4�k�d6n�w�x�C,|w��c�"d^(�.�[��X�е�h�&�e!i�
k�)��J�MuSv���zơ�A̶����/�:^jݽ�e(��@Fn>R:#�	R�I�RLκMM�cC��J֙�wK�Z����.	���Ը�o�â�`���P\���q���h�hŠ��c'��wΙ�ꋵb,ӳ����yٙ3z �,����^2,�M9�z�����CEQ1�?�Bl�e3�+���ÖͿ� ǋfN��~=a�qP�)� V#u�ٷ�Φ��Bl���(�[��P���K�����"��7^{��N\5�F��i���$����36Jd�26��۪B-��4���fP�g�l�Oo�J��8��mD�8�_gV�2ɤ��'����:���Z�5��T2A%�VF�t��#��l'��-�Q��Ƥ��?��(N��ƍ��F]} ��8q�=*���+�CGka����%��9pm�r�x�,6����1a�x���4Բ�1������K.� -g�	�;i�,�Ҁw�`��f|]>|��8t�
�Ο���"<��||�r�d�9v�|�!�۰�?�0t67�l������Oջ�\����8�%�Z�矌�����	����f���Ơ���D�.����8�=�VX�n83sN��U�l�ɠ��$߷f�3.+�G<BMiJ^�7���� �V#*��a��8�D[k�O�^�EEy9�v���67Pu�
�e���c�Fm}+�;%FK�I"?ˎk.��*�[vb��#��˭�����8��A�4�lD���J�,7^�Sq`e�@2%��,���ɚ:�[�Q(��=��`ׁ}H�b���暫Pѳ�Wm��cu�;sЕ M�����=�5���5�_��¿�Ie�*�!O{���O�kkii���eiB�H��Bs0���ԏ�M���(͠L.��3�gp�ffJU�n�&�a�O~�R�t�nmz�lS��*������L�<��Ɛ�������y�;����D�L�E�:4=�W#~T�dᖛ��������છ���sF���]���
��.��@8�ǟx�G���q�����ή� |^��z�����Z�?�<�<���>�h8uJ\�F���C�����qYx���0��=�f:�|�k��V�7�X��{��y��T��9spѥsp��ψݱ��DB*[�d$����qD�wj���G���:ݛs�"(M��Oi����͖�B�U�6N]^�I]S�U��cj�4�|�c�W�Ct:�1�����7^l�.<|��UY��������+�@g�9�.����o���S1e�$���'|�t9���V�:�q���ùg��^~ӧN��߶a��5��kEs��܌�/��a�����	�Ǫ`�P�"�.Z�-Bԡ�9J�d*���Æg�{��_ g^l8���7`4Y0�����H�gžYq\J��?XR�d��P\���F���g�S��44�.Zy襋U"?i�7nZ���|AW�;B+y?��;��1�H�ٜ`*<x�p�����Ma�]�p�L�0^��S�a�G^a^k�����S���}�YB]x���P^����ch?u
W�>��.�MMM��B޻�r9�-��@����^�Yg��O��*K�0�1n�H���رj������N��}�pڌ��f��!�RS['�P�G�����a\y���Cq���x���{�V���ږ�DH�#��У�w�(�4���4�T>���tϗ^��͠�բ/��H�F:���Jo��d�'7��hASfhq2(��H�S����zc�A���(V��;��3���Ep�l��k��A|��r���`���((*��wޅ�����K�#�ڊl����?G_z�U�Zi�+�3��-7��E��nԣ���ykƟ3�`��5<p �����bdf�%��"��<��+C4��天�74��됝��i3.Ķm{q����qA�}��;�aɒ�x��G`qe�+�C�S��1���1m���J!D�S��	��5r��;}@*����ƫ�=�W�����Eְ[�y�pe��To���1 ��J�����=�B٧�gP�}M���@��Ϊ�U�L�ɚND�����n36m�*4>������r��/���X�;o����$�j؜^|�~+>������Ź.�������A�{�Gz�W�gz�fԵ�����z�{m�L38�p$���|	I�G��$���z�@���j�+�}{Ѫk4����?���+�@��kY�J+ͼ��<�}�����d���~O|�Sp�}ǐ�dp���f��x�������x-R*��`�ݛ�(��L���������������J�;}
����UPoT��>�W�����w���{Q���&N0~q�ڰ����:>�o��n4 ���3&l�/�KG3��M�cfW*���e���Ѡ�,��}�l��������wy�U|;���eM��&[��{�p��.B�WC������G?�1���忍���[[���߃�}���:=�y�E&�Sŝw܎��UDSIQ\s�ո��ⵯz5��˸���`�9�]���"��.ܻW\� �	��d�ĉR,����=�Hӣ��{���>����j	/������?���V��9�sy��o�$`���:a���@4���41m��{�M�L�4��'��ƃ�s@�S��[1���h0Mj��Hg�y����6�<DIN���	�*��l��k�T����iX��#
�hɽ��!��MT�fH?����W4&�z'�xr �&i�t`��������5p������ʍ_�S�y"n��M�Ɨ�������4�]x�����+����x�*�Kz4���;���E|�K_��Ñ+�]���S���;Q�����]��}��p׽��{'RCHL�������W�q.\�[���dmC�nW�l�5�V��换F��e&���Z��>�>���}^]�28�b��uc�F�s�Z]�ų��m4�0Ѡ� 4�?�7������ܤ�!�cN��\c.5hS����H\�M�*���3*}�~O�H�]�e��������8y��?��}���ԧ?/���A$3g{��!�����c�69�ӄ�\��\��5//��ԃ'�V�&��j�-&��h:�J��L*����e8p� ���c���yE����6fc����tِ4_�y7�z�d�����#�~�����U����!�Y�M~3��f9���Gx.�͠?�Ӽ�}�~����p�%��G͠����z3��@F]�o��]S�?�R�����0r���L:):C�.H^;�����z,Ξ�џ?�����J_�ڷq��A��!�?���_�p�.,��,���	���x�{���gf�����~�E8w�n|��_�r���	;��#��-���Kp�E��Q�W.�jZ�d�p����eEHD�Y�eTr~aw�{/r<����ݎ�~��Ԙ�p��y6^���կy+���� 4P@�� o�v|s;��#�b}�˛&��f$;t�*W��1v����!5w�I�A2�G(J�\��8���-ܸVMeP4Fb�AL'����{x�s�Å{p�|މݻ��k_�6:�-tuttG�����x��(>�q��Q��Wu� |񳞈��ڇw�����I�W�̏~�<�ڧ��ɓ�#<�q�%������VJEݳD�D[ن�N�##�%T�5�I|�;�Ef ��=��_�k����g�������� �����\n+̸Ӵɭ���g֟���W6���/�u��XO�ti
�/�K���y��F8�Drp�#�ȎL"�̢�u�7oWd)k�t��"��>��l�&B��D�y�e�=��N�ݨcǎ}����p��/|.��
Μ�žCW�{�w��M�����mc8v�Ad���w��?�E�i����{'���|�#�4��+��?��ݘܾ?���4�{/�;��p��a����:�	M�VVWP\]�f`Ϟ�h4�Ҷ�r��+�p�5O�v��~O��,J���J��}�Ƈ>�y�����Da��� 	+���T���\,�ю��]�6DMhU��z�u�ie��8�hv�ǠЈ!�Afd��c
o�z��!�@0B톕=�a�=
"���E�&FŐ��lĮ��'>��������j��0����s*���~#�T� �W��~S�M�hL��G?�1X\^�ͷބ�|���o+�u�|�A:ؿ�z�{p��U8w���<������;T\��a�x�T�kr:�}<W�I&��������c�T�S����Y���oĽ�ާf�С�x��߃O�F��_�����at�It���C1]��bM��FS��G4RM���� ��NSa��y׻脺Ґq}�
�2ٺ��]�X~�^ �vG)[��u�� ��2׋Q=̸�h����ng['p�5Wc��mX�/�?�?��,�Up퓟���b,N?�ַ�����\����ӟ�,d�c����pӝ?�^���?�~������?��{ޏ�[��ˏ���&������4!�3=�3'�)B�W]%���²���H�,S�FҐ�.�4����'�ܢ��W?cxݫ^�ºT^������m��^|�]�Ю��RW�t�\D2Ѳɠ-*� �9W~��~�����Ѷ�8rD�?�;)ݲe�+z.԰Ǩ�fx�3`p]9�r��ެ\I���A�F3�M����h��H&�u�
����C�����Y9�Mn���h�TƹS'Q\ZB,�UF-��:�>ʥ5��m������'=���7�\\�Տ~,~tӭ(s����½�b�".��B\x`��&JF`@#5U���̜�}>���[��_��~�X�7���
b����׼����ׯ':�8��I�e-�����23�3ä$F��
��������H�qs�����L3�m6�L8��&2�E���&^v ���Ed�N�����z$����L���xMё�SAn�����x��<,Ψ�p8�#�Y�1�iZUt��x����]Y|����U�\�/~���G?��\� �c�(�4�"�}�6��)i@��I�޵JEZ�f���Oj&��Q.W�g���!kE�Z�~ҵx�k_��g�|Z�`<5�P�^����u�?p%���fN��Nv�4�-N��gM#C �t#%同���8"���9E�0+��1��%��|�    IDAT��"�i �Yv:(-,�8s�jٙ1Y�1�thV�2a����M���� �8N0[���=�$�u@��%�|�(5�̇��d��2.�d/~�w��P����<Ɔ��/|?��O142,�,N�xk�z��TV�*K־��hT� ��r��q�ܹG�|5��~8�P"�j��l&�k���Wxw=�N,�v8��V���ڍ�(�s���c#��� �hY��t�&�> @	KM�3�83��i�.W�_X����^��:Wj��ϕ5N,ި�9���Q�&��`2�GKp2��/i����7��5��#4��fj��n�!
��C�� Fw����uOz4�oF.�ǹs'�կ~'N����8\v�"������nQ�Ӯ��[��o܆��ujk+�;��߼�p�~|�k������w���f��c1��S����-صm�Pxj�|�]��bD>;v�3EQ<x�>��\��e��
D���_��������{^���Oo��#[�̓������&�=GTПL�_���xj��i%-�Z&����6�m�8ʯ� 50�@,�N/�ū����
يb֢∛�W��0e^_��D�^�e�ĕ�+�l&��=w��7��-�ʞ�����Y*Up�Ϗ�?�.��9r@c�^ �]�g>�eQ c�^��k��#�x���Ox��x�����1=�3�ϩ@�����ub�.܏L&�Ý|x
W����0̐g�&�<�/.�Moy+N���w��������oB����x��y��x���f��$-j��3?Kv�l#�_�\sw�f��~ׅ�i�N>�~��r����P��j"�Cz��H*�n(�&����`�n�#h��h�z4R 
G�2i�Aj�ր^ +@Կ�I<�q��`\�J�O���?�)���\�k{�fw�w?��ek]r�x��/�@��z_����X��08���Y�����;���>��Z�z�������a��(��/��<���u|�"B�DǯZ��C5��clr�h��sx��>���{xؑ����!|�ù�ge�s�W�mo{�����_����{��8qoc��R�p�C�V��\�PW��ԅ��v�(���V{�0fbT�q��I�S`�l�É���g`0i���(!�����~�s�3s}Gf�A�1����{ ��'��e�y���8uz���c#��5�x:���gfJ���� ���C$@2�Ce�,.�5���_/�����]�߻o��oŎ�;q��yi_|��Ш6P���G\�|.�^+�p���|�&Ct��g�GO��[�������8|ѥ8x�0�����GU�\|�E��w�3>�_�����W#�EW��1xmw6P3$�,[���k�%����I�M l
H�Z`J��H���)���~��wi %#�8�[wc��EH�lA��n��|�S+P�p2��ٳ���m�-Κm,��mx�2*k��P�Y��եG�2��L:|���U,�=�~��L0�UjcR9�� [��G(��� ��}7f��]y�����#�y����k𒗿�NɁA�M:�z��Ȧ3B�eJ��:�j�ټ1R�S"�FM�'���ӻQ\X��̌���?�9xի��}�G�ȏO�R��gZ+�AZ��+Ge���\�s�f�**��g��*�=��ck�A�� uh�p��f,���n�."Q�{�&y��C�}�řY1�������y@8@F@&�H��<YΈ	�r9IExoZi���,�B:�|�&� ^���ث��y�4�<�7���ʕ{�޽H%b跛X�9����Ǉ�w�n9���i=sŕ%�Yh����C�bKx_�2�:}�DX�3��o��&l�9�7�����#����S��ˌ��9�s�.���j��%3W��7�;�.�C$A�}� �Mtæ٢�������(lf�f� �'���0vG����&��I�{N��zv����L:!s�R�ѥ.8�3�m7����4��@�@@��~����X\qxw�q�[���o7~�3jv�މf��cǎa~aQ� ���N�rY��,�x��� !)��Ne]:0'Pk4�tF'q��Kq�S~��|�� ��k�R���%��s�[gZ&���Sv6�ʑ��2�Y�cd�љ���������:eia�\�\�$&���I��<�.��ƽ��P_+����z����:�Lp�g�V����i�q�M��"�3R�OϜԝ�,��dp�c	xu���(�!M�<48���Ӯ���?;'򪭷�8wv��H�H$�����"V�e�X\������=��#7ށ�܏G?��) ����uQi��t>�GSڛ(F'ưR����r/�E7�B�n�~��F��:
3��g4ҍ	���9�@��w��z�hkicgd���F�=�����ٺ���"	�QE�ިc��T��:yfڤ^�7��M����f�:�D-a���:妡Ej����4�u��/�61���H�c'O�~��(���9ڂ�p��1�����욉�,��Ȓ�YL�٬�Ҙa���zy[����o��z��O���z&������5PZ]�葫���Ɓ]{p����I3��h���~O�oKK�X-���ma~e���w%T޳�0���On�N�E�_�"<�������y�	LN�;%���I�/]��k�&���qHp�B�Y����w��*"Y��'��}| B*- ��Lġ6�K�:� ��H��Ϝ2mS��I)?��hR�g\��MģA92��3�-"w=R��J��Z����@V��t�ʑ�+��όWY�ϻ��r�x�;���|
������G?��6���JLo�D�Q��yܯ�$�#�JHL%��ՕJ%�?q��'q~nF4��m�ߡ\'���_�Cc����{	M��tGtS��j�g��}[���8-�9!:n6w����\�l
u���E�8Q.֠4f�E2�N�i��
�,2DgE�-j�K��y�L�F�3�V�6�U�b4*+���tР)�NRi��y������ry,���gN�G�+�C<3�H�����c�d�x���O|��"�\q^��W"���R�`zz
�z���v�Kgp��!lW�/!c���F�RG���R��^����9|�s�ŷ��}dص{����h6������� >���C��"v��^XH�]Dg�ɫ���gA��#g�u��)�7+N��H�d �E}��:l�C�̆z�!� i���;1FBbq���鯌Q�D���ȩ�\�7Q���Rf�"�N�����B2�ƃǏ*�.���b���PB�DaY�P�L3�����q\�oo|��̇?�l"�]����?�CQ�j�*vM��#�z�"MZ��F���>��;EW��!�Z���Z	G����gΝA�\�~�N��x�,�i!�Wt�_��K���4>��������*��}"�I�8��М�Q�m��������Oz���?�Tf�M;��!̢����^��G��N �t�m;1�m��m�P���Z���L�`K�	F�а)"� z-N3i"C�C.Sc�,�0#n85��LC�Vp򾟣������j�8AŒ�s� ��bBN�wkK���K�����5��7���\�� ~����oL�d�mVE����ӥ��'5�f�O�<�[�q)� <�V��O*j���*�C�ʎ�,}��_�~�x�?�p,��qQ=�.O����S�(V6U-�ѭ�u0d3,l��0�۬UP)C����!��3`Y��*2c�=��B����� ��ۑq����J�W�gf���Y�p���۠Ġ� �8�zM�	�I��:zM�|�30[xɋ���?�Ѣ2X~��1���>��shtT�-�5׫X[�9�V��ԩ�vΒY���uB&Y�wMk*E-o$��m�p���j���m(���ty�3���V���O��E4�nY�A��tkܬa֙�~�9)���_qݤ���bԯTL���La���a��i��>p.������~��S[s=�B�&��-��1-��V���;Ad������n�ΉE�5e�ʯ�|�{�4l�ѫ����sXy�c�8��+8z�r����kKo[�Z���r���)|�;�"�������a�
���8�]J3d��t�YmTZ�s���R����ŗ��}$�Ē:[=���غቈ'f���k��LW� �l7M7� �t��XT����M��}���dIД����ތ�mˆ:�}��Fy������d-�"�� �1�$�}n�@I:����c�$�C������QpR��̻ �ڦ���A��!4je�q��0=>(/����4n�IVS5x��F�ٖY'�a�����h�����>5��w ��z�4g�$k�Pвm�z��>��>f�-=���vX�}��n��|iͼ-B��`��X+�5�����(�ø9��[��/���ɹǺ(�y&{p�ޟ�l��n4��Vs�L�L<a�}5��پq���������N9�t=�5����%;H���-gsP�B�Ŭ_�M��rL�م\,�=�i�^�(	"�L�pc�09l�t:�E���EC�br`X��Y)b"���^���c��?�'=�Z��o������7��1��12Yd�)iՍ ɇ������j��^˥"z���H����v�;w{xƋ���2����ȏM�$���]��9M�C�G�?o�:���e� X �?���0qk�ps5���>p����e�/<R݈ ?������ :����l/����a�P�:������H�27 ��X<�d<f���{d����e3)mD�Kg��g>Oz�A|�����v˭x��ߨ!\<ǁ"ciq�����j��2��6�Zu���=sZ��D��_�4Ÿ�+�'. `��"'���wbx�^����j7���i�)�:i���:Z��
ɉ��j=h"��N�,��
T�+��фWZ��}���C[+�O,ڄ��g������)L	I�O}$�Qxݶ(}�d���n�&N?��x2-$,�@���vmY�w�0iYy�߰��u�Z� �H���$3���y���m��]���o�[�cߞ=��?�S��M_����P��sj���;�����.��\�U,.-cf��;��Z^���f�L������P��-��+����w�k߾���/�0}�P-�S�Kn��i�ڗ��;�47�p�
Hט���^�63~i9l
�T��Qp=Q��K(d���,6̀��Q ��B�
2�}�@cZ�$�5�Nwe�؁��=�0���s� ]\�E>?�`7�f�S-��V����n�CM�W����!���^��}�N�9l�܂����h�U��auq��a���u.��Js�ﵶ�f� ��lJ�|6�c�n���������P^\���5�3338|� �����>�Mi	����a����o���sb[?Dl���7�-W٬�l�y��NŜCB�/(��sL@���(�!�5�@tl�v����nTh��5� Y>'���,_M5�)��$}����^S.���ģʾ]�V0RB�Ԯf�c��	t*%=P|j&����K.G,���i�=�� � �@�^����?��jb�XF.ŗo�ʫ9�N����ѧ3�FGF1���������1x4��D�eb/y����31R��ĸ4V�bIV�̟my�ߡQ��D�|����~	:5c�8+c֪��9$YO��s�fr^5��&��A3�>��v�9- �s]�5iR!fNvT��C�̱ؤقN�M}�O�!PG�Md��AU�3���j#�H!�҂N�#�)_��<�g+uj<;9���E�2�_��,���p�����=�SQ�.�rp)s+°lH{���9�q��,������;���� �t�qՑ�1TH*_����_�jS�é)��\��l�� �w��g�&K�J��}��������x��e���^6�}h�����fp��f�f��ivd�=��a^?6�֬s*���k������?��U�}S��d������^8��g�u'�?�1y=I$-�, ���v�ь����o�eT\8��C���A
��/O	>���,�gg�i2+gG��u��b�x]�{�8*�!�D0:>���v#�b��V��V��@s:�v�u�6��`�ك׋�Ĺ��YF.?�H!��]>KԌ�klM��G���f0P�?�?s(	�)]4Q����r��7�,��"%�����&����.8��!��Y��8� 0�n��`�� 
�&021�f��.l�%�PCA"���a2�P�4*��_/�A:4�E�g#�	�m	�P���)ߎC�0#�:mdx���j���yԛu�6+���A�G1�m�ₚ���ݭ��i ��p�iIz�͎�8N��/�m�q��ƗF}�H�XZ.��)�9g��~��Xh����݉��9���[��	Xv�X'��u�7����0Ju��Fx�a!��i����� ��ִ��7�y�ߍ�&��@�Mǟ�7jN��h@�9��#2�j)�[�D6o��_�Ȯ�CA���Vb�!��S��ɩ�r�|��5I���,��a�\����_EԤYY��l��On�`�����)�ۇ>.qp��C��ɿ���D ���M������j�b����3��D���&��&b٬�-����	�p�#�_��~�F�����J8�fPv��1C�YD7϶Tk���,75��_�hU6����F;��u�K{ U�Jqf�Rs�t�sȪ_���Oo�-+7�f��1*�3��׺	�v{�C�}�b��63��1Ԏ�j�]s/z�cp��05Q���g������x�DR���rk��w�juq�Ϗ�V��O�NW����ʜ(�k"b>��K��A5��&R�8^������ڷ�˵>��|��d��p�&s�2y�0LC��t���Qԁ��Z�LH)"�]�Y�d�N�H��t9�����@�g�L-X,D��4M�/Z�+� -��7#�8��]b�(W4gP�ra�^K� �cQS�@˲=u7hO�(���2'[3C��*�n��<�
��U��\��`��T,����v��BrC�~3����X\-aq��s'Ϣt~]fD�>5�G?�q
��[�65.6�l��}�T6��E��Ȗ����������巢�.���vgR�vO�.���5cn��i���Cf��N΃B�ϸ��ړk�%�k�����C���7cin�g��#�dB�^>���c��B���j�4a�QX�J�F$���=�V=�c4 :L]���aN�j�Ԗ�gk/�u�hߨ�Z�+��z��B>�L�H$!:��JI̊�g����&n��f��$Z�`l�����\�(�ɱl� ��`�&,48�����N���}�F|��A0�FfpL�E?ȌL�����uR&'@
������9@�\R�y���6�'#�XM��`�repr�k���ň��Rˋs謮
���04�S/��T&��%ڲ�=�ې>�N��`��0c�0p9�Z�6/4����4�uh�vw��#,}@�@|"C#ضo�
�XJ�g������h�1���ʋ�;��W^��V16U5N"x�C��r�#�>���>}nU����j���sϮi����G4 ��y��՞��I��(7Z���p gΗp�w�;�QTAz`�^��8��!YtXyIO'�DC�}x���ak�tY����q�/'d�$�6���� �4� ��b�y���d%f���E�����ekt�sv�r�s�	�II9H��(����R@ �2�w�M�T�D}����Vs�F�YD�)v�{<d�1����l�ZK��z�G�G�hvp���|�����@:�3���j�X׼�����uzXX.a~iE��c�b�ev�M��[�Z���^_�b��o,�7O��I�/� 3)�о���\	�:φn��pp�9�/4��Ӯ���B�I5&+������k
��qO��9�@ ��cVq���U�� �2�5���1dY�#��J�V\^ƙ�'�\��'=���8rc[����.���Q����ܿ���3qx`�2�<�9�#��HD��1
)72    IDAT&c�jN���h����c�x������AE���/<���R""
�1����Pe1.��j�E��#g���Dey����J�Ұg�
�u��j��C�=5HU�Nг�4Rs��#��~"a�7c��
�7�<mzh�%�aO{ ��x4�f���p����L�8d ��v�ۃ�#18�LacۦR3�F�g_��~��p��N�����T����H�fm�:GE?�gcNvA�pTN�̔���z����&���,΅=�<v��,����s�ˎ]�/tn�N�BpE��nW�g��� ��V�a�7�%�[$B�rF���Ѩ�`ut�R��Sl����~M�QB�'�~3�ZtDw@��'���!�̈́i�p��Ѥ�͵Y�k�i��v�4K�աo���=ӹS�0��F�"����3�+��]_C>���Oy���Ku3����z}�uf/����U-��:�o~�'���?����F���#W�Y�]�魣H&#���`�I�e<u:�&ђ;Sgf�����;�uDSCBÛm��:�x������7�M�5M`x ;T`#���h*rCF u������T�z��=Yo<}S+�D�7�B��t�R5I�X�PC�Nn��h�@��A�\zh
��cDi�&����� 3ø��`l5�yuM1���|���Ο�W�c۾=����œ�y<�	_�a�Š�5ՄY�W���<5�|�˨u#&r�Z�%]ES~A)��{5�(���VWH7.<��i:�՛����G�FO&�Y�d���.��洃Z���Vu"�2d�|T9T,l;=Ov֜��A��cH�
��G���k/�����jhI{0J��1z�vy���!���{��DÉ�ERiM9	����`��?y鳰*�x �(���l&IGm"���� �� ��.����n���(�-�3��k_�*ih��;u�=s�3GjL4$��J��ٕ2���[qϱ9d'�Q��V3�E����E��!�	7�u�P�2�w��T���D���u}׳������鬵�����EHMR�z������RSh��" m�2ŜKj�B!HZ�-�gD]��ת!�YC2��#/� ;����g)��Kfm���	i��fK�(�V�|�y�=��M7#_ҫIeҸ�a���8���&�iҤ[-�8�@uh��nu���[��S3r��� �d���X8S{b�#�,�^�i���eE��$��y5�S!9�3��n�AϜUf���J�e�;w
s�ΠS\�)P4�����x#�ȩ0o�ir�81�Pg��>�i��؂�x����I���=�L �k�UZ���8���~;�w�:p�v�A<���ٳ���[�Y^B\��l-���<-�Z��{-��-EDlݱ�� :����:.��MÊ���ٜ&��WTK����g' #�L*-�"b�dM>��N�h�\��Qȏ!��	��:��凃s�!�ϣd���mw�4�y5R�!!�\s��S���H�H:����,gQ�"Jkњ2yB��P�`�Og��w.�������'u����,�B]ն���_��FQ��D瀌��ަ���5V�`P�ʉ�VY����1?7�kM7�f�*M"��:吐FT�hz���pc.��%)������M��0���b\ A:����ޚ�t���]]6�|z���+���UE�?�p �����j�M���p;�k}p��T��~ز��1��AqĬ����6��&252 С��<��!Н��u�A�c�v�o�@ݳ�S�N)C�?*;��Ж�(l݁ s��DM s��`���%� �d�tYU����>��A��p�h{�������v�2Wr!�j.C��'kj����Q��F��������f��(�1�Y7��\�_Dmm���R	�9�n߹kke<��(.,�f�x$As&I"F'4��pZ���ء	P��$��"ڴ���C��kQ3Ȧ���D�t\�>�5��LJ��lț]b]�s��ڃp"+#�F����x��h����"3 �A_��2xx�C�t�a���	��X/�bj���*p�	3�&��/��s��gD7�q�q�ZSR���i���|7���t����Ҷ��e����S�y�RCk#$6۞�d�\�������`c���섺Qp���ʸ�r-Z�'^�ѧ���Q4K���A�r}��QrcM�Q���uyn���`"Y�����d��������K}��ܲXʒZF8ƅ<��uְ�Ñ�{�5�������Sʤ����+w��G6�ŝ��׾�-,-- �Nbώ����+0�� 3�]�KgQO)�oZ:�NsKk����N"@/��h�%!h\���>dB���n2�9B��4^Hk�mNGT������꺢ߦ2�qa�:u*��Q��wh�k��4�imT�w ������n�|}�ˈ���Zhm"F��.vlF4���)�h^��B�W��'�$�N�B��Pw�u/��^T�E�����A�ޡi������e��J��i���s�[\���*:�za
�)7���\q��Z��[3�^��"���7X+��g�B�
ǣH$S�d�rB#͙�=OYR�L)Q�\�~�:�k9���)����Z	�JY��� r�S�y�fPB]Sɘ�Y����T��R.��ߌ�yx��&�6(i@��D:G��@cuc�b�.Rt/��ѩ7��fZf��I$�a���(�<NnA|����2Ξ�Aqv	�7��09���`Jt�Z�������QJ�����4j\_5��4F�P�!�Fv�P��ǟ��y�'�(Z����>Y۞ubV�Q�n��V��<B"����LGC�ԇ_x�s���&�ZNQ�ݤ��PY����K1�c�O� XT�gE��������i\�����L���d�^�jE�n�DV@^��E���\�JG6>5��°�!f�&Rix�6�x�T�U�z0Z�Qy%�6��*�����j~��Βj���<�pq������+�	Q��!��lm*���t#�Z�5�����6�N����q�4G��]�!�aqe��?���9����ݺ;v�u~�X���MM:4iq����,����"�C�V[�#^)a�ؽX:}^iI��p6������Lg�0;�3�݇ţ"��,�@�ߒ�[�єnMN�|Bt���j`�	Th�P.i?�6��E�PL��x<%�&:��c!\<�Hyf�J'�Z.Pƽ"A,��.�@��DhPq��D�5ew�/�,�<Ր�Ϲ��}����i�>���c�P�o\N\8'��@�L536!�����%�,3�-߱d��(�Bg��S%�M��z��|�?�e!��Mr݁����qa�/�R?���Q���D�W4���KV�[�5mb��!<�0t��Cʝ�A�B�c9��;1b.ꚸa�T� xn@V��{`@�&$ꗻA�R��4a`Vq<$>i��l2�ѿ�$����9v�����5��A�V7��=q�ӏe�������vGW�^��oth�v�Ď�Sr(��޻1;Ks���x���m�n�o߉hfPF#�@D��6��?#!��c	P[. �1v&qlxZۣ����skE�s�-��� yH3���	>J�P��5Q�I�%�"!���\�e�	�R��2Jf�k�kK�L�VCev^�"k�V��p2���ݻ�szZ���8y�8�M��Jc����X�c]��{D4�@,��=�� ��b��izؒ��^��e��.0o5��3)����ʛd]B�ϨZ�'w�ta�ۦ���t������P����#�HFU�z��i��m���"�A�����M�b��¦/�V��^��WIg�� ����fd�tٔ�[�e癳��y��c��#��Bl��'��eG'�����j���l^��Jy�������,���&�dt�x.=�����ː4���4�#׽����ĳȐ&ʑ(ǣ�]G�5"!�D��M��������X'��ͭ�!nj(��7����As7��<�PL�9�U�l��T�e�]F�it�M�{@Ԙ ��JEc��-[�e�vt�̕�X��)�_k"O�x
����c(��V[���cԢ�U*�X*��i ��.��f3���~D����������͖��`�Ŭ6Hg_�	���RȤ_t��-���os3��"P�߬'ڙ_�]ѡ�ц�s�����a��m3��P�C�6:�*��ڝ���T�n��U�+e4��*���;?2����R����e�^Z��! �3���8����W�Q���FS����(�j���UH"�u������5laNg�n9�;��M1���(�m��怺��(�U�.�K���ZĵθW8�`�~9�������F�t�D���[��E'u����]���L1Z��O�J����2��M#�/�ص��"���j2�h5j�JXk ��i-��΢�,�� ��!3<����ۆN;�ٳs�?}��<��c�����1L8�A�S�Z!�$qD$�])��'��}�WVoL]�L��e���笃>"������Oe�O�1��p�/k��� N����yڨ���\�1~��ěÈyy���VNsY���SSꮁۇC�>�<��p���#��6�ܗz!DE8E���g��]�DG�x���!�y�s*A�\�s@z����XaBc#fvr�'59�VF���m��F�?�nC3#q?��D��D9Ͱ��(=顙?��i��xtol�����0>��ӌj	aai�O�B}i�y@����&w����vMDˍ*�n���&ƹ�R*aG+P�n9��!��UZ���?� ��]���&����"��̙�8q�=�-, �b�'9}4:�G��u�DV�m��D~j�vMax똨��E���>,�;�� �;��)�uF�p��mT��l��bAI�)�D�#��� �#�>V4���P����lz��P���� v,�����'N��TE��Q��47Dة�n6m�&�-�{�}P�x����u��nB�	� W�`n^����Nj:����o��ph�F#�q�k�� �O�rF5���4"�+amWTʇd|E���f��1l�_7���hgr�t3M�i6��9��>S��S|]�@(�#6���>,ٴ� ������I�<̀·��N������f\��!��u�"_�c�k�H��ol�F{���A�Ȩ.�����X�=�ȬHˏ`lxT@���<��g(��i����il�ޅx./���"<[���k�&�=������)���f�b�}ƺ�(9!˓�B\���cwV��'�l� P�?��f���ܨC!��L�wK�Ht�m�;����� �R+'��Ӭ)��k����ݻ�ubR���ShTi8U�`G5'<R����(�yNN	�d�2�NS��`���լ#	!���=�<�N�����#q$	���1`���WSL�#܋��<ƶ�����w�a�]�N��H��L4�l,��@>�B�Yé��\��R�����Q���G�(�Ů!��A�x<"'`2l�Q�k�DSݜ��<��k��@��QF	����=����7��k�$�7Ǻ�H*2y���y`�۬��:w뫊X����=I�%A�H?�'K�12��[���jtb��5]צr���O_�f0��Z���T��Zy��f�Ɍ�@�q�:����>�P����%�����R�*�T�*v�!�P����h��n��8���!ǺX^��<�ϠY\R������0�u�� V*e�>y���A�:�02��-��
j��7v3�`3H]���2؝�@Rp�f ��t`����_����/}�5�<�E�F9�7��$�f�j´�Z6��gnB�h�������	�}��=��l�0�Ɛ�)�V�YZ�v!�_j3���J�@�Y�Q|��zl�ϟA��M�b�4��cȏ�c˞��4�XYZĹ�'P[Z0S
�I�p�upв���%ƦKgh65y�dX-��a�E�BUb�_@3U�*N��a2t�Er��('��YB���J�ҚyD�E�.L0n�,��X���{�nQDB�$��M��s��@�TEu��p"���}�ځ^4)�7+��0ݤ��K����RscgEn���N ��x2��('#D��񸮡�޺]4��?}s3'�mن��!�C�\S����it��@�&M /5񱄌����*;�[���l6�� ��~1���BǦja1�(�5v���H{�v�{=�~&�k�1sLɅ��1�I��������>�����j5]p?��/傹�C/~�	�3�f�R��§��jV�X 	�њ<*W�`7,��h0���{A� \Ӽ��K�<��(��6���XT~�Ō�� q�.�]}+=��J��g)`"C�j��W���?�g0j��<@��h��������A��~k6D�a�Ѩʖ)4�����܏�ب4�}�g�kP��c˾��ڎ~$�j�͚M1铤��A��w8J �����.
0n4P�9�_k�EF��e�.l۳[����y��n,�<�`��x"�P(.����xD��n�--r(�@?��=��?�X*�Jq���`��	T�K�e�\E4�&A	^��cJ��z���0z�\�0Hg̵���` ^�"��P ��f�� �+q�QG��iE���������Y�J�"�%�W�U�Ϩ�d4�Жl��̳��4ՠ�Ì�s.5{�ǯR�.9Ɛ =өq��'��:��|Q�+�%�sS�v�H���]�D�K%�>��67�u\�_KoΏ�ꅷ�a�gPi�'����M1�צ������;rl�ĖҭJi�	[��H�@MQ��@�V,Ӿ���GB(f"Bc$3�y��/6����(����k�Һ&p�)��wC4�5���jk��7�ew_�]�� �f͠��^�,��`�gl6��{��s��y�JM(AI�����9I��X[�G�ZF8W�����2���0���h�4S�㦬����X�j/柍�k�8>���g���5A[Q?�_�M�=*�!��a��ɠ�N,x^�ZN�h��L�^��?�`�~
���HS�F�҈�\:u�R	��"�s(�$mI�s�w�0��o�|���3X[ZQ�}�{m8�D.�d>����)`0s1��F�'��!)ܤ���ի���]��0YƂE�r~'��2�bҭG�qg�BM[ ��MlfI�H�T&�`(����F�-@�n�k�E�x�$#A\q�!��6�-C��ݹ��r��f<�b����5̜,#�*K�,�����JԃfSJ4�g�w����U��](c��B���={>��.�����w��?p��İ4���G�.�(��5d�.���jrx�W�Ъ���WD�:6��>Pp��ĳ�۲ӻ�F��� MӔ9��Aj[�_��J�g�ZZ��!{�:��6?{�%�-�>�D�z�Ք0c�-�qS�kݧ����y��S��`;ȍ�VR��k�--��T�F�@ �Dˋ'��z����մ�x@��ޅ�=�ᡏ���X[(����v��X*�L������{j6L3g%5*��$���7�u�!�������7�.�d� ^m�{�t�ڇ5�3r-���f�>mD̀k�K�ӧ���|s��}�՟Қ�_"�������9� C4��Xl���\_XK�CGᣲ�����N.t.Cȫ�Y\�Bkn�V[�'N[��E*7 t�����ZUy`�����lI�s�<mڲ��v3�a�%^M+�Wb�����S�|��6p�u�����-4��q�*��Z�����(
ҁF��CRN��ӴAL��c���
j��Abt4�\&�V�T�E�8~F�H�m;0�{?"�h���΍��A2�!�=��	�/�?���
M�A@z��y|u�Opm��-������0y��͞�ܩQ/Z^�ѩزk���
fΟ�WZF�Q5�6���j�C�$�.�QV��Yp���\*M�zmϹ���"}Y����q�U�;���a���Z���?S��A����l}[����(@nϲ8C�
��*�ia&	�g�    IDAT�3m�	Yv�����)��G繁�!M���߃�y�N�~��� �cFcfQH�$N�����:��������p��t��:���T���|R�LwU�̨�SK���81�ĝ�-� �;e�B�24�爚�C7��OJ��k�1;���A�F�RU q�b��I��7��m:�&��8A��>�����u~v�N�Bse����#��؊��%X%-�h7��>���{�L�U��Xa�r�>�EN�&Z�"��\�����Wq��h�.jbb~m(� �7�@�A��.��F*���"��"��ayu	�EqI��F����zM��i=�F[�(q����"���!3E`�3��!�z9=M�v��C��ܓ��{���5��3�q���)���cǯ�+Mۨ63*��3���B4�4����f�h����$RH&��!���kuQk6�P�)\F���Z|�� �.Z�Ō3#���@!cp��^K�D�1��~�7!�������S� s��l͠ѽĆ#��Cn/dqPKm�(�ZbCOM��\(`�7�����WÆǇ|�/�דͦt�f��9��j2�n���=M��gn�2�p4y�U�냽�e�f�T�n$i��3��6�&'6<��I�G����W�Dɞ2��5�����1V�6Q(���d��[�]�H�{P�ݫ7P�_����X[���/�Da�4�v�D4����D�v�cF�pÙ�ن�Q7��1�$k&��<˨�7�Pcf0]F�|�U�t��4L�g���,����f͠"p�=$�dј'�n���kq�ĉ�R'�����j�e���Q/�X+�Z."�Ib���رs�fgO�����k��t+���8��M"5R@_������I�������Aڍ
����0�k�&�{� '@ؿ�~�F��Q�G5�	��t����o���2���}B�<�?���v��r�3)��K��ޟcl���>�i8�w�Պ�X���f6=2�z����}/~t����h���HS���V�/L��q��}��6�\>�V(���-��sh�R���+�z�N�|搎g�sH��e}5�V^����\��k��p��p�C�YA���ji�z}��v��d,�u������N+��1[,�-J �@ntv]pC�:�NV�k�A���F���bG�η�W��s�Ry����!g0"*)^t`�q5)A<��+N�	�M#�pQ�Ub���.%��b Hsa>AHDċ�b�r�B��R�	��P(� 53AZٮ��˳X[d���V���P��!;4�l&���e̟<��yR8~#3:���҅m�u�II�EѤ�FNXE���d���H�[qHدj���b��_��s˿6����M��f�M��D�}�G+�d�e�9B�M��V�^�B����z4;�7O>����eʹ�P�,������VY�d0�#�Z�������:^GFrxc��A��D���q��R�z��s����G$�'#�gϣ�&7a�,z��	*�v��uS(]+�D����(�"=�K�,�Z�4'�4R���wySK�E��<4,T�ܥ��,f">Z'4�	 ���[[�������"6f�1;��H���} 3���:x�a,��3\�'�(�B�I�x`�昅�QUYR|l�b�?��&s~�1	 ��P_����chV�Ф�0��]{0�c����M�=��:BZ��!L7�,D	m�zѓ��l
��0z�:E�*��S��Bki횉2��nC�˦��FVo���-?b�MT�p�a3����?�!�=�w�M)�i�}Ά�lI{T� g�ƞP�7�n�I�Q�@E�	"��~mM�<s�9Q��~� �����(��D6�E�F� �H��ЗW��R�3)MX�3&����h	9�6�Q7j���I��G�����ѥ�B�c0;C����R?ӦaH�iRY�
s�0�&$�I���d�V�dN�<��.�;��W��Dyi	kg������ѥ�\��@��>6��8��㎁m��m�AY�f�:s\��}������8���u��ċ�'���1"�ޭxB�ە��K�b���Q��F���V�`��QT�G(�G<�W/#ԍbth#7��r:�E*�B�FO�(
[EW�Qc�iauy��O#�h`0=�d8���9fQC���CN9���)+>���v/��r�n ���Э�U�}"��@v�DZ�3�#:n3׫\^F:G2�Z����3^�Ӥ&�d*�&�t��䤥���r�h���{��6�P��G���dqi��V'���	��u�b��u�ϖ\y��Oh�i���� T8 �IB�{�"Ȏ�	������XK�?m�c�M�n(�\?s����)�]7���`�I�FM�NwV�;b�>`3$�TǞ���?�	���`��7�:W�nhX�A7`�x�bk�%�9�A�3��s��_��͟�{ܞ�:�i�����ȋ���.��.�N��E�v���Z�8��׷�w��2뵉��F*�ҀB���a���D�q�Ԓ�̨�{��YZ�W���Pر�S;�,��(g�?�{��?i���(w�@c��<4���Z��4u��k�Uƛ0[��˒{�I�AM���b4Q�o�yrc2H��x6m�>ksJ��HCW.����I@"��i"�X-cmik+E�D�� ��c��}عk��,O�<�rqU��+s�y{߶M��� � 4:�[Ʋ��8�� H�\^Z���,I)������]�c�ݏ�Sg1s�4���X<{Cc�(M �F�΢ʍ�d%�
!�� ��!ʌo �G��������<��[�P̊�Z���c�6\{��}rzfL�	C�q�,TJ��w����TVZXZXF$Pr�@?Vb��e�v$��~O���F�"�B�������&�4�#��Qk��A��u�؆"�_n�e���g�Gsc�~��^+�^�Gue�vC����,v�cd0��B�i0�tѕb	�O��g>���:�$��!tC	NLa���Ȏ��K�>S�n28����{�U����>݁��S�3H��Q8JӶ��WC��
�QEc��6�0.sK��s�a/ō�y$����F�Z7���~��~��,���X�j3�h�v���\l��AjLD�%Q�h���F��%��̢1��C(62���v�ݯ����"ә��M$)�cӻD��0���_ h��DIY �
;��C��ʊޕ��k4���ulnIS�k�5'n���Van4w�A;����4'���}t����<��]{�A�0
������C����8=�z3��r�`��Օ詜sU����AqFIH�(�:-��^�~Ƃ�b����~���^/�Gxۀ1F ����$�cD�4J���ӹ��+��޹������a�O�tw���{�=��."���Y0*r1�B,�F��D�&4���yI�l�����FGF��(�I$�կG�mZZ[I������>)_n���be��i�[,ֳ`DA�V8]�H�2Qu2��c-����|�j�����a�$��=T+�]�o��C�-]I�L�E��4>&Pu+�׍��y<���#�0M�|k�"��FFlr�.<��]f�*k;�
՟��@��,|�A�>���4�ʩ��J����f�8����Z.`ca+��./�z�����$���h�P-
e$`�%�^�(��
!�8cI�Ζ��sAR�C���2�h�҇ߡ��Y*ǚW�_k������5�[��S1���F�LQ6��¥�BM"=N&��gJa�U�}j���a�,��k���*��T'6�*v��Ux��<)��4��CF���-vR�@�j�Na66�2�Aza1�G�YC*��Ğ�����ŷ��:�/ s�~ƹ��q��Q�V�w��&R%���׍|��z����$:m�5�J��Jp��E�"�0��,�n/ɔ���K�T�mq>2O)UN1�ZQ:�L��J�2�&v���B�@S��Dh�R����4*�<�����g<=�Z��j�#Ub*��kU�c%R	�z���PX
���wMa#��s��Ir��Gpy9��=��Zʜ7��H%8��fѩ����QF�QZR<�D6_@����Y�+BW����\hU�pw;Hi��[�ϋr����}NQ�>(4����#�j~qY*�G�=�@���"�pW�|빦xK���-\F4Ñk`yeKsH����m5��F02m�Z��vm��ب��g��l�
)�2+�@���N� E�*�������p~.����W������R�fw��.��d������2ۨj�R�ʻAUz��!�X�ầ������� �v�O��KL���	���|�QA�J��A�bwel+�sqd;i����R`����K��C�(`�1@���nr\�
�H��{W�S�x�7��.3�W{����5�"�7��mN`?w@+׶��C
aBQ�`L{�����[|6y
i.fNRv�pm�X�
!�(�C7���=���E��.Tpvn�8Yp���b.�&I�	�G8^A�/���n��<���Y�/I��sI��.Z���S;L{VE^+N�4Q�?�DY��H5�L�Z�`�߳�ʱ�`�s�J��:6�VPXˢV*�ƨ7�$)��r���g�]ˢ�h�Y���B2���C��F��T�K���)����d�p�A��!~���%����_�2�võ����ǥs�𸰱��z� /u�y��JUE`��J9�z�����GG!��ĂN���Dw�tF�	����`v�>A�hY��F~Tzm�:sg�\F~��|./�jͶ�SQ���l,(�G��r�'m��G(���]�� 5��H�F�f�W���8
dfU<�v�͵.	&�e-ث��� R��s�e4
k�f��&31��� �ݷ�S�B�%SK�CR�Y�������#�½_{O<w��8����R����q���Q��z���}5Q��Zp�_�[��7��ǅp��fHZ�0�&�̌�%8��d{�^F��C5����:u*VxT$��ʊ>��/6�/�/���.��f$��H�L�!Q��+�T�H3�
hh�fA�$n�hjWL�����u׃�u2��Q�b�����Ю���"QL��-�q�Ǎ���X>^ٲ�$��1�S�Q������2�V�JR/�*,bg�{ہCdx��OA�y 7N]m��h���[�f�/�� x��=�_o��C��X�*����b*��`s�Y��4]�J�<V�/���"�X�F2��)$�	5	�Hb�Vڎ� dk'�Y����*�^.�|�B'��\�χpE�E eݛu�}lw�qa��=���8��),_�_<�p�<w��J�3�굺T���[yi�����v�A���M#�3O��!pb��SbV��Z���:*�<�1Q/��O����M>�O(|��s-bF�Cs�Wn��+�̪:�)I�ת�8��0��F��yⵅy,_�B
)��H�X\��@�]Sz��]=%��=�}ؾ��:�g9�Z3|��\�l�>���~>��jG
��D�g���]d���Bc3B�R%�ד�q�n:�bY9�΀���l��������2R@9�C��f�P�x�^��x�/�� ��]N������d{׋�DCȌ$%qO�#Ȥ�(U�����A��`�]�յ5�6���Ql�����R�v"�N���1�d�hĬkn����ښy�ZN3�Z���̴\�z1qJ&�ɤ06�A Ȏ)�Ĵ,<��y<���h7[� �
9��.��I�*�,/J�����8z��כ�������Z����q��)�߻K���D�ef���e���Ezd�F2��/���bE@N(q����~� ��&Ĩyqi�x�Zs��8x�0f����}����'uyuA��#�Q�
U<��7q��)�"A�b1Q1�>�Eo��ϡ��N��~�]Y��f|dTfz~�����@�<��|��k�J�.����3����2��Da��|�p�q����O�Bv<�B D.�C�V�"����>�L*%�u0��znKKK2k����g�y
��OU^ҵ�9��$"�(FGG�{zG������g>����\~�s���W��2�3	4�Zy1 G��J�Wv��s8H�Hg���V�V���Ba��̫J�&"^F	�2�̰�O��ʐ1P�3�ë� �v),k�կ���M���YO�2��E"��Z�^���~��.���u�b�@6E:=����)h	�z3��fs�����Bm>Slg�g�rӥ5�Y�����dMܐ��V��T��'2��=_,%,�V��3_i�b ��	���$S���%^3�gy'}WY������D1�� i��VT�I�y�i1E29I)�Fr
;�o�ޒ��P�U��rB�i� �p̦����"��,��2�./}24���kbrzB:�K��]\E>�.�p�`��"K c�Da����#i���^�ɲX�A���fv�2��,<�"^���p������~��sֳR��\���~T:!m��c�h��/��\�K�Ǣ4YdA����86����р_���� rϡ#���FrVT�ZbH��Q*��@����)��
�,>�K"H���m���+@���B���3��hgQ0�Po#_k��q����"��'j���k��
��0��m������\�\��9���+�U
�,���,��d7]w 7��X<w�-zRڒ�#p�Z P/U+��o�>�0N���#�D��A����#�11s^_H�o$�rA�W����ky��t*�U6]h���q�T�i��mU�[����
:��uxHh�$I����H
LdSII�<w˫4���	"Abf	�nm�|�[�a�M㰪r�eH�Gx�e}�X���m]x�i,QX\D~i	�rY }0Ef�4F��dQȭ� ���
����0B�$S�dF���Qn�Q#i�i�Wf �$����əM�>�4\
�8f��0����(qU����W{c�������ѡ����L{\i�Љ�$�9cR�.���.�s�X�p��U�`&m��U)r�T����ۯN�:�FF��[0=X�w<���3��I��Ee�n{��u�]�@�/���sX^XB�J�/��Q+#��s0&�����,���D8���4��߅�I�;}O�|���ᛘ��ރ�Ǩ{DYA���S�WV�Z���	�t�6�H�9���	���!�CU����^7��"J�,�W�Q��Х"g3��(����AB6$��̬-���f|���X��_�RkЎ�>�50�I;V�M�a�_�-C�kh����_m�ف����S.���>���)-S�Ep��
���w�o������x��R<+�Bͣ�vj�r+r�ɸ|��䄀�b�(3��w^���
9�#,��E�Q9�R��k����)��i��e���(]A��"�8����l4Q�5��M�m�VA�U��qbrL����~���.��"�����s�&9bP)��Ay  	rx�����d
�����r�"�A�*�R��u��b]-��P��Z�'��%�'�;�LeP�Tú]�v�Σ�<����Q��|Q�Y0�lV�>	�I9�x9{�B�x\⠫��ٳg���ʌr(�䊀���	�-�I^�g���'"1Y�Ȳ���JUp�3s��ք�Ñ �oQz�ǵ�
ح
����r�,,,�������V9,�J��t9�tS|F�8IY��(�orr�|9�*%�}��Z�!�W�Q��"������/<��������(\���2c��-�)�$ð}Z� ���w|X9N �����l��ƹaP"L"u�~1��_�����F�r-���Mk��F���Ub�e� ��҈�]��a�'kە߳�X����("����Q�-���F`ŰY���_T�v<��Ze�V棵��Q�7�)���k�}��x�"��=bQ(����HICB�
*�J�����ߋ'�ᣐ��3h���<�ʬH�� [c4���h��~��E�;cT.�p��S�3�����s����,    IDAT:����ҫ#7��U,�=#��6����{�1���ŋ��Xˡ]mbmyM�o��A�:tZ�pT��i�Ҧ��E}29��n��z��l�,�Y��U����3#q<�E���f���ڲ��<�|�� 9�����t�Z���Y��h�ĩ��R'�ߛ��C{�n��X���ݳ��0�w��(�Z���j�̋z�&�qwϏv��]E7�duԊ9�<�Mr���5�hTIg�7m>t�a�M��^��5���<����Fe���~����X�:PsE��&�t����>ŀ��m����5I�:�R=�v.^ƾ���f�|�^D|]4UD���W�w-����aq��wZx�O��9<;�of�z�@ߌtz�P�x�ģ;����m��׿_��ۉp4
��AJ� �����&�r[�f��E�.��(���W/�W���x��ǉ��u���XJ����VVWq���8����x~�����/�F�@�CF>%ν� ��v�"AZ��#_8�3�MCr��kK����bk�R���L%1>5���1	��\N��+k��v!42���3c�;�(7h0O�>J�õ�Ii���d�]"�C<��!ˡ����{Sۦ���(�
Î+���y�P�~8��
Y1VC�P*c�ى�Qf]�C�A���ղY�.��[G�TR�GYM5���F����l�ȶ�h)��UF�D��$e����ϒ �l/���4��?�k
��
�//��+������}�P3��M �F�LT	UU]J�����`$�D*���T*�ܡ"S�1��3i��N)�Z,af-��L]� Gf��9!�E�m� �v�����(dY-\@9��.�&����9���ô״|��@������C{o�y��m�i��5�����U�^x@&{�	��M�����/s���j��Ch��:D2L�6�rv�yQ,���x<����_�5���=��+x橓�=%�C:��&�s��&NN���YԢ�#3H���R���5h��7Be8�����O�逛��PPfO�1'H��t�(���K� x�k�#4�9��vi�Bt( �<��&n;�x1_T	m�W:l��c�$�d��<���X~U!	�t���n-�i4��VK��$�B�f�T0���
��S�3�m*���XY�
gr�L���ɣ}��X(��-�a���_ 8��tﵥ��g�������q]W�� .W�$�Z�p(��]���B��}��\_]�����>���Sԥ�D0��{z�֛B�����Ϣ�(Ͻ�iVE��-R��Q�{���]���5��M���۵�l��M��9dʣ70;;�������K����5B�1Q
�t<�t�J$�?'���+]��^2b;�5��Y�`-�{��%�6�w��Y�F��,޴V�W�GB���i��Y;;��5T� ��}�4\Ò�d�aͨ����mk_�Y�(�%���Z{l�r��H��X#��$���y�5��JW.�2�+
��%[_���I�3t�_���I~V>}�C#ܷS9ݰ����}Q渃���Y~��(g�D�~з?_�SI+գc��ɡt�ם�K�7h���Q�~�C��x�qZ���{��-T7��Xb�o�RmZo�<8p��;�B����E��/�Z��]k	�039�]���ő���}V4�3��H�C�YG�RFaeY���u���v���D�_��7V��Z.�ya�	'b�%�R�c׮��㐖p�w��h���(����ㆽ���'�1�NW�<n{�+q��e�"��B��
Z�Rc1��>��Qx�!��^�v]����u��+�,x��(�@�"=>_$)�׭���$����DL���p�uy�q����k�p~������\�Ƞ剣L&�u����!�3g�S��Ӹ���F#.�%��Kn:��tH���&�p�e)�v� A*���o������7���ٿ�3�F�D��Ǿ�'�NO"��:�pH#����yE��~���D��f�>���v-l"��䀴�J��
�+��4J{H��[+b:�K_�b��U/š���N&DH��ɕ�5\�����>�z��8��y �Dj�!�GfP�r�Zg���^��J��Q���d�Ig�-�d��!��B��(�,��ϫ9o<���i�OO�1�_\�ʥy4�%QD���Fr�>x4l����4{�}"C���7�o�2K1{�g]��+��;+2��^��:���A^x�,5YK��P�C����HL;;h��� �/]�10_u��ZV�I<�L��""�&�6U�wF�Z���*�Ծ^�K��1Tq��6���sn��TU���K�Б��/T����P�ip��ij[�~澓7!�{
�H�B)�0iUP��M 22���b�q�*���A���T�9QO��_j7o����@�k#���z��6��� y������N����d��M�<�mES�&��}[�����*8T��Ϋ	8ɭg�W埦:'ל�0�KMk�ܙΧ,�v�ɬa���������a��PV-����0�\~�. �����b,��>򿱺�?E�^#a1�g�A�R�(�td�F��:m�|L0��A~?�=�A�hQ�)�+�]T+U����mYi$(�l!)S��d�H������ҡ��S��)�pIi��E8I�[�B��C�#fόHE��B�е�|h����c����rϱTA
U��ϋL&%j��xB�J�|�JU�"�)HW�!�H�����̫�[���=��r�������"M�yQ̆����D��!Vy�A���\�`�tT&jT�~���j!��4*q��}J0�Ϡ�N(�(�pS
R\���ɼ��0{=����z��cIC!YshV̍�Zr�QE�V����ו}��b��o�]���e|���=���5�v�Fϳ��r�.^w�R���Nb���H���F�	���� ES�!Oe6u��T��hwE*l� f�$� f���l����ڧx��²"|�(y5b�*������m�RS���Nr�R��Y∔�dz;�,wd��Kb��B.6wE��?�8�wC}Z�wH"���qq0�
9�ܓD旡���F\���6Fl�b���}T��>f�2��Oa,�dF�=�
��-ŀ�@�����ib��Q�mp�Q��ba�0�F���B�MKv�c QY��7�p������U�0�/�:�` ��g�a}-'�|�|IXKӻ0�oB����&-�k=ǟ(�bf[͕#�"���D��f����6��*��kWp��ØJ+,�-�%}��.aupF9��ˌx8@$D����˗1?�9-�06t��Z>3�+o�1g��5���ʡXG�߀�ǎ�
(S��@��C���h" _�0��k'Gк�j���V�)��i�Q�m ��*qhtl
.��Vc��#�g
UQᦎ�{hE����B�D�C��ſ>��\̢䈡探��J���"oǩJ�<��~g1����"\�<n����_rGwGd��ө�O�vqw2�sc���-+O�D��Áǟ?�w��b��@`l
ْc㇑�LK����` ���*Ԫ�1��ߕ�`����3H���v�p?xma�b��&�uL���?�s���#8r`�T+(T��V�n4jm�W�~,����=����/���z��&��@�A����,�)���W�:X�{�.����f����M��F!���r�.�a��±&v�BblL�҅\k/���@��m0���nħ� ���M�����'�@7b`�*桋���B?������Vp��2m
�/D��:MԂ��_�\�`�Nu�sS&P4����i�p�b�X��Z�Jş��	%Uظ��i�,�~H�ܟ�R3W���ق�~�>T��Ob 5t�D��������v3����3���]@��� �\	C H�[����=&v�WQ{d��QU�V��(R���G�B}i��H�>�0r�v[�s��z\6��m+��#h@��P�u9[���;�����h5�)(ѥ���	�����K�����̞�C1���5p�iҢ��SW�~���ϴ��_�&������ ���$��of@D}Onm�]v��\{�0�-��$�g2f|Z�y��3g�����Nv��B%�
?f��3�=�`��6����Eݖ�C�2���P}Դ�?;jN�xQ��
͍����U,Į�G>S<D��N#��ˢڧT8����/ʱ���}yΦ���%�p�i���Z�..v!��h6ZX��'�X�h�O�����tO=&�r	��؜R�	ިV�F*��1 ^k++��j�s���D"rfWs��y>:��M�Ú��A�א �v�ץ:Z�A����(���B(�k�ń���`,�cN�B,��3x�rY�n�$���X�����"����U�$ ��v�Sp��_��P0�� ���'��:�N�PGC��$�����S9.�Tf�v�rY��؏�o�	���7q�Գr<�#)x	�9�<����'�2�,8�D���#�o��?���46j�G2`�9�s�C�I�!�:v�U@IE�xK���>Y;=lgHV�q�ኈ�3�d�J����:ρ�G��l�<���Rk�a��h��c0�qÂ�yљ���H�m�x�v�y���j�Tq�1{���$���	�f<bGҮ�:�fU�M=Kf�w�������P�MI��Hf�����G
���(��{e��;�eD��3�K;rjt~\0-�x����W�w8F��7� ~mg�*M�*�)T���=t(����zťe4��(��U�R �>���5�3���eԋU�T�w`lj
{F(C��@��h���YG�sJW�--��ێ �#3]��VA)����yTr��w�8~l�G�x�/ ϙAgOf��)�v��#D-ΰ�Ҙ��]����p�V�V���a!���n#Q^y˵�;� JE8�U�I|ц+�F|,��]38r�Q�2I���
�~�h���3�����ԅ��[s�P��#��Y(�k�T���0�Q���� rhVDuZ6�<hu7X��]Q��;1�Vp�rz?u	k� �^�U���(��p3�a��Vŕy��]�}��x���	2���4@��@�r��\�zFl�����˅3�xߟ~�y�4FC��/0�Lf�$��>) �3��`K]�
o��M`P:�TR�,��C��UC�$?��Ұ��ELd�x��^����?��ߍ�_}�h/�=&E�;�Bȹ�/����G��O�-ΜY@j�'��	��h��T�B9�����ܾ����j�bx�<v;}�.<��(瑛��v��Z� �$���)�GG�n��avM�z;�.��(�#HO�B(�F�Z�q;�x
jW��/_m��r��FIy}�+}���L����-�/���@�����n.VZ|�Ψ1n�řCֺ�BL$h:Z0�sߡS˾�񴊍6�+�tc�a��a��q5P��s�_���P�<ʌN�F�B5�AvT|������D���}�PǺXl���"� I �C�Y��Ln8��
ल-�/�z[9���*fJ�d����2��̾��6��`J�C�HZ�P��l\^{�8��Ū��[��I���k����.�yO�7�N��Є�d$2iAJ�ێ�a�Sv�*�D1�M1�`�6P�84)�n�ږ�G�o���+<��"-3�z3
[�O�%��I�K�>1��6-���M*n�FE(��

��Ԋ���](�x�P�"��\{u&�]*�U$��L!Ĝ�>s���zr�C:�����fʀK�e6oem�lV �P�@m\��3�<-�+A��o��n}�(����uM���D"�={fq��y,�-���(@���X!x���t�a7M�i�",��S6;;�J���g�H W��S�g�&ۺ{v� @��a$ �6q?FGGX]�tY,c����^J7�������p;$��5���?2� G��yz�ژ�M9������:99)��k���9@n�x��v��%�;{�����	=����Ȥ3������vq{��W��� !��Ç!���;��7A6��/'����H��!�x�<V�v��0�o�~ͫ��o?�'�x\�}��Q;[�J5�F�},���lu��m�߽� Z.nz�K����Sg��E ���GS��*j��*n$\�A�3QM'��M[5�I��n;MP�mc��3�J�&9�ԶHh��=m��r�������a0hfra�q�>�� +�}J����#�r�k�6FW�hy�XwlMˌ(3F�R��Ԭr�N@Lr��h���	���]��?�#���,��'bC���s�b�t -�B�d������}��b�U{��V��k-���8�f�����!v���Z0��9?M�9*��ϮY���]�Cym�,�y=�}� �:(����X�4�F�*�d�06=����'Pm�P�ǲ׋�r��d�n��9�(� ���ؑ��m�P+l �<����������^�L���2J+�\R��I�7'��y��(a*O��s���Q����
�d��spT7�ûq��}��
�S�Mt:U�l,��w����q��ƣ�h� �b��3;�j�����������?>�g�@�^��8��tW��Dc����&P����ۣD� S� gځ4*��}z�zn�^� '2��j��C��>o,ܺ�j�%�˄�S/�����eaV<�ٸr�%�vqF�����Ч-�d��Q�_��������kPC�n��4R��Pt�� 0�O��N��7�~�K H�d$�������qa��0hva��U��n�8�Y��u/��}�/bb4#6i��(�ĆɆxJ	O}��wσ3s����}��� ����aDR�h��K#GN�+�U}q�V$;+c ӥ�"�<�
�2�����kÃ��06*R��-ΣQ�-'�J#51.����be�����tk���#��`|�d
M��bB�pTjCN��v���ۗ"���m[�� (�n��z����^m1�zeO+�YG���=�ω�V�� u�3�a`B�!��$٠���K�{fE;/L"�����;�A34nY��-�Nb0٦�d=���J@aqj��6.ޢɪ%��b5E*M�j&�1bL&��N��)�k�-���S�W����`�*YM�2^�p���@"��ꞌV�LHEu�`�Ɍ�Ii���C�:Lt��'A}u84/�+Kt�pmZ� xo�՟gp��M���b�� �l���|�{�ٜ��n��4��u҇����M�(��=�8��<d����RVۤI����C,F�͊TD;�T7�Ѯn�ժ�۬Մ�/H��ٽS3˴0X��z���t�x�:|XLş8�$
�uD�	$�q�9�<�H�w�F4G�����*Ξ;�R� f����{D$�{��*���
��k�.d4���v��B:�	�H��H%Sؿ?N�9�3ϟFm8��%��I&2���[�s�(Xs���\��H�D�����&xj������t�
cdt��r! �O@�8� ��F<�T�$�x�<ʥ�t�R�$|�^w��H�GDY3�]��?�4X���!��sXZ�,���䌜}v�]SSS���A%����JE�8)��ߝ;{V(C�n������ۇ'n�m�5��������`v����T���tFF0(���L~���F��޽�B�=��l;��/wg������./I���K�rr�bw2��`$�Y� "���V07� ��P,�c7�H��g/#3s o�Y��B�e����v��3dC�m���'.R�(��\CV+���13(����.A"05���w��[m�4�b��_�Bm��:W�׷����F�v����U��j�����`ʪl[�fU��C0�s��|�6pT
���^��J�̐-����ϠG���}�^�w��5�ʼn$wa��G��I�šr���W<� �Ki�B8|�����Z5�Wq�YX��va2�|2�׫ʈ�[��ԧ    IDAT��_��^�ᐨ��=x>�ss�0w���"Z՚��e�����d%R��m�"�d@2IppNPt�t��]�x�H)��m�])	\8�|��;<������G�YA4����"����N*|KT�y��Mno �hɑ1�GGU���B:���Du�2R�6F�D�=D]��=��^^�+��-��{�;&�w���^"� ��:j�6�U7�QQ��z�[��������翆z�����Ѩ��
{�W
w�u��r�L��S·6FhGB��=�i Uwk�0���e�`���'��'������N�����Y ��hVpx"����v̦]���)�e�M4�f�Y�6�a�	3�R�z���'��)�{���b�� ���ۈ�0vS]:�#�U`��7�N����r D�@Dr�F]MR�N��_����ex��kW60;������e��@��<���t]�;���(��C���s��`km�+�~�w�'V�[����#p"���u��a�ܱ�?t��Z�-w��mb,�8==D.sKX��C~yQ�VOcq�ܳK���6WQ\Yc�"<�p�>�{�l��̿x���V	z�4H�@��p���׶&��	�eI�vّ���;,�����u��ް4��_t���N[��Rq�eP���}��A3���1�+V�H����S&>MB%Tz�$�\<Y�3&��l�%���	v�����F�3c.z������R��V ��%Ҋ9�0$�`5��R0m �qT�y���6E�|��ʹ��I%��A�^�]#���-M�ҡ�b�⋬�8 ���ϯJ6�M��8t5IgP�#�$
rp��o|�Or�A���<�����C:#2�*̭E&{������}�KQ��I�xVl�7�l/e����L�B���� !@޿�[+�v}�?�׾-��\��F@F_� *�B�T*�X��)z%������kp��pu+��
G�[O���w��1�ٻWd�9��̗���( � �V�cbbB:�Ϝ<)�RiU ��>���+�#Q1�͗J8�� .vR
�u��>$���ϢZ�];���5�p`jz���Ԍ��ml��饋���!� /u�HM\�ʽI(�j��H7�x+��&�P�ѤIz��XYl�ӹ�]��3g�S��%��4��&�q��q1|�XϣM�BQ�Ov�UՏ˗.�Q���4�x�BIb���NLNNam5':|��S�4//�p@�'nK.��˅T<-kW�T�s�ss��1��rv����î�AH�"��V*X�|I*�����KWi��tǎ]#��j�& �����E�J������u��E٦щ	��m,.,Hb����n������Ӄ� ���h,�����΢R�!C�t:d�s||S33�����H�3X^^���sp�<�%3�=r-���8��g4�"�<a�[u�-�	�.؇�};HU���λY#]�66k	�<e�Z/1ʤY��1i����Ƒ��(���Τ���I�J&3`g0�Y�� �v�A l����*i�r����^��J��+Y���t�d�v��:�ۥ �����z�������bφ�!J�I�vĺ|��&3QRݞ����J���!)�p��%W���}�ܢE-�؂R�Z"$�1�1q���#!�s�]%�E~e��K��*W�'0{�� 2�Y]^��<��Ve��R�صw��Q�=T(��r�w0Go4���������B�y��t�k��!����+���S�6�8vxGg'�퇿.�*���Գ�cy9��'G[� 0E4�e.7\�&v���z��D(�W�yn��(ܝ2�/>����(����@��B,�F�[�'�Ǎ/�o:!~�y�\���������;�������/��������6�.���-@��SgQZ]���#���+��x�� �>���F�-�:��F��%q���7N^�ӹ��ֻ����F�4�Y�>����d���w߅}i��Y�dQ����W�<Qs1P@o͞}r=��v�<r�~��|uD�jG�LM!��b'���~T8��1z�o�<�x��qm0�����6jT<+��P�w��Vq���V���c�0z���IJ(�M�%����GV�0sȼ���S����x��O 0�3�E(1�b���Q��]	�mZ���#@4tM��b�W$Z�����l���[G�D��E�WVС�.��!�g&�J������ŋ��gUe��������L����b���#�1M"�a���	��sV�7���%]����v��.�W��%�JgRy{�|�T!t�_?ߪ|���`���I��ZIH�N*rm�s(�3%Sh]W+�g�?D�ͨm� ��s?����J�W�
^�3���$}j�vqt�Aoh��
�hW���#�c�ㅊ�r	��b�KZ$�]�����qQ�ރFK�+�zK�����y�C��� o���?�J5��s����E�z6����K�Rn��bK�C�IE�퓉����-�i6w�KTלm��}�m+�;���?0���}�֎��������3(�t#vdA����$*lka�>������Y,�uU����aog��D�NUh�.��5�|^��a�?xD��i���Fvy1� �#5���N�Ξ��Ν��z"��`��+T���C�q����X*tf�Ź�.˜�=��o��	�ņ`jj7�ԿiC���.\���8�;X���"~�A���g���ؤ ��슀Tv�HO��a*=�BXZ^���$0�@P�*e�޵�tJ�6M�Y%��=UCy<�JI�$��C+�@@�jKJ� ���,���}��(F�_zRMt��%�M��N�������������y�k�����o|�J��HA	ٶ�,^8/]�H2. �@�sD��N�ލ��]"�C��w|���c���|��y�w'��`��?��#Q��G����<� �h��Ǎx<��'G��1��(搴 ��� �jƍ��rRzYw�}d�^�E�/�P�0�7
�',3���3�6I�`n���޼�����1P�VȉJ&vMą���X#��t�K5X�uR�JC��&-�h���%�3V����E�(3s���/��bz����� I�,����-�Y0�Hb�Qv��">#A>A����6����g4��H|��/�nӄ����ߢq��\��{� ��B�4{oޫZ�/۟7��P����m��~�s�Qj�u�m�R�~�,4��0l��c��sb���}"V�1�Gam��eѰE��}����/��籺�$Z�q���ٍ��8�c#pz��3��@�@O5r���`�e/:dj5U��yG�ZM8)�D���5\:�4����`v"�'��(a/��	<��3��� ؇v��z�,kZ d�7�ѩ��,-!	㿼�m��7ߍTԃ˧�g>�!�/\�d"_������\7���O�@/��F���%̝;�jى��Q�Gv�������"�^���V��A���7��w������������)��_#ݳ��@4C�R�ŋg�ȹo�^�'���D���p���W�{
��]T���u����#Ζ=��,�����h=8�%���;�0x�L.*�;9*�;���"�7ޠv�!^)u���c'���<��x���Y����Ș�3�Y�K�D���u�TM�����ub%сV��/4Q)/#�t�R��Oښ!G��gނ�������-ȗ�2�v��UL��yE1J����r��R���G?�w��'01{��9�It����h��m��o�p[�Z^��.m�{V�J��M����s��ĵ\@~a��%����BA��f06>)�rސk��*�6:���S{��u���.j͖V� ��?QҐ�A=S�瀞��G9�7(�������R&�8Si�nfA�^+-�����A�?]B���!����)(T��g�LB�m����t�1ɸ�Ac�n��`f�U�a�a��@Ut0��h�\�+�#P�����#0�c)S����ܼ:���=Hp��� x���	��GŃ�V,��Y����
���y�H ��%� Z�P�l	�ۜG��r�KN�1n7�]�4� 1R�CA��~IB(��"l(��R�����xi�s����W��4*�4�w�e���+��8�~�w-���r�R�51T�'��2��6)���wf^��F:�T�l�en��_C�V@��C9��veN*E�HcU�8�6_����|���26V���e�W���� ��>��=����8/�}W�����z>rU��ԻXX\��*~>O��� 2��>�ܳb;��y���8��	LMNcv� Μ�$��ބ*�R�B�*�r쀭-,���"�&M�+��3�{�[^$ �ԩ�d��&�h*�4� ե�EQ�����K���LOᵯ{-������p����!Z#�L�ʇ�v���g$�q��1��O�|>�M�X\X��?.��z�*�T�Tț� o �d4!�ORty�&�������e��|�}���{�y/S�sffF�䧞:�@8�熢R�g�_'����-o�[��Bw}�'��/�+�QRv	�4?��ȶ3�R��v,������&����_�|_��A�^3�8Ξ9��ښ�d
�TkR��q�129#�p$.]�|��/(�*���k���ރxvn���H���J>O�����'������[`�]�籱,�NH�R*ӆ|g��0��DMtP��-_�������(�-��ڂ�yu<@��I��j�Vf�r����;B&��;� 6�Q��_7��ij�#B�&v�?��w�N:�qZ-�_����4�(��[P�3����k�ag���+�l��]sѠx��*�U�>®�;��6ڭ�y�j}���
��~�3{ .:�K�QG��M�{(N3�P�1�Z{$ep�rK�(ndQ-��Rʋ'����{���F���bmy%
�����0Ñ�H��M
&I�Z�mQ=�q�_}�4f0(��_��'��i�%�C�ڕ�>�zv	3����8���HE�M���s�`yiY�Gr<�n����U�G�+x|!�I #�R*a�����ފW�y;�:.�z��؟���L:��������O��kn�	Ӈ�!>�T;�S���#HM^�\������g>��X/pF�#]na��"q�����_|������>�W����~�q,,^�~�n�>��O=��}�S���[q�^�b;?���8�n|�_�Ņ������E�*t��3��t��I0�[�Lԍ��[p�@^쩋����o�*O��x��e���r��Z���~��_!4���4V׺ۃ��1��,���"
���]]U�FRRy���� �6�N���Wω� %Y;�"��!���"~���1"Y�AJ��
��_��T+""�tK�c-_�������#�Bf� bc3h9<谽�t���p27�I�`�j47�o5�����eh!a;h9�ht�o<N��E�����T�9��U��d��id�2p:;ȭ�c��YT�s�z�;�Ddr2���K�DB�������})j����c�9�l"�n]�IٹB'���ܺ��px����͋Ӡf�Gr۶���pm^�n��6��� 4�Q�E\��fA��̶lZˇP(�3nB˶G[�ukӟ%�y��h~�߲}&�.��꿩����f�0�a�� ��V3QuKg��V��AQ�-=�,�V\Fο��J�Aoӫьe����K+�B�u}�Z��-"
Ξ���Pt�E2��S��m&�n�7���ei6/t����N4h{֙�S�,��_��ue�B᪥��"�`��-�H�O�g��c�b(�<�"pcA��C��D:M�iV���&�Q����
����"!Z���{�����v�ӣx������~ �>��$��sD@B`��G�d$�	8#5�*����_�/�����O<�O}�Sx���/L!����u���Sb)A@ş�A��ܵ�o�=���p��MXZ\�?��x��j&L������gO�� �K@�T˒D��cx׻�+~�'��P�������L��m'=��#�<�ĘP8(�&%�c�#x׻ޅ׿��blOJ�?�A|�;ߑ��mJ��2W���ss"��D��p�� ^�җ�C� ������W���?�I�H2�����7\/ ��o="��x$&3x�|�Cw�-��=�}/^t�-h6����>�O��rn�zf�w�y�Tӿ����r����݋��~�*UL���{���?�SRpx�G�����lN���ٻw=�,��iB"V"S?#�^��W�w�{v�������'>�/}�˲�33�8~��8w�y|����D�׋6��� ���7܄7��M���-갏}�x�o��uc��cٻ�V��t�f�tT���H��l����@�g�������P��-ǵ�ʭ"
��<���$���U3�~(���K�>>�Y�e�-�Jn�a
��~��z�� #0=��ظ=9�k�� ��an��;}L�';��y�F�������&5�-�_�ym����>�n�� �R��8��Am�����(GԆԦ������l-�kU��f$j�,1��0�>��1s��=���j5���_<<��A�/MO�f�y��`P��eI0��.<�T�d�ח����#+�ޫT䯊:w�^A�������#�q���g�9u+94��\,��wMab�DFF�B�&���V�I�p�2/���0�;hSW�PD��G�`�Zt��^<���%L�cH]x���!�aj|Ο���
\>'�ci8�]�׳j�#�+n��Qi�xC!�\]{�^�0���SZA�4���g4�Y��n��ND�Lv�q��u�ފ��Q�F���7[�;}�v ��n��Z	���%��o��Mڅ@���z�8=��ٍw��]x���ǧ?�q�߳��|�kx�����;n�����(^���׼�ne�X�y�Tv�k������
]:�#�F� ���P�a|oU��.b&��^|=n92� ;~��BN�YU2/.~�>�=4���\ۼ�����b~���~����_�ؑcp�Ɛ]�al|2��hЇ�����2�pB������ *��V��rspu��\��K�3�����ێ����yi  �Q��<��*"R�������b_�������}t�Q$��#91����6>i{꠺&�W�����������ea���*�#$P3f��v�nAΛг�P@ayŵU�y��ģH�݅ə	1�^�����˨m���+�@lj7����Gcpx�"�ߤo���24��2��-�]p���.2s��RY�2f@��3j�c:�;��Y0��yOK�ыz�ze*�;��:��e_�KA��l���B(�T*�b�y���7x_�t��ؙ�|[��4�jeQ$�v�x1�G�8��9���i���8��zA�(��\[�Y
�x��(1O����v1�Ԫ��~�Պ	����/�E����A�wW�jh##u|[��A��c������C���`��>a�=l��_��z�dGi��4�^%}�gs=1y�r]��ә��̅�]Bz��Πe5H%OEȘTkB��B% e��ЩPί��ĤZD�V@��g��^���EI������;����[1>9%�*��˿�'O�D,����u�]' �k_�����ށ�(#���o�����4���?u��S���N�RZ�&���Z�ٳ�<�O��xN�&Ďr)��܊���� 7�x.]\§��S���|V�G"���m�B�ar��cߑ�%X! d1���7�'�'p��Q�q����G���e��M
|�z뭲?��w������6U���53�w�����d���{���w��Wd���=���ŋ�>�<��)]z-�!j���o?�Q�-.,�_�����؉�q��5�1�{��E�
zպ�^��V���;��9����?=�x����M0�7��rL>�����色�}�Ӓ��u:q۝/���	m�*�?�~����:���p��A������=�x�q���    IDAT"�K&�b�p�P�y�׿���_�G���x��G>�����x����Ͼ���wp�}_�ٟT&�8�������|����?��q��㈄����}������n��v�9zN_^ƹ�58��=L��q��d�T���l�i`�:��1i#��
���B�bǙ	���l����Ͳ�*a��d�<�N>�}�f���D�)˨�!E^wr��}"�D��~�Y�m���n�`�{H���6��n-�q�8�>Xs��KICcz,�,3�#\�$�\s8f �`frp�OlL5TU���h�\�o�om#o��'�=��Yj�V#�?t;�iΛ=�&�6�	F���|��e������0��F�㯍�C�����qN��X���Ɉ	i�2g�baW�e���̈
�ۢ�J�\@�����Y8r�PΞ���˨��P����Frz3�!�N�립Ę�r��<k��.�.Vq\�r�v�u�k������:�37ꨮ������i�-|��_��U����d�8z�5*�<�˓&J���T��,4���#z�`z|�j~���SB��F��F��D���Ӕ8q�ݷO���\�B	O?�$
����|'O��zn]
��rUj;8\X\�ʨ���f�#�����̈O��J1��7^��V�/�����p�����Q��et�@
�6:x�g����O������_p�����L/5x�jhd���p�����"��Wo�GeT'%���;����K�B�t��Q�}nn����cg�c���QhzWcc��Ɍ
=W
L7��d����O�A��
M��SJx�)���I@'\�ͣ����-C��^��1��=?�W�qB.�k�h�uY�&c��m�KC{'=]Ȗ��?|�~���
#6u ����y"�8���k	��خ���w�ܺ�ZA��W�a��;�i.ʴ2�c]�nʰ��PX^���e�*y�a�c��Ef4#���lK.�Y(�6\�0"�HOL ���Wh�FA�l`�/���+��'�v�ٺ�;1Y\8��|��� _bط�I��av�`h��ή&@[	9u8퐚� :'��C{)4E�a�X��fEi,�1f�X��p�6/��`�XOl�)ff�V���[�h6L���D6i���:�����9�th���	Ba��̼�N"��`j��R���E�_nz���B�{6�a�I��ݢ�c�φ�M�I_Rv�X���t��W"E������/�Wn����!�}9&!��Z^6M�q�|�����$>f�O���M�#�60]L�\je�U>�~�|3�"���I��-�2ER�xW��E��u�Q&]�G�anW�.?w%�V��v�m����fYs~�����w�2��ѩ�J��[���+_�����M<�,y�=���;�@.�C���>�<���r��^�≛N�E/z|�q��2K�Ed֐`�����{<./VV���O�>��O�&Ҝ_�wr{n��&���wߗ��J��T&�r�$ �݆���=��뤓���G/^	��o<���O������'O��gP(��v�p������]�+;��<~�7~'�zZO�=S�Ӹ�λ����'���O��M˳�u��߈���wP*�Q������ğ�ɇ��\* �L�o������\��|d|�|9UJ)���dP*�D�=��J
��ݍ��ر����$j�<�15��/��g�'gY�_�{�^�M�@
��"]T@lt�*(�`�,X��?ԣ"��p�����!!�'�{���3߹��y�yw2�������μ���u_�ˍN8	��G乓�}��=���w6�c���8�����#c��091.	^X�\H��#��+��	'�,�_�����_��GyN�s::��}/��=򈐺��ax|j^�럝�ׇs?x�}�Shhh���#����X*�ˏ\��+���X
/l�,�2.x��"˙%�$(�?�dEؑ�9�*��ڿ�@T�`�(�$C��U1����h����g�Qe4�2��M��i�I)�E�� ��#$�6���!��_���fS�x��k�_�Cvv3~���:a}�x>�ڭ���ɍ���eX�tMte��J�ʳ�ӣ6�ٗ	���37Tʭd�H#MI@+9l�@�f%��ph�i&�cJ��?�ȭ��]�a��̬��Y�9�N��;�&��$�FV��C� �	�C�U:�C�p�"a������V��84�?�������Ȅ܊xK�y�m�HS��EIK��*oR�+�y"�d�Ӓ�R$%�:U�EJG�ς�0��<�k˧19҇#t ����лk;"�uh��CS]����N*�0�'�sHO��Ne�t���C��@�!����8�إ�;���M ��$�~gI���W#�ފ4yF�!�s�v� S�i�r��'���5���esy�O384���sڍ����ً��Aa�$�s�o ��^L&P_Ǉ.9�-H��G�G&؀��i<��aMyk�(��(��!4��̭T���p"�'�� 3�o~����S�`Qk ��,B�~"3
���6�U�٠ر��ذ�Tȟ}w����ρ����9�k�����N����G�A��zH@7���
�HKP����\���Nbx��=x��ǉڀMQ?>~ѹ����!����i&QI���|�2��qW�H�Z��7��x_��QrG�X����Ȼ"������������	����3'���]
.j*7ʾkb=�)��"�.'(�
	�c�s/c��$ƥ��o"���Fa������ R�}�pE#�56 ����E&��r���C�l�=5s_�s[:z�.�=Ν����������gt����)Ɍ�5H�Pf�Ԍ��9SNGCc�4��:����|�Yh����P�
Zi�����	�� 9���3���ֳ����i9�6I���5��)ɲ���־�Zo6��c�Kɕgk=��YJ���x��k��kzy�Z�D� V�A�h�b�e��YI�Wu4�L�!?��_M*D9'kmZL�Υ!%
,�!���Ղʄ�X_Y�Ӷ��w~[�KS���{ѥZ8'0(S�����f6T	��/I%J�
�����3 #�
Fd�$�2�evQ|�y�@��R��j2��G1�D(��?��J�T�%8�3D���p��?49ʘ<K������I�~�{J�09>.����pƙgJ"����ĸ�!9�n�� �صkq�i�IW��^G�n�vO>�d��	L�Rx�����#�!9�D����[q�Yga���x���
#*;����ʟמx�t��Ѹh�mذ�����R�	쩧���s����v�.E1O��*�b�ܹX�z�\]��ىT����|�8�w�O�݇7^�H�cC�5��y2K}�eˎDOO���D"%�8��PB������ �n݊����ڊ��n��#��o!�p���`����>c�chln�)��"���6���}�=سg�tuy]�ρPT����xԑbG�������U�Va���N�D������$��C~f��V��iV�CV̮A�Ι�uW]-�3���� v�z��]���|����t����|P��6�/��/"�kO<ͳ�c_g�z{/��������g�4l3��1�|�,s�$�+��40��"�)L�nAv�lH��2�2{ۼ�J�M�~f����O�?Wf�٣9w�]_�t�F���[`l�q��V��>�o���$�*ƱR�;����W=�տ7'`{>��j�q��V�Fu����#$��y+&��_��,iM�b���%a�*h��16�G�濕Gs9|�c]&�)�4*�7�����Dw�X��{T�þ�*��ϔli$
y�J�Kn������uhjk���^�������H��6��}�2!5,x��ƀ
�˙_!���@����W��Jin%�Fd��*ޣ4��3�C,p�)��0�CXs�,_؁�7=�w��,��u�i�bptHf�yʹ�<���Ҟ1�t9	�0���8��"j�n4�<�9��b����1Ľ%��ۣ�;��$r9x8�^,
������%�W�ly�ȦsH������K������%Ǻbu���34	t�:���k��)��6���"�1$\Q��M�rp�m��(jd�0U�#S���&a��3��L���]�
�Q��938�#p򪹈{�98IV��蕜Ȑ���P�&�L���'3xu���=���a,<v-�r����05�z�BA*pyqf����)�U��1���/el#�e���G&�T���lnÃ]Hv��|��@[}1_	�=�x\����F�$Z���=j���4�`�~��1^�{F��{��;~�k8}1��]���E�:���pz�9�Y�%;LQ��g�ഒ<%Y���Y"�2�����6��`|��C�s��i&��0�s#�(����[S�X�,�7������v��sb��"����2DVF�)�-����n��9N��+6�ZK���ʋ��z�,7�z'��*H[ـW' QI!�hg�;t�*a��,�VU�K%/���e�*�v���K`O5����l�n*�Vae����T�-v�jES��g��3�R�u@J@��Րl<2ɬ����v�rX���1�S{�[[�Ȩ`��gvU�S�Z��\;za����\����w�9�sc[�3�������!��W9 �:skul��Z���qɗU�֯��rֿ�}�0�?w� ���v
44���}=��g�(��9vE�(:>1!τ��#&���?���X�:�I��qѼ#��$gQ�"|-����!!$.����G:Ok֬��O=-�rd�ܷo�T{%Hv���1:: �>/	L��(�z$8�ѫ��$f�;;�l�tuu��7)y��Ab�
�s����@L�YLN$P�܂�N:~�_`��fuHp�q����(5��RTI���R�p,.���;��l��꘍���&,��ó��vmC0D����!�B>����G��>o ���^�}�Ad�vک���'���;��e�*��?L��]cW�I��ؘ�Zƚ����N.gF�}�Yؾ};6n؈�!�� ����UrɔHX���Ec��:���2��Dks�v�z����I:=	�/��؊�!d3�7�#�	�w����]���^$4�xs+����T�I��eΪ;���H�tFXT�������%q��7�8����D���D���5��@dʶ�3Ԣ6��6�I"Mw��6��*�R�#��b�B��2$UL)ub����͠^�c�4�!��$h�@Df�l�~u�sɠÛW�a�[�K̯�St��8ʠqt�m�Y�������#P@�N�m;<l�X=կ��y��2��ӑg��bW5�C5�$ٓS;�o����y�~}�r�X���c0�3i���@����b��v����&{a\�"�Q�)�Y p���d�TH��e��k���4+6Ǘ����%�\[$E(�{5[�z��Grl���&�Z���Y�,:�*�����ڵ*��$�L�H,��k[�Fp�i�GQj�eu=�pR�r֑͓Id�e|l��98鸕p���C6��#[�`� �GF��׋d:)��,ұH��R	)��@��ֆE��>^#�b&��P'��ax��;'ȏ!��!�B����G��.�$��p��֑m]xG��G����c���lYj�&�ʤ$aN	���-���Qt;��ri��-��R "aͤ;�l�	�p+6����=H�0�!��n:�ݘ�0���� w��]Y��*�y�����Z��r!�w4�!�V� lP��B��%̐�b&���R>*���[��7�=�7�D��#�oF�x
�Ps��!�i95���
�q�rp�p���7J���������u��N����+�11և�p���0��T����ymu�̺K1��Q(���q)�1�S�I��d$�.��#�����q���.<��z����i��hcrNf���(�ceBWCT_��	��1сX�0!�xY��T5OSO��ہ��w)����� 1<��d��x-j���>w2�$Ɔ�1�ۅ���������Y�)���-gc���[���ړ��M�pJ_����a�
�'?��-��U�=����'S(Z����i��d�։����O�~Ϧx5{2h�@Rn��w����gS�*�����~M�9PC�`N:�	fk�AIX�*�	�!�P�:S^[9/���+��\� ��Е��-���Uv�̚1�@�FK�5�!�x=쯥.�C�)�����"=��5kǼ���L���h�y��}#۱	Mpi����� ��yt�<j����p� �\�Ό��|��fL5�5t)��`�E,AK��p晧���}��[�wu"��Pb�~�S)�2�"t�D�IbR��(]A&T=�=8������cbd�p�_.��|�HD�ı�	� �\$	��={�`�b�]{"6m܄��w(B :0G�l�T.��(a�E!:�������124��x��Ѕ��<�G�(���N%%0����(s��eE���s�oɤRx�X�b�$Y�����	���KF6�����g�3>2�h��I���"�ڂY���yp/��!�Y�398]�9���B�@�D�`P��Ę���X�m�;W�KgWRɤ��j�Sa�&M��'Ii���b�hD�Zi���qs�Z٬�F؍�f9�v�ʳ�q���,�6�Q$G� ��Ȉ����l�����7��֩ۍH4*��T"���%!)�R�plbT���3�ϗyebד�um�8뜳q�����-���o݆Y��� <� 2�\~��B��A�Į���&��+���T�DǍ�J� �A�$P!Ru��b�.��d��$q܄�>�%�4���<��s��/$�q1���R�E(�{d:ؕ�oJZf%r朕SnC]�9��]�X���lҖ.�h�WuLŲ�fLC��2і�L˚��S��A~>������A^�B�ͭ�&{R�ݖ��YO݂1�{iӡ��sEf�)�gzxu�V�4�Yy�5��j��И;Zv2d�&���RH��im^�@�����iĈP�)�5�r9����1�ۋ��0R#Ø��Y�1�� �؊�ˏ	J�8T7�X�(�gΟ�x-
^HX�0o����S���Y%��[H��MR9����	I(+�5֠.i�������)��uV�*.{$� �����1�%?����6.K��,��Q��H�ΟGԙF���:�a�K�X�xc���z��L���l 9�n��n���Ã��^���5�R����YL�?x}^��֡��	s�΃;A���pH��8CH�_��rN/�� J5��
�⹷z���^�|M�tős��.h�lr�}LNW�g��E��(5���|��D����8bN">�&�ma��0�ό_�<z�y�x��x���Q?k>�-�xɍ�|	�p��p��J3Ȳ�L�(��G�|��o-��������!���BΑEbb��n�4'�&����$좟��C���3�q��n'�jb[g�)�d2@�D��� R�<y|�{�ϰ�{�6�g�mD�B�93Kٙ*>�âE5yfgs��O�Q��2Wƥ�.g�6�f��;�7�|����@B��S����P��*Lt�&m�x_?��dӔ�"z[�kdbв�8<�e��� � -=�����K\�����)qi�~����V;>W5��
̩2?�yXU�X܂�����[�_KaX�G��_�_T�q�DԤ�V5A_������OIv��H�����JH�� q�L���8,* μ
�Z9?���Z�S�����ed�@X�}��%ڬ~���H�;������̪�ȢB�ߙ���RP�i�1�5h���(���PG S������Rq�	���w�
�5��Y����M�{���@[�R�T=2����BR���N�ɱa�8��M�����s�>���Wxi�Fd���i5���&���#��H$FG��l�st�T��D����d�d'���`I�n�b��H���0ჳ;:�� ,�N�j��    IDAT'bш��Q��t%`�d��s��$�0l�2`V{���#���-��M�&ߎ��LT`�d���Q�d$aa"C� �Ϗ9���c�I
;;�����SvI�o�uBF����C�PV��Ԅ��V	�6��.%;uLv�؇��zS�@9��L����q#Q�3&E{jɒ%X�d��+��*�6k���?��h�ؽ�>�ǃpXu`�Q��<w��±�ȤB�#�&�����ľ��D��I!��l8�$HL�)K�?���Y��NiK���c���AM$������N�q樀��Z�7�c��0�Ҝ]	�/g@��Ӌ=�HqҚ$C:��s��9�`����#W���Oł�s1����l}k;�f�G ���!��=2{X(�՞c�A���2WE�,+��܌>�42Ԩ��,Vi	��k�'��T�`f��w�bH�3�g&Ԅ1��M��������[�_p��T��t!ۦ�K㻍�Q�H{l���YT������Ԛ����:�MR�f��f��?KT�������!EZo��%&��\�6�,&y���p�9�	Z��mwArZ%�m���:�d�63Ư��C�y�?,�����V�����c�$��l�$R�8K�#�ݤi#c���ӓh�?�;�oD�E"ra0�d���I�8�`�1����3�Xqgk�9����RE��"�"��S�(e����ҭ#M�'9](�p����?�>�8�����R��!�-1>!������v����� $5��ag�~7�B�EXq�4�6�A�0Ffk�W�XS��Hy��/�� :�wblpT:��u'�r�L������A��jkk����I,;9
g)��!v<O��7�Z�
4�-����!��M/��A��G��2y��6��ُ��$�٤0��9,�ӂ#��F{}5 I@��1ɭ��
�<R�	�@� v�ލ�_܈�d�m�5��D���'W0�h�^�W�9��N';֥�+�ɗJYW �`-|�0�� �Y��s���!$����G4��P������uW����n�8]!#�aE�ό8Vs��z=�s����>��P���"�u�p��(8�(8}l�J���i��%�
~Yv&�N��U����\��	Ө;W@vbc���2��t{
�����Z�$���7_6тHiT�Z���Uq�RE��r��̚i�NLD���Է���NM,��	O�K*~��ѵUqfOW���}���+��NaN�vږ|Mɷ�J�馔�"ڽ��bXY��O�x|0k���9
$E���ʿ�V(��iP���hu��t+ܿ:~��,A�qUQx��SC��^+�]��,'B���R'���M�g�[5D��*N����Vf峯�j�|�m�F�d-!��e�!�Qm�i�*Ō�g2��b;L�C}��`�tT�x:��{zsT�^�n�e�۱�::Q}	&Ԟ6l�*1��b���΂���3�y K��՗_�L&�ͯm��-[�{���5��H�K���$d��ܲ��q��cP[W'��A�j��d29���fl߱]�j������i��������ғ�G���?m�-�Gsc��F���$��-[�o�~��,�H
ԔUI&�-�&PII~��$��/y�駱e�f�S�X�h�@0�Fǥ;Ʉ��	�h�~��8�c��ˉ�&2�����)�`oo:���fD�a�%&�I�I��0Ijlj�)��"	4a�|�r�o�w��sdt##c�����>�c��YhkoE<Ac}��<&�Ԑp&����nL$H����� �G���H@Dqw�/���#u�q���#9�@<>�\&���>�!�����a�˘3{$]hko��3p��#�7��r�@���z��>�N�g��l��w�UK��9��v	"9/�/9�����Td�팍��-�E/q���x}�B�@Xg[�:;EW��V��&�@:�@Wo?J7��0r��2I���H'[���]hG<TOe���q��/�vc� U�U����tv�s��s�J�k{���hw���'礫�&�P8�
���� u"#E�þ*�ؖp�.GtJꐖ���8ꠖ�=,���x��RmNU�]�5=S�z�����_9�֝8�>�����Y3���@�ۈ�9����]����i��M)�� �-�;�>+�g����|�f�5�˔��>�t���3�c�L��Y�h�~
a�����;J���b���93+��D�Xt�
�kk����ʓ���>�^esi��1���h���Yƍ��b�����v%v�@!�<�S)?���	d&��L����0:�B(��dr\�>/g�I,�8D����-�I�%9�����E�B��DW��y<�A{s�#���Ւ|�s�L�o)_>��X-��:8�n���dZ����bs:5����kHJ��SBkk����Q���	�D^P����' G��P#Ɗa�s���K!l�X΋�+�?��D�֨�*��q�Y�) �; -L�$��h0�Ƙ�[k��0�H��ў�{q�\%�I8=>c�pȵBY>?��Z�cB<D�"C�x�"���������	��\�,��4��
��"�+�a/����	dǇ1�{.GMuԆ=�&�� ��l|�C�#��E���\�jgK3��b���d]Kg��c��/��ۍpm�M��5�� GNO�H'1�1���یE9 5fw&�1eԦ;j	EW%wy&�%�$�zz168 mf2$j��֊��:Y�%⺑�ə����*i��dD��S%6LB3�؛n���0d�,��˘ _�WӋ�O?��6@�FL�%˂��s.��Nq�悄������畽����J�1���W$-7�ڵTO�*��-y�|r]��v��[5�~q�K�ɰj�*e.Q�-�k�ĎM�ݼA��Ó:�-�q��K�]�-qJ��O�o��<��R.�ƪ��ʨNQ^ۤ%��ٟ���L]�@��r�_KbLy�z�Ha@����M��Z����թI �O%�Ê';;Vy��*%0#�lk�y#;!� !S�
"2L	O)��~R�X8o.Z$�������Q�G�;��Q_BO�~�z �dSs�$	�
�g�إ���K�w�^�(q��L��Xv�*Ѷ{{�n���IB@�x<&��A��ɤ@{8Kx��C�c`ǍIJ�@�8A����؄����EI�8��d�t�d�d�|�2
ٴh�uq��!���m�%)e2ƙ�T*#��`0$.����DbQ�!^S#����q��	%�C__���0ybW�<b�N�U�ϕ�adtL���?���.d&�T�d�?�K������T]; 9��8���U�XyL��477!�ˢ�P'�51q�C�C������f૩'����e�R�f�$V�_
9Lvx���ƥ�J����ظ|�z\py����\/P�������"tU׍���]"*O���C1��R�to8"�L�9�*:��#M$�����d�lw^Jj����*3��@E�Qt&�9EU�*�,��������įr��b�tQLa�&Ғ���|� [T�f�lSf+���:�~f�UC5+s�`M'��A���Z��;R�]@C�b
xҙ3�5$�Q,c�W��c	Hg�"��������5`	]Dֳ=���;�e�DuO==�gŹU��|��ڊ�VB����0��J+�9������դо˪Zg����(�T&�1U�-��'�^#u���%�I:���rzP�C:�R�)3ϱ�:�77���EAŝNdX��b.]q�Ί3C����6���ev=oSdQL�jDE�}�_)x��+�R��x����)t�FOw�S�qx��	ߧ8 D��HB�� c���8G��چ��!a����#Br��2��t��	IIhI�,R�	����8�'�&�u#T,bvs���}<�ĳ��jpĲ��(g1>6��n���R
=�1�����;��݅R)����	�ׅ��g0�I�1�q�՝}84VD�W��;��ӏT�$u۵�I��4'���������	D��"A�h��JR7�Q����\	Ɍ�m"�A��	�pL���l�qf�/�!�����p#��%�}�4�B�f��!x]!���P���p���D.5�HЍhЉ�X�=�q�G.����ֺ�d����������5�g�^zm~�����/��E0ڄh}|�d��tq��!5�@��M���g[7�|�5�m9,����{�r
ƹ�."�M�S(!��"�p 5:&�	a1OR���5l){��ąm{b}��u��3_�ubl������u�Fh�r~v�tmI�� �����D�>g��0�8��˖�S�B3�a�K�P�����6Pn�\��޾��_���oj�D\��*h�wa%5�o�)��P�z��.�,E{�4]<�K���{e2q���������<+c�	R�r���


��)��<��J?�g��|����B�*��]Z*�"P�,U�7,��b�T��+D'�Tħa-�N�Ru��LH��/����y6yRGU���� ��zS=�`P���V�tA�Y1�=�J���\m6p]e��]B]�,��Yd���=p���L!��䤆�3'#����&����H%����A9��b��L")�a�hL'c2�F'�Y8&��X-��mK$e��	� \s�l%����ʃ��$!I�0EHa;#s�tF|#��1�b��D*�L	S�4���c�Χ�8�(�$01:*�PX:V�#��!�}�?��&�i9��dIW��h=.��)�(�!�w���z�IJ=P���V�_����r��E!��x022���ۄq���u���ȅd:2���$\:%�\*VV�/v4�]�l	`�8}�����f���4|5�ʿ?��N`8���W�LL C!�XD��F�!L�GF����rB��Og��N�e؅9��Nr" �/�p$$�w�s�$�`Gi�lI6BM�B^���j2f7��\^FE ��Yr�4Q�.�Ɍ���z��Xѱ���U��	i�Qe,M+Qu����L�9-Y�UB�]�7�ٻW����b�-�*C���FkVa�?Ӱp�ܵ�=�3���ǆ@�6.!�fU����~�*��{l�Z)J
+���٬�YuN��U��T:/�ӫϕcZ6����l]���Q1Ȕ�C��E�$A��
ʕ:lf��4�\z�Vd`է�-2�@%�םA����S�i6i�S�9&v�\R`eǒ�� -~I:���g֢����:ŨAFNQ��v����kn��*�l�r�b��d��F�	�z��ﺻEɷb~W	f5cŲ��Gv2��x��ž��D �t�LZd�<.��D����	s:栳�[�xS��O8�����׷`���X�d��;�.j�@<Dj|�#ܨ��a�$,����s�'E�:��<�^?N<�d��6`��MX�`	����H<Ƣ������`6n|��u��N�Ho?vn߆X̏��ZD�~�''����p���ȸ#+z�9V�h�5H����S����R�T21�?�7\�S,��!��#��od�L_�g$���+P����r��D(Z�`0"��>��$�` C�^��t�8�p�p�\wk�{$�pM+J� |�ff�q`�[!�L`l�_�d\Ƞ���l#ݨ��3O�Y�����!�uJU;�����n���x
/m~���3x~�f��k���h��02!��޺<[�n�<��MY{\-z�9+/vm�g2�ӛA�+3&I&��`<֜���� �#ȥ'�y�NW�9'aʚ��mp����A]��l[�#fh��}�� j�6ؠu�X�3a%S~�*�� U�Kc꧊zWT�4L��͛�YV���d���I&�!W�I��2���c���(�ɛ��P��&Y4�t�k���I�Y{� �?��.5�izgi����>%�ٖ��TH5��<7�U�gfm����k����)}L]�����Ճ0���w����W�Y�i�z�����ʊ���fft������9��lk�ٺǪ`*�2sV������V�/�6�W��9 GQꬢ#E ��?D.��$�3FR.��-$o�T�bf��WI�$�O�e���qI��x&�G�`�ѩ�-؅�1(����H�%���"2{�LM
�@0�GFHH��v���&^###�� ��rх��.�d}drC��)���0�NHb��r� ��pnϫ:T��t����?�OV�3�|a�t��䘄��I`�O|��*�,��qn��aO/J^����q���
�V�hΓ��n���tucttu���=ot�`,��$.��SOgH��6�I�0!�g�zH �N%����!���={�$|�A���>�J���yqv�V��cQ���{�{�v��`ъ#0w�la���섇��������L��3|n'V�9+W������_���^:��%K1::���A�������۶m� ��\��qN(�x��R���d^0���"ͽ*�)#�?��6�§،���q��`��4J�d��Н��߮���dƼA��l��l�"f`�*����h)��8����#l���Sh��eA���_�w�u�]T��r2h�Z<b�m�U�L�J"�^O����4���M���
!���_�&CWWI�}Lb�Ȅ�b�M�p���������,4z)
�#����YK�����&w6�Y>{��*X��,3$d[�#
�/�Q!�Ѵ��{�#~�R��9��nDBaE�B�'�(r�PX@��o��7r���;Ħa�BCܣ�z�r�D����o���Y��h'���$�}�I����J��?���!]�a`���؞��:f�����Y����������/�c�<�p�Iعk76��2.\��ǭŖ-[�Ź��QB�6��م��.,Y��C��G�@�wub"�B�3y,f&p��⨕�x��װ|�24�����C��û�<a�jr����>�$�ښp�qk�����ۛ��5�Cݝ�s`?��-D��eJP
F�9Z��7:10Q�;T��$q���H�3�J�\'�\����懌��@�o�ȓ<rٌ�?y���Z�t{	���g1�%���B��d�G�K�2	�9�<@������V�qp��v�ӣ� ��A�H�'�m$'F�I�!�F<�E]�/�,L��VuN?�]X�`�83�ӺEL�&��ӏ׶��'�~[�ډd�	��H���$��&g���<qg^0�U�k���aSPJ�YUk�$W�J���� ����4��n���s�E]����Nd&'P�P�4��PG+�+ș����My�=��r�
[����ϊ�m��tml�B{��7��W���.����}�S����x��*���2Ϊ�#�����%��L��0	@e����rj-3D#����7� S����~i�g���+�&I,/2K��,+,�l���,ز��� �r{f5��h�t�O�=5�����$Q�7^	���u�
՞���yS%�]���S�:Ȭ�OI�*e`�mo[�Um.f�"�'�N
�\s�����}&ϟ���^�����k���)�����9䲊���q
#g$���K�O���'�~�z�Y2+��C#1�TL�<�l�h�X��Z��Ϛ���~�����y�p��!	a��xk�[��_I�	����̦�&�q�2#H8�K/��-[� ��c�e8��K���&�"!�@�H@V��Ԏ_��V��q������K Ey��.��$Q?��]8p�$#I�p�Y���3 �{�kjp�ǡ����[�r�G�+������ރ=���}��p$,!QMCC-�{�YX��H��uK�j2��ʫ8����g�E���/��~���H�c�k!�$%<J�KJ�K��ŋq�9����t����1�\�a	���_�w�>�Bg���8�����K���SN�?��������{ ���^�I:����{1LT�%I�X��$I���8�=��?x>|�'������N�wv���\���n��w����E6�]���h�c(�"q��tV%2����^V��q5�b��EsV~�N�Rd��t3���`    IDAT��Y��:�i6I��ӏ6�w���4�4�bfհ�%��<	��4���FfL�/Y�G}�܏��4s�\��}}<K�Bw�T�Έ�k
(=�_6���P��+�4��6�R��%+���yo���L��-�>̐�0B�����*{���j܄��5(I�)V�L�II�b�d���FfY�bE�Wbq,H\��5"D�T��
&�	��MR�d�R�����^�� 1PȲ���+�0*�Sn)��lm���[d��@lj S�@#[uaUp���dP"p��|���I|R���:���N<f�p����t�5��6���aI�6b�=�+�F��ΝB���T/v���s;�����غm�0x�Ysv�كW7������GwW7�ZI��?(�e2����QG!3�C#�H���m,��d��VlЏc�#Dg���
̟�Ɔz��i�4;N>�D���"ʸ��=�y�����'�A�=g	�d�_{&R�`BXq��>ԋ-;���E�[�Α���#��8��A�0�+��Bt�E?X!�h/�$�5j��qm�K(B&�z���	��S�N�"��I~�tfL�B���E��D�Y@}Ѓ�X�|�'�W�@�~6�N��y¤�f�*�q�Y�+����M&ٚ�Y�hЍ��:x�%S�/�FM,��mm�;g���C6�;��aǮ��>_��p-\�U�P$�21�fh����,8˹�i�A�1��Ѝ�1��L��@�T[�s=ܐiu{i`8|:6&�`:1!�D����rk��@���Y�_�2��
ԕ��ڨrn�N����P4��)S�o�l�#�4ݗ�����W�)�_e�Q��� �:\6�oL��G*�S�<�=���� B:�v����Vee���q�?̐nXiƴ��IvfJZ����Ϝi���4�|�*#c�~d 3�P���9S�W�ɳ��^L��{`1e�������L�o?�=Y�f�M��V~�w��<����VsYt���3��mR�){:tV6��9(4�z��ῤ�.!���_��X9^���z�B�(��(��S�Q�����\pƇ%�ػo������[;D[�ɽ��<��C/&F$��7N9�4a�|��g�������T`�����O�4v���@��g��^�w�����??�x}V�^�K8/����)�׊�2ހ@6s��Ѱt��9��d�^������C�xH4�n��Vd�)|�{����G:o�HL`���$J���s��	'���C]��\�x)^\����c����܍7"���W��-�"��,�LE�S�gb��)!!�9��cp�9�ƣ�>�����/��/č7~V��}۷��߅xS��122*3�ɱ1)t^z��him��~�SIXc��$��Z[g�ҫ����~��H%&��ÜY�P[S+	�T����l�R�~��hnj��;������}�1g�"|��J���� ����s:�"�
�����ġQW_'���1�}֙8�g��=�'�|Muu�z��H%'�_��+��x�_����K"��SO �N�s7~~��~�f�9�\z�ex����p����\�O�S�O~�Sؽg����8���p��$eH��ۻv�睏%˖�:�h/��ãIx��7)]��n�إ*��O���=o�DN32ڶ���3ݼ���0���~g�r��W��3u����VG��X�͈A�+��P�o�@�^�d�)vQ�iڊ���Oo�ٹP][S�~6vO��:���3�>*N�#Z*.P��&:%DP�E��F[���R^q���J9� ���O�͌�j�p*�p����z~�X �G�<U�ո+� ���d�rꙈ�<;|V2���?P���l�%i�(�7_�e����-8�8��*^��DM�J��ƀ^�[m�W�u����?�P�,�NJ6rh�㌓�`��ony˗,Dǜv8xH��{����c�e8���0:<�\.���A��555������7^I���6��D�`�[oan�l,]0_55uؿ?^xa=�^��0w^-^��^�;{v#��(yL�l�n�D���9KXs�!�z��M�;wb�0^|q=�jjpʻN�..�����FsSZZ1>2���z:x���GP,d��ڄY��p��k��W�ڛo���mF����w5�iMi "�d߱=L~��C%�h�]��g��"KO��r&\͆.Άk��Q'�)�D�vȧ��OO����8�w��������<��;
G��B	�@^2���B#���W6��,f�I�#�A65��ω�xX�d�0D,0!I�s�=����0&S���e� ���?q�>dܲ���uUǈ�*�ВЫ�L��vI�,�]U7F�2U�
W����e\���d��%�7X�n�e�@�z�Ol��	g�#F�9��H蔡�U�Wڔ��b�`=����Z$��H'��Rv��(��4Z:�h�퓪9I�\�;wUn���&�;O[����U�A�f�ic�$�V�"F�Vu�l����]�7e��w���W8+�1�}�d[�Щ��ٹ���<�25��d�e6���@�W�k榷��r��6,F�X=�Ҧ��;�2@*�+CF�R�v�;}�4R�9[�
��xS��b+Ag>��ؔ8��P�[g�_���V;��@�t�Q#��R��Z��jڒ@�9��=�{ef�}L��Ioۋ�=4�7��j��լ?!�a%��S�yR,Hg����`�׭�����+7߈�X+�;N�8kj��1o>����,�n�&ݷښ(N:�q��ڱ`�B<��3�뮻�d�R\z��t����hlj�G��K����Ef��o؀ǟ|
+V�µ��,�z�Y�����!
��眃�ٳp۷��R&�c��.�Z���������O>�/�6�"��a�+��x�"�����s��� ,��9��������y�������`w�va����裏���[��ҳ�`ɼ���7��͛7�{�AKs+���J!���O�"�SN9]t�t�8��ꫯ��G��я~g�}��Ǳi�F������lĕW])� ���w���.��g�%��p(��7o�ow/N:an��Rlx�m�h�zg'~���h]�a�m��~���Y8z�j��v-Z��P_��;v�?��	>>s�:,[܂���<� ��k�G�T���Ƿ�^��y�8gA�Yܾ�m��������H����3O�UW}/�����2+��܄��	�~�󟣩���^s�1(�hoiŮ�;����a�8�3���h�hǬ�Y���{��n|�;�	��W��5�����N�g7��
>���H�~��=8x�6m��#����D$$��S���3Ͻ�C���E����5!���	�y�3��U/ 7;b��f�=����)�U�PjjD��1*�U� c��J}n�b�:�:�M�XM�2Cg|�^�}�T�V�vw�&:*0�
�8���e�E�DCKU�Sұi����Zut5X��������]�Hy{\��0]�/O�
��1!�Jiלd�˫������r����?jB�jɠ��(���:h�d��AJ1p�7/Q�$��1�4�,E\�2@,��X�I��
P�J�U�8%��$'��s�u�m�̿fB�"���6�|8턣�u���S��v�Q�108���&��߉G��-^�מ �ռ�c�����6���㨣�`��ױ�w����b�j��� �y��{p��._~�����w
�65���kעop ��{Qr{1��``x�|��5X��uQB���N�x}V�<s��Ɓ�{Q����[^{S���=f��m��׷�F_� �=�DB�ٵ[�=�I�ve��UH��8�?��ۋ��}�i$sNdn8�~�Vʘ�^���XL�8�,�t㶂�����uכ�;��p����bQ�)�_2��."щ��qz���<܎�������`���3t��=�_�����O�	9
d:��@�"�q�G��'���� r�C�Id3	�)��u]a �N"��7)F/\n/ܜ������.□rb�	gP7J1ߨ*<o����&��z��� Θ}%�0�?�k�̛��zc���|��(���-)&R)q��o���Ð�K�M���y��Q���dk:�d�`&�YF�p��Ca�ul$��L
Ž�t���2�.��_]�F!K4+C�ojm�|�j�>��T2�9��`�Ӈ�2��O��mI���M����u�z�N���[\���L>i���i���FO���3S"�eȋ�_��aP��&�3��9u�S���\�I��&�fϩ�P�fed�Ք"�x�XZ�K����t敭�����H9q������G*��t_�*w9dQ�I�d�!ݶʈ��ʐۋ�`P��(aę�a�C�g2�'��iT���ƛ�Z���
�?�W]z1^{�9l~�E\��KD7�]����`��v����0w�B����w����~�Cر�-�Ι7�<��������#�~T���ӟ0o�\\{����`=��Z�q�?�x� �������#�I�B��?O�?���r�^�Q�q��x����2w~�~�	<�I�hV�|�c��ŋ����^�(�yW]u��F�v�w��؄+��JXD7lX/���V��?��O9�h(�3�:_|�$xw�}7�zk;��[p�y�	D�7��uuu����b�r�hRo劣d6e۶m���$tl|��?����sϢ���]v��(���	4����GC}~�ӟaɒ�������/`�����7����wv�|w��k47���W\)���}�6�#q\zť���os/�v����[��.>�K?�΃=�5]]��Z7o}�P]�!��;�555�첏�����v���q�%cbd߼�+8��cݺ�������N�PD�ʯ��
LN��G?�>��[�K/�8&�'p�O"D�_�I<��?q`�|��B�,~�ܞ"~t�]ػwn��d�y|����ȣV�k��E�db|�����{8YMo�������C�A��n_�X�� J��-�3�\(���LE�o�8ŷغz�$���k��"��)d���d��ܣB���SV��n8��Li ���5K�B���]`��+�b;��Yӿg!P�'�EX�ʖ�n�U<�FGP����1v�]�
�f���)w��jMVb�%�}2���2��I&M��.[��8DB�Yr��k����I�L�2�FQ#ŀ�d�@7utb�!�����DR���=�+j,�����Z���/U�O� �����$j\{�\�Q����q"2�29���tH��yl.1��-,����+0V���)��i�x/�Ii9��,��3T!�Ե_(�f�p)�^�&�]�P ��IL�6^�Ѐ��I<��&��f���5�f���_.����믿#��T6'EɅ�����6>��4@�>z-Y$6�3˛7����~�qhmo������8v�;�}���U_ñG-A[K��'���7��y˗-�QG-�D�Jcc�xc��Z�p>:f7����}���/^DM���}ݮatvDs[#�f5a�@>Sz���@"��� [�T������N����흉��>�V�&0zz��FA���Ap�0f��H��XXΉ�b��\@cȏ#g��Ȏ��Bpl�+=��&���g�	�m��<�u�Q�r�Q�J���LgIȫ��	 ulrٔ@D��p	fZX��(�NV;<B,���K�(9S�6��*� 醩��t�%�2fPh��T���'"C�Ӆ�z�I��2�ahR	����]�HOI��L����R�Z�.�`�i�f�y�C�T ����B�L_Z�*g������:M��rN��ơ��jo/�XeT���8{��|��)'���t3�S�?B�'%#��}��=�1��>@�����T02��D�{�I��m
4�$��&Y���r"g��*�&�#A���TN�m���r���`;�r�\%�b���Hb�܇�$�i�`B�]�vPy���S�-W������Nu�_��uW��:X:�����=���Li�u�l��i��#��2�����L��`�ߧt*h�\.�
j\��Y)��t�=7%B--���b��M tcݕ��m������>w��n���f����8~u�=8j�j\u�5�:ԅB.��d?�����ЄO~�K�H��靘3w>>u�����b�*\}��شa#~wϯ���p啗��ڦ�^�u��^ݼ��oҡ�3���磶&������]s�'���q�-�b�����/`||_��e|��u�P_� ݹ�_~Y�_83s�N��NI�>q�'��ݍ;�{f�����?-zg?��O�x��5?���'�����^^�k�H��|��ԧ�����/~�ڱ�3�8�ݿ��h	�����������JX�eW\!A�����_���}B��͟�t��7߄۷�7��.���Ĝ�V|�[�B6��O����\.���FB�����Y�p��7a|t��pf�kp�7
�<?w�����-�l���&��ً;ﺋ�8������xq�7���׏�?����z����'?#b���_���.��ݻ��?��L�x��Xjt}��+064��~�[X�ln��&����kkp�g>-���������b�ꕸ���ɧ��C?����8餓������q�k��c��W!����������76�5w���[��ۇ�W����E�4�Zκ*t���h(��"�J0[L��Y��
1b�r��g���F�\�k�p�>DDu�S����w;e,���Sɡ�*���~���"	�sg4�w�޵شUgA�I���?`��\��2�ב �:��+ff
�d��Mc!Y�f�[w�E[+��H���QmW��<���)��rdekeJI�7�#t^�dOX7-t�1�L�� ���)F�r iM?�
��H�ZRm���JS�4e��q���L���q�'h��Uc�|&�`���SI��xu�K�[�*�V�����8���=d�V���m�_9O��E?9=5�&I��d�dF�gD�a���4���d�ή���ꄗ��?��ƥ{K7O鉰ߋy��D� �'�EC�v���#�H1���
'/$�&l��F �,�������h�|CcK�d���Q�a�e2"D?L4��H\�]N����F��e���B��E��r/
�,��	�[�/"�	��J?����y��_�ZE|	��^}���I2��s�)'I �i�s&�����e�!
&�1B=Y7u*iNA�"'j�t4�aQ[�7Ԡ���1[�c4�/m�׋?=�߸)W�`��� B��PX'���V��H(hI	�r��b�nu!�Pd��V'�°���P�:i�y�m�w�Un�.Y���Om���6�1N��fpX�}2p�6��3}2h:UM��S�Q)����h�0�~0ER����Ai:�������Ns�S�346,�Y��O���9*W(MUO��
����{oL��M��M:ZhO��s��\��,�S5�'�
��^��]ӥ�㥍����j(�=��h�j��_��Z宛rbg����4�T�PS%���jZA#�3<檎��.5���0@���3uUR����8q2Pumʙ���6Z��\���4��|��#v��>W��JJ��W��2�<��n��i�s�dPh��W���O�U�b�u��y����U�i��2�6�+�0�gF�MB�����&��f�*���G{ę�g��9��Xf��"�,��\���"&���9���B�� �u������ҏ��m��עh���t�w��OV�$i������;�Dk]=.��Z�ݽ[�7�W�o�	^x����Xy�Z|��/b��q���N<���ux��Ǳ�՗�雾�m�����2�F��%_$]�_���+�������W���h>������~�/�P�6>�w<��'�$%
�&��+11��/�K476�֯|���׿���\�u����?�+W�ēO<-?�[�o��������1_����'��/�&�~�������[����  
#IDAT��gn��� ~x�����DSm-���&�I~�k_Gms��i?u�:8�Y|����EI���~盷�.����"���y��^�{��B,�{�y6��:��_�
�:���߀dv���q�������~�X(�k�Y'�{�|�{߃�׋���g���w�s/��\�k�[�7�����F(�O��N�}~\xх�����H�@�n��W���Gck;YU��ގ뮹��C��[?�/������ϥ�}��W���#����{��;mooğ���׿d�����֮A67����	l�_B��>p.��ltv�J �gw7֯G�������xO>�*��G��G��Uɠ�^і�q�g��Q�¶��ݧ\{7H�,"�,����qt'F�W�u�4���-��XU:�*�Tǟ��g�Ea��>��J�E�`��M`��y��儙��k���*��i�m˾� 2�D1"2��c"Y$b��c$�1�_@HЄDA`Y��l?���QH�D��2�ց�k����<�s�mD2�h{{?��9�9�9nj́<�2e�!�g�~�@!k�\>+M|]�C�Nk1�6�D�F�
L�8���f�5��C��(kY	�*�I��[!c��5ǎ V�W4ǘ�A����g s$a�x0++��Q�Mt�0�����Q��;�WJ�
C�`a���(̂���(JH�{����"G>�#��#�^�Z�զ$*̀$_P0h5B��� U�M��q���K�7ŊyrcB�h9��u��;"�X<�����Z0�P�T53R5�LVFϕT�*#[4@KH�/�3r!�l&#�b�.~*�䔤����ޮ"D=I����H~|Iaf�6aN*\�:��ҍYI=�d�T~���D�׉�'�KI��)#[���d�y�)��*�=%���xc{X����ME�o"�u�������� ޔ��&���Z��**��1>�|_��~\Ι�k�H&|�T�0}ZfLW���Ō�*LK���Iq+"�+��pn��D�/��z%T�$j�鋣@v���찑����1�NQ��s���@/�3V�	�T���}:}.C�4py��].�(��ߕ�d£Fn�U?�-��hf���?�Q���Qs�)�5���h_�~�RL4���Z9&y/�x/&�/(}H+֠����0_���Y�Lb�Q�z��I0"H��낥�ߕ�rC�Yq�Tj�n��U2�%���:��C��\��+�3��>$6��0�m�ˇ(`�&9��|N��J�"1���u�1@պ���\�Ծ����,���aX��@C��1W�"V1�h�%Ra�# �d	�wuhW�1�����X��mt*���e3&���m擅/g����;���*�����E�kpGD��J&��9wEQ���O��l�܆=#!��Y�Cq�nͲ���9!�l���������T�i��%8$K��{���� ͪ�bc�a��ƶ��hm^�n���(��ɓX�v-n�����_�̆f/�y�{�bg{;&�91`)'p��7"m~�	��}gz/a߾��a���3�;;e�eK3��a����];q�� �~�_���^\�?؍Tr�~rW�^�ٺ����w� r�65m��g�1��y5S&��kZ�y�߾�Ml۶7o���C2���*&Ý��%$���#�4.]��={>B]]5�ߟ����c�Y���6d��ػ�(ңi�n�*��G�����(�]]]���䬙X�~���)���a���hnnF6��ׇ�"}{+W�B2Aӛ���]�Fr�~�9�[�`�l$���]�W_� ��7��18t��Iㅅ%T���?	�[�Ѐ��~��;�ځu��A���ٳ�ŕt,�Gò�hi�"�;�=��/cɒ���;�'�mJH�I���d�u}zN=�T�">��y
-��@o͎��e=��sȗ���#�͟��,��W����?�ޮ�X�rn�}�{zp�L��F$S,v<4�Z)��w�v�L"�ʗ/��+�x������!l�Ԅ���0}�,��ˠ�t/���EU�T�"�֖	k�OL��y�tW���-4�g�[�C9"��� ����n�^<�����g�EcE������\�@m��T��%ᡥNֈ�A'A Ǘ|9�;�(;*u�[�&kl�� T�X����'aC�A���g��8g2g}>�*ܣLv�f���C\L@"�-����3p�^����5�#8�Ջ�uRf����� V?W��p>���0�ŉ �# ��iv��y��QL�	M&�Rd�f�k�:7Ѱ��5g�Y�9`hc5:s�UPIG7_�'��^<zJ0�S.�T��+T���J�%��Ղ�=�2hx�ՍUN�9�u���q�c,�Ԓ~ɔ/�#>�őJT�(���p�1��ʸQI�c'���ȋfV'=!��i#��C��|��q��Ӫ�<"�zJ^#�F;8�Ά��q5:���6_�7�	6���C������r��&�e.�O_Bt�y	Q������!1��k+��5ox�E���[�ʬ�Ӌ�&�QG��M��6/{�ޏٓF��YK8�	�d�	���ȳ� �����S��    IEND�B`�PK   �i;YM�f�  �  /   images/54318eec-5d24-4037-8f7a-d01382cfeac9.png�V�;ӏW�\?m˭޳I
#�{f�X[Y���r/�6J����7��P2���Y1B���܊>��>�����y�����y���9���� '��s�b�"�,QRB䛹6"��`Iabbj��bW��Q�@��{��k~�Q�B�bQQQzW���^�������[���$�:bl�Es��%=]Zt�B��6ɱ/�W����M�Aa�9�)N3|F2^;z�N2ɪ+߻n9*?c�������_���ᵦ����c�߹�ƅǖ
w��nN<��Ech~4�~YP �1�0ԀT�); G���d(��c�Gb.���g��z�1[|>���2G�-:�
���q[i��AW���HqV��<}�[n Y�"A�̉������pt����s޿ǓBBB�>}��K7����T�˗D"����5�ꠎ��s%���̱+���Z�5ŮՄ�lo�&F��xҰ�_��wZ���n[��ŕ��/588��)zL�v_�����v�j�<_�!�w���N�0o��L��TWa�CX��6Vœ<$����N��vW�Gx�ܧWQ]�(s/�T�A��׺�|8��Qd�����6� \��i=>�Aj~u6@�%XY��B�ßh�ɔ���%(�6�D���8M�Qwg��DJ6�О��}x�#S
n8	.�&`��>bޠ��*�Y�&�p��eк�ʝ_�=C�6�$��c� ��Um㕧�(X��P�.o�&Oēɏ�����xx6�A��Z�@O�_�*Y�� 9�*e1�iW)73q5K��O"@�0�%�k�����&{���Vz>�ھ�k%9��T)*�).�ҦY�_4�����^_�%-�G���{SSSc���d���V`%/[��@���ڭ��N}f^�^??|�Ҿ`ۢ�f�N�8�%!���{�;Mr���t��"����b� �]�f�X�ŷ��p���(�N�aN傛_4%>�qf���S_��S�-="
ԭ�����Q��������ez���`z�,Bx��dF�N*C��������Ȋ����%��ss䨅q�;������Ro%W0 Z�A5QS��ve�+����ؿi�Y��������}8	�/�>��4�C��m�φz-u/�=��9???^^^�^bw��� ���=� �"r�"�c��Q�{��,uA����9Ǳ�佖��y-��=�O� �����<�����qgɀ^�i�o���|K�F�O?�#��v��CIA,fq�[������IЌ���Ƭ�%�'28�&��tV����a���'�ß��U�O����ܞV��H�mn.9h�A--��C�b����,�����
vA�V8/ӌ��9���R��C�o�GrBhNd�*6B�����pn�Qq2�}��}ƃv���+q�w(�qׯ�Gm߸�p�(��`H$?��v����ɵjĢ��T���)��K���/0""Qp�~H�ֺ�GOl���A"s֠�	���ȕ��߂�?�}�$(�/�;KL[o͜�j�IhV��#�u� �"/]��f�=]x7֧)$N��T�ds�<�op�\��6��nÿ1�Z'���~=�H෸�.x��R��܌+%�"�YZ:c�Z�HLx�Q@�O(�Ä6��y4�,
���ҎiN��>�:�(s���%�}Db�t��o�96���_�Y��^:�.�"8s�885鋢�b�rDQN����-7䁫�����IfPK�!����#qu�Tm��Q�,u�4I$����W�嚀XE�E���ȲQ�-���?i������y^T�)����^���	�w�[S�����c���f+������Jد����R�_a��y��]N�8Jc~� 3m��p�wW�NO�ɫ/g�Os���%�yz�J����w��aK��}�;�{$N�C��W���4��N?���~j��	�o0�9#[�_��OP������a�Oh�Aȕ\f��\i�n�������Ⱥ����������J0*6+�������Y��\'=��C.E��**/��GT�2"��\X7.��V�
~�۪<_-���_�h4�6��[;'y��o�@$���P����\�ǥs�^rl�Ƅ�Ӹ��1�!`ȵ���!n��z��,���wwTL��Ve#1����b�h��7���=�Rrs�a0� �EH'���|F�{DX-���g2#Eg�,W���P��ukM�<v|v@ !���� ��|sO�{���rg��=s�s�T�/&�PK   �i;Y��N  +Q  /   images/55dfa5c9-aad1-4e65-bbd0-3dabf009b856.png�|eXm�.�FJB�[:����HwK��)����������n�l��;���%��f払���5�)+J�""�����H�������߈��O��f��uV��S>J| C##.����$��\Ӎ{}��<�����ߊ��5p�۩�|���P�^)7�)����_�����LcH�4���?k��"��W�r�<٦��[�!x���l��4]�r��y�C��$Y��,���y7�����KA��Ɔ��L�)p=��_�Q����z�������a����^C/��_A�� ��X�	���o�N	2X� ����9�a�XD�{�0��P�H��腈�0��0,\�1�&0B�eQ�t�bX`��^`�/��` b�"�����C/��s���.���x��>S�kֆ+�����Z�!G?1���3ϚjL%a	�<2Us�=�����5R&��t)atRB.�ya:~Q���/�F������Q��v0��weѳy84m��!��ܺ���;t �ڦ^�D�w4C��ǕyH���f��W�{���g�tŻ��5�^�W�#��TSap''&������}G��[�\]\�%u�j����%˩�'���jI��4���_3�/Q��,d��L�{���dz���}.G�.���Ԗ�B�H����1���$�����45y���S��,����2>�}}4/�����p��97o�P�+l�_��"wq��,�����w_��}��K2������	q��JE��5�-늶ke���:]q���2$���~�Uh��l��Q��ݏ��T-Y!xHHq|6Z���*�����E$� 4�F��paFV֗��lRRRS�£��5�')�6��������~��	�����/�2�N�4Lz#� ����Yݘ����ȿ�i3n�?K*~L��Ws���.:�ޣ�"
/OON�����p�՛~]���*Zc1l�֑�艟���}Oc~CϏ��GI�2������3���kӫu��iR{��󢖖��I�ҙ���Q���=�(«�Xa-JPCs�}tZZD��fɒ8£�g�y��i��;�N)�@��uFxa��5ao4IKim��@
�餮p�>���U���dJ��96/´}�����ӎב����ԡ+�--GY��U�^ž{�������6��EZ66�.�P�cx������ħBj���p��7��Z��T�s�U.�w���/�3B��>~QT�255e�ȱ�z�ED�y���S�T�u5���yK�T�Ik���
q���n`�5ե�C�DD�i���!��Dd[3ssRU|���]�`3:<<�ƽ�Ť,���� ���z��ȁg;�¡���}Ĭ�Gbb]sk� 7x���i�c�gNXXX6ޛ�L��?ߘ[c�{��Jɧ�Hn}�,�����j�^�~l���af��������#|>��� cL4�\�J�b��+���Y\^>��:?A��``f�Y1��IS,\��\�߷�Bb%�B�cN*|TȠ�QV�cad�a�1��]����!+'gȞ:bs-��Y5wMg2x���������Flӥ�pttd����"cRG}eA���F��abe�z�M���V>��izzZް���4��p7��b��v8��A[�N�k�FTpX]�Y��G�`T�������ق�C"�����έި����1�0�̤}�n\�;�\dE�Ř=�����A{����՝]�1L%�3��EOLV���F��g�ǧn Yߜ��u\����U�t�:���"7�,�AU�cxh�J����7ď���S�h�C|9�����RAA!@e�`��w= Asfz�)���g%�}x�7�UD-�o���t-�+/��b~z\�hA��-�$����F~|0AW�U��"IOf�d��H��M~~���5�G������}��cH���=(>!�����Q���$P�S�3OCK�)�ѧT�=�'=�>~�2|e��%	�+051QCSC�]&܉*�Q�����I&aފxi��k�?t6l�]_�j�c��ǝ�Yn�&|�͚��"����~}t�j}��)}}�jw�QX,3s�|����_����s��B��Vg%���#���Nέ�:�-��F���=k+��Czn����ӕ��j=��+��)��*�Cu�J���WjRy}��K
[�ml"�Qļ�������[���yS�J�!��M��8��]y���o,c�����®%�M+��gpY*�����g\�L.Ԙ+*�^���w�Z�%j��o��r�^0��&�G��#O&C�u�[n�W,�2�Ӆ�w^�!��b6���������PZ]{A+���@B��S�)l�6Y~�%+C8�č_9z�K�=����N�gz)\������Ǜ��S��V�l��fX�����9×�,��ڈv�v�`c?��~�ŮW����sH^.��Kj},P,ۂ�5��v�:]��cg��hNX��l��[��@K��]Vv��-=��Ii�i/��xg0���[��IuD%�Q�����X�Ӓ���J$���Ȗ�\���DF���������+�����R�V�;�n%,�ζ�Y�#4>��M��uy���f��\f���i�G?�+?$�p��R�O�Mң��xZ����+���\8,ZEos��ܿ��e�L�t��+�T�]qtx�1�g@�g��!�ֿ���(s��F��a7��SA�y�����!n 	������!5�a��͂;W��r��؏�[}d�(�>����<5�z�>\h"�-ǐ>Y�H�lp�������o��La��}>��S�����M�)��F/��?�@( ��1- @"D'܏�+!�ߺ>)Ƕ��Q�0�����H�y+���k�\�^��i���H/{_х~���қ8Dw��Ǵ�6)V����*��pΥ�l��P�"���N2�u}{y^��~��
��֗��ծ��kG�/iq�D�M�7�_�z#	.��lpT���L;�[�#{��+C�|o�:^�����DFF��vd�,~_�uL�8[[%|����ҟ�E_��ooo;誒wp? �$ewT��&�s���گ�.�v#�D�2��`	}���~W��3����%ڀ�S�lp�����vɭ��f�I�E�}kzf��wyy��P��r�#��[!���i��|�R��mANG9d�S9�;{��-���E��2���9�Jr#QqGs����D��
�t��	���lh�B�4XҀ�p��Q�H��������
P7�������>ٻ�R]������㙱&B D�5�վ::w&́C�~����h�Gֲj����H���
�ÄJ��O\��x������F�ĽT�y��#��&&[���?#�k���cl>�*���6`��I�O4�H��6��ZK�M �M16���jhj���ꛚ���!:�����K��Ͳ����nŇ�$��踕V[[����Mܗc PΤqggGx�h��f�˝��;�m�� ��P����g		��l� ���;�1�޵5;;;*���#w�!=���Yv�W��ᐚ�B��w�e�����D���%<�LD�@�����g0 w#F�8xH��!�������V'j�L����0�,�1�%���1���!�D��rvyY`a���{�E����ϟx����˦�y��:�JKSS����,j)٬U��RRR��XG�kj^rsr6�<�()�j��W�~N�3���g�`y�n��K��l]S��ܩ�*x��I
5E`�d�A)��v1�~Q���T1%�=���z�B&nn�888r��Z�����CCC�m[�y�D�vi�����5��H���R9E��lw�˱є̨gff^
��]F��54(�ED���p(E!�t*��?22�~�܂�V��\��f��\��q�@!uw,S�,��J��0���������+U3�ݱҒ��+Ñ�L������>����Ij�r4�gY��B��vH ��R �2*p\�qY�
�97]K.t�F��w��I�zc���ML���^�F t
WA㘋��胠gp y]]]g��u�t���X���V��p\��n[i
��!������qsS�h`�׵�p�լ����l��9�,��j��Uq���\ N*�/�!��O���@i��O��8ʝ�����,����~�:%��e%�<q{@c���+JII�K�u�=8$�EX��e%%q�)�Q�"�0mw��7���/���	Đ�\�T�,����@r��^5��"d�[�A�1&X�-�Zm:�{+UոlC��c
HkU�_ܖ�v�ғ.y��F݂���^@B:e��VNa��=*x�N��J9���(�ݏ/���yZ�⳿O�$IO��
�<�>���0�Z�ڶ�RPl��,KD�i���my�
9|�[\\LFcc�ڀwp����T��dt�g�*	�&<6�s===��}}gh��90ێ����ms�ʜL4A�r삁C1�[/&�&��\^U����\4��8ܚQ���dW
j�$�V���qHO�L������,`����C�D�4��#��y�4w'���͆+5!)��[C#1{/f���G_���4�Ŷ��j6ˍ��2I�����z7+�C�s�b�BW�_�^>�AE%%�삂�}��@�Z�o ���e�gt�45��B���@����� p�L��Ì��G�� �qV��V�k��+ �����I�B�ݭ�s�G�h�Qw�����k�b�X������Tg R���0�$�{/��B�%��������ZGAu��8	7������A�D)��Ǵ��B<����=���,-	�����8+�lȄ��[[���� ���'�C��${��p7i8�Q��B�8�n�*���~��mج ���fJ����[v��̑��@J�MkO^�^�Tn��+��r������S=J*�qW�NY�EV�8��%Q7�oZ@E�3�{����v~ciii
D+j)ѩS�qh���b�	X`ro���Gh��#z�����x�ⴕ�Sck��M����zF��y�-�4Hi}�#��_'����ݑ�;�^�'P|=�}�nT�fy��#S���vS��i\�x��L<M[����prO__�' ,���w(s� �>l�;<::b���c�n}V 85�����j����`�p��6��x��+��t� p���:q		�9}��6�gT��]�U555u��
|i!G��b0˨֞�ʯ~u���nH�봭�+�|�g��3���"j}�J���q�ȗ�+��'4T/y`��T���Jm9��vssu}blc���[�Z����,E,��2yw�WQ�`S/.�H�.ۑ�9�K[�bÕ��e�熓	�8�P����	 ��9_����0��HX�г�5$��Q^�٢?X�G,"�H�^&p�=�z���ݪ�8�Xq�k�+:���>NYYY��j���w*);≗�=a)��OE,x#�d�C.�B�$���5�����/�#�ywQ��p�R�t���I
{�hS^�2����yI�"
ZƅK*T���!3�ND�p�t�������w-��^�ݷ,�05�&���lT�YtY5K_��yxƝ�����1�qq��
�~�w9NuQ����5�T��Rca1�zG 9hR�G�];E��KD����}�w��\JIO��.�ݙ,��}�@���,I�pH]O�����k���KyIş���i�������&�����w���9��t֌W����`���S50Ķ�㐋�N1d�tH��g�ɿ�^��k;1���	evk�\�@"��g�v�F1�{#���hi����g$�f�aX��>�y2�����'O������`͕�A*��2xIHH�,�>�~����I��	-���u������Q�	�G�>b�q��eZw�^��h�G���>�,o��g�jWO{�W[�xlu!-�0�mOJ˼y3kX[6.C;����f�x����u�V��(W��
�W�X�/L�rs;�ո���]��_8�\��\>����m7::ZN�|� V������33=���#�c�,;,�����*�F���W��a=�~���ѕ��)3�������`#����6W�P�ܺ�7�g�$��'	���uȠ�{�zf<F��a��]L��g�'���=c;{{s` ���f�b-___W)	^M�𻟂������������*����|ݰ�54d�hۻ��2<�4���ܴ��U�;;���ust7��WԽ@r84Exh�-hG�[��(�M���21u��4���p�����j�$��
e�~ߚ�����/���>k �q%�sM���H�}s��9� =���B�v���V�S�kڲ�Ŋs����kd�v�H�j'_�SC�`gQhEb���UTDWUZZZ������Յ�>;D�)貯<d���t~w!#�=��qQ��⚚����u�wp�GҊ���cn}$��N��7P�������f�x�`��P��k�*K!-;|C��ތY�P�L��A�ZPH�R��_E�<,�s���MF0���U,A1���xk!�BJ����e-�%t"x���T{�.գ����u�s�V#�5�,��= �s�������c�$�;�ZPsssmR�˿ZI5h��f8���'���'˷��K~z���ڞ�2G�S7�q�d�
2MLL���l�D7-qG"�'Ψ�̓�T��~���D����BjuY��t���Yx�ޭ�i8� #�j���z56ZA�L�ZVi��J����1�����J}=X�����9�Ӳ�6d;_�g*�RuP��L���n
4��Z�:i��Y��i��&ͮ�6�/�M�{S�X;��p��o�umE.�PV�wT�o��6!�o	���i����jI��h�6��选��W���y���|�e3�pNަZ��~Q��T���ɸ'��L�jSCI�/]#���9?j�<���*?���w��(2��(U����W���S���p��~E��%A3B����(#�P�AG�(x6���)� ��tD�Z�p�Q�F;�f;te���R��a�}��u����F£�H�U%Nƣkg_�2�-/���{FA�'A�^�R�8j�( ��M�J��Q�^Yy_It��ˈz��,�ǒ����J�;�C�De �o�N����\N�׾���Č���&�[L�H�<�y�h�&�����L�s4�9߻7�a㨴'��0��EUn=�U���f��H�R���	x�:=&�%�	����E/�:�
k�ѥ<)��+~����<��y��&����\SHK4tb64X������S����R4fwx����{��~���i;?�C�@2���b�ȅ!���d��	�(u|�FǝˬJ*��`���nI�%޶��@.������.�H�=���#�#�oX�耗���-�&�!Kx�����S��2[���nf�H,xŽ��zI;�n7������J,l+zK��o���"����j����[N��nV��
���&(Ă+h�A�:瓸�f�JWZ� �9Wa(�<�!�L?M�V8����W�B�`��JG�x��N
 �� %u[T[��T��|ʠkkj9�_�Jbѿ7���/$'o�(�J���Q^@V�������$���RR��<��� 76w� |I�#�- np�*P�N�>�i�L�/��,���9�C!L�#�;�\[>88襦�F�@���Q_�ηz8O��^O����z���\MF�~��C8��A�#��mK�P�����������APJ^>rza�^1�-wF�������ߜ��d �a�7د���z�'
?(+N�S4F��^-���|������zs�x.��*�ReҧZ�ψ���}�������<H�#���AY���D Y� �����>˄k�|s2M���t�Qw�
/K��ȈON^޶!��}������"��c7�f7��|�/��пd@�.���p���D�+����ݶ�	¤���Y��~���{���g] �c�<f�����[�.��"��r2/���d����,���)���L�Rz��v��,0g�E�3IB������$��`��J\Wx�3�����_���93ߣ��=T$�n`L<�w.��Z��!I.�Uo��X���%��F��g�ע�K�e�F~j#`g''_u]���o�\P�C���`!#3�����l�.�	�}�VZ�� �\��:tڢ>+��x�W��8�^NH�A��;:����Q��Գ��ר��νe&%v��ſ<�ǳ;�&�yt|ɕ:Rn�%!�U״�G����d�B�y�J��ФCpd���(#�ݬ;ul��ր��Q~�B'ud�gII��v�q�<��7��*뺼���&�%�XZ�5�Ͷ�'O�8�k5�ư��"���(ư��+"�#��Ύ)b<���"�a���W'#yKK���_�ݗ���.��/
�@��u�!��b��٩�.I ʅ�q���2��P����&�R)��P��������������A7b �kI��TV@���7��݌舢��`V�����@�Q�&~�����6�@35ӆz�sr��g�R���B�F�ݘ�#W��(d��BFAy��L���G�<���S���DS��d������1�;*F�ϸ�� �I�Cs�>�D&B4�aj�.�M��Z4P��@���}�s��o�P�נ����i�P)��}⊂�+�� ^|ԽP>�a�_g�4寂`K����MV����c1����gG� I=蒳��w������u�7=M�m9��E���$=�*WRT\��Dm�3���`a9�"���N����O�͢o:%:^�b�J���ښlnm	��sqs+�����Q��N 㾕f6u16�D*�[��X����t�>)S톅��bY�Ŗ�NNN nc��`�@0 n�m���Z��[6,��&�qRSS�~�������Qf���-����~�X=C�v�n���<=�U���h|�b>P"'\TTT���Æ?�����/?9P�V��۽M��>�DBB�z����&'//�ߑ����}�  g���P7j��^���#v�DB��+@��dkƭ�	�M�3�+8��
N���-��X.,@�h �ƍO� )��������<���G�uh{�, �K� ۥz}N�Y���d��f�]|��9�k`SXp�*o��L'��_̀��)E.̇82eFX5�|���裿f���u�b!�������-� ����geg�G��^�+j���^QQZ�Vę�;��w����M�`g|p eq��DKd��ꏉ~C. ^�w����}���[�c�hw~�'��/����^�F��p �PGq�a+�~;�1|ݘ�n�����`�_KK��z%����=�m6�����
���L�}F
!ဂ�`�N������`G"g��}&���Z��̔��n�h�X~~Orl�=!,����6�M6.��^�<d�p3�?a����;��	���7B@ߐn�������^�u.LN���w�!d O� �t,���[գcBo b� ���䡪�:)e���¿6�
�6̹H���uON$L��0�"�5���Z�X���vXZZ:��xp�	�����17Ncӂ�bp%f�9)䀕V��@u�t�)�: ����8��"r�d��l "nt���MC�Y��������Fw��Y͂|zzz܈Y���d��X���{s��w��c9tȆ�w;�������������|W��$J�����EE6����s����=?"�}��4�(�&�� v�CE�d��B�!O�:�:�ock��'`�;)`@��Ȥ�LL.H�=�3�<�eo�s9�q���S����������1kW�o
���x�P�`-�Z���_?d�9�0@*�H�{{/yEE��x�y_A�c�p��9޲��	���1�88mٴ1�-��MԘ�䐐1yf��yf��g!��j��)
4��u�em�cf\R Fp|�$�f@B����=N��d�S}�x���Y��MRZ�8	��hϖ��ϻ��,#�GhVi������?����#��r�X�vo���.JFV�h}rr����&Jn:??���`΂�|��`l�\��f�Fi{��ݹ�� -�d}CC����<m��/pUY�-r�Cw�C�wraᗁ���̡S�WS�w�vr{U�#z(��ͅ|utt~#�M�e�}̸J{�&o�������@�X���tTU)Q�5�4�t8%䇇�D�Z������E�fa�3$/
���^w� _g\ul���~`�G㓹�6Η��D���$����� ��e�7��b����o�h�F@���h8.�=���T���qM��`$A��}���{1RQ�(5��3	�h�����#���B 7��'{Ef���~O��$��@O1o�...����/��F�yE�LY�qAp�P���0�Fd�W�7W����v��Pbb��/"�m8�����uN��͡.^\p[`ցR���)�^Nʱ���0���sX�B��4�-{5�'�j'm�M�Y��=x��!+\;P4vV����f"UR����rsO!���<���I�:H ����}K�{�qa"eYq�,_�B��s`�� ,����~U����A��|{v�D���ŰI�Vų~^�y #�����3�����u�ż�����\�fw��ɖf�:C7��B�#i1d`+n�z˿O�{�"ݲBZ��M���4FvXά�?<������Pv^U*%��IHH|/d|8�y1���u4i�����<�FAf�&忴J���e+j[��#O%��#	��.?s�4,�"�f�`N�¬FZ[�LHH(X�c�yWc;Y�Y:���pHx��8O#��+YL�����E�������b$�̜54�"L��������<`�FZ~�:)�F��UVV�#���m-s��6N��T $m==��P�phY��C�X^7/�E�xE�6 �'ĕ�5�;��UL0��F�5.]����\!.@t��^���T��ք�� �]�8��!dcA!D�����^]:�Vs����Ѕn?m�@}��aQ��]Nb퍦��C|�:Ȏ����G��j�^�������ZB{� �YA�����~���X�x�5�L�w�n��a���y�� �0���˃)-4�mF�R94be��AH�pZA�������I��ssM���@w{�~B44�����*�X;oðh��]g4���9Fn�n��\/�����x>܍2��t�� �&n���� E��)���j�ё���v%��2����|0�M{|�� �-��|d�B�|b����g��82�-&,�6��J���e��ݕ��K�T�PH�����"�-U���zCBn�+�pp)�Q�<=-���w�:x7�ڷ���uߟ�����t�P��x?]�u���p�c$K�k���t��ϳӵ��`�dOKk�nQ�}�--!�c������C���������bd��\��$u�4E=��I}QJ����HI�J%,KZZR�.�O<��l�i;��$w��=����/��s�-RGh��Z��b�f�*�0�_�Brrsw����'>%17,�\�Y��`�����:���9���7�V����6�6UU�/�pf�vTΜ�T�\�d#��)�tz��
r��������)eQ�c�*�9x��" �ǾfaT]C�'??��XT�R��
� @%!%��}��17Q���෡ԫ"�?E������7H4}�i��\?*���m�N�.��a��6Lol��rL[�>.[�]����<}W+T<Q����է�]�)Į�-Nd4٦>��G���x�1���v�6w������_��:��r*^�+�b3��KK嶏N��?ׄק}�l�fCo((�m���D���~ȋi�uj�k�75��W�_�&��Y12�'�P�'\�p~��wlaiI ��C:F�'Pܟf����x�J�j�]7��������K�D0��/��s��4A������tN�;` J:��D����<U�3(j
ulmO����ן���6zw�g�z�Z]�����g͟�)�$�E�~+Gsw[��RaP6KH]E�9��($�`�To���V��.OJ��蜩#N����Y�g��@��î����{�7��9���	����Js��G3:����K/>*Z��N�@��N|���}�a�0,Tzh�(�u'�|Ο"6xEł�[��W�_��Bk��z��&''���O�K�u,i��1�!�ظ,�[z$�����\�Ƽ-��n���;Y`��bĢ������z#	j�R���|�~VTd6��eK.�A�����k?�P���[���'4���N.��CZ(��'K�I�׮_��T�t�����c��[\�f���Jf�D�DK�A�m+-��e(����>U�� F����O�_v�c�`�h�5�^}��b��ChR\nr^Z߰�j�����Lǃ��7 1(n�@���+++�����)
��H$��x�O�C#αew���hրQO0�#�o���:���5b~Ko�6�cE�����]AQQ�R&.�Pb�v6x$�h����ڿ�aD��'$�t)�����`�/J7�Oށl���be��!� �-����"�e�+-����r����~&}�,����_K1����T��>�eu2bd7��E�)&����=�|݌�-�����$�`��v�T�HK�|�������K��b��u6p���>�WP�}�H�|Eĭ���d�Fbi�����#���.I��ܬ\v����TyJ��7&1{������k�#n�E���;���E������ ��B���i��su����8-E���?�;uh�_�jɹ�;@ޘmR�ؒ�z~2W�x�z�`,�+nȤ�;�V��7��5���zðw�K�8���ĺm�Ϻ8�ǰ$�Kc6e#�h-V�?u�$T������xfW��6�{�S��b~}��@.'	L	�EV��VR�#�=�k�쯟H?P l��|#�ptxH��Z�e�_��m�|������(�"H/.>��J�t�Z��2FJ�W�U���� 뇨�'ZGߔw��>&ն�_��V.��nU��-��qГ���p�Gcퟀ�p��(5����hʘ_�E�<k	��"(hЅ�@��ywx�l�G;T2�y�{`.��*��4�%�1��i�Yu |u��$}���~�c�VxR�/���}���|1��웵 a�Н��8/�v�e�M!4s�K7[��p��b��1c�ȡ;+�z� �~�$�=����|���o�0ؗ%��z�^�����Y�Ɨ��̽Nz\�8V�ϦN��Q=�yI���a�$c�J�QDJ$B�I��(>~����=`gg���ȧ�eb,?T-��w밴��J�0f��T63�����۸y���5��]��Ͱ~��q4t�9(�aZ�iWS�u�S'�H��M������F��U�p��dc�=��O;c8R.�6����Q+�Du�B�`���i��dh�@��GS��}<�Ct� �J����1�0}�D���A7ɿ�B+?�}�� ��'���jJ�����ɣ�CF06@��v�&%3���,m�&D�� �{�~�7��W4o��Z�I�qB@'��p��;@�%�sD^We
*��h������g%1�T���p�fpY]&�.�O���[Pc>&4������ǿ#&D�^:!	@6C�Nu��c:��Pv�@�x|||��ҁ�wcI��@m3bmM�lόZZc�F��k�:
��lf7��4�_.������ՙb<��%�R�lS���΅����Kx4�^������46�JDi �~�n�*T��� ^�k�dll<~�NĘCA�.www7$++�9! 0r5s��]�Cmѿ6I��➍����ޏ�"������U�}F�{���'q������TX*�q��� ��J(2I��EQr5��:@��+"G��/nm���Z� ��ƒ*��2����38w�C���RBQ>�a��F��"��iii~����y~#hZ�Q �JV.���	�@ǥ�o�z'*wD� ��H�� ���`�x0)�ֳ���EMǖ�v�ֲP���aeb
����Wlq�"�H ^~��
���YbN?^�Z"[�����	p�g٣��84R�Fm�X�ttt��@��X�����s]|/?�uxxhQ�#>�]�t��^�S)g!�	w[��v������^�� (�RB��f��Դ�����
D�x��S�4y�o����i��lq��rvz�uӚ4�1{���+��Q��o ��rx+G�]�5l�8�	eb沿p#�Ԫ�E�Z� ��|qt�k9۳���lp;��J����0��G�#����P	��$��5��;��ȼ9C�'�S�D���� ��#�\�����v4� Z������n�q���Ė
(HP�?���������}���d���MbDLX�e�������Fs)��򖖖��+(:�""�� �E��e!�F�k� d�m �{���E��m˨X������2���4���T�Q2#� 0��,,��˚�z�*�9C�	�I���gJ4�LXӑ�G�j�S7�dُ->`��A���af���b�<�[�!�,_w@=ҭ���^) 0�
��Y#�0¼�@y��F��	�ԥn$tt� d�6F�u��e�%Ň�(����S�Q�3'�,OP�������v��w��-�������&f�� �~��M�!7a�K|��w�j�	GeW�KS,T�[�YYY7{�V��,-N�|���5lJ���浀��('�Q}�㛠�}kR>�03	���
{m� F�.���^D�DM�Q�D�L10 E:�����5�¡_I�h����?X�� ���*6��?4�cu#��ZuH��\���0���/����;OJ8xxR`�3_-H�SHH=A)��t�����Z,���s[���Xꁟ�عM�V���~�[d����~˷|y~�z�,~R033��d4�|C���������Ɖ ��? D.% �z����2DI8Tm�ụ%�� �G�(s}��N���=|��5���{��V���29�Ǐ[��Z��-������ii��3z����𑑑�mR�|�+���H"Q6��$ �_� B"����k1�U��x�&[:��_o�Ʋ���EV"�q��^A�OB�ʠs�O��1������Z9r?,�t�����fE�A���AZ�f-(l n�fXB88r��*%i! �z�<�$T;�+$� 6�V���Aޙ�e�h��Ht�/��+�������Io�W�^�FD��N6h����,.�\y$e���5�Mꥈg�*��Ӎ�����!��
m\  l�B��ѷ�6�\+����b0��!�����kb�y�2�� �.�"nEh!����:�����L*H u���7Ŭ��`m�y���J$��6D��@����ʒ��]a���r�ׇE�E��5��HLu�UQ�H��Z.;v��G2
-����ϖ����L&΅������!OC��p�s�(��E�1�g&��I|���|�]zC��.�Z�S�	$�ؕ��'#��VO�땥q< &P	���"�V0��
�Z֡�6Jc�`��B�y�"|
,"K3�/��d�CR�A����K����ϓS#�v�)�+V��K&NH���H�A�WEDZ�ń�^O����#�c.���*��JAX`����Fnj�S�i�G��7be�
1t���m>|��%�l�u)ZL�Ha�-{�Ck���tĮ�c��.}f�q�Ե��N�$#{�M��O[�)� �j���IW�XV��Ώ��_]�da���^�C+so���v��?g�ߤ|���	?Z�D 2J^^�`���FƇd�W�9�����	�!�U\|0Х܈�c�I��''��jı%�Jg��x�i"z�U�͸Rd���5�6?�?�>�^��bB�T�t4[ƾ;�,�(u_|�����8c���T877W!=�cٚ���7������N#�t~탠-XT��O1�v7���bkd�D��>�J��ẟ�j���-*���d�88mV._����)��0��	φ+��eNS��UK�d����(,�r�ƴǻ��y�{Xʵv+�{�����1h@ ��k���s�!N	����i^��G�T`���,;�,@8�D¤#[�����+l&��U_&����8^�������*�bd���*ZAv^�f�&�����2����y�v9yҊA�$&܈������*��f�Q�7��=DI��=m�xrp�&%i2 �e��l@�nMm�O�lptQ9�j;�:���������������p�O���u�@�(�On��7���U���8&�q#8������,������E�YXNˮ���j���=�m��O憾V�JFY	��c��^8�X�a;pX�e��/�����U{���6�#�#��6�Q�"L)�j'=+��YMu��8���8��Ԡ���f�~z8�9
�[5��d�D�+��}�ѿ?��Q�ǟ�A�Ӄ��$�xԪ�tU.ƀ��� ��d666�:ߧ{�m��>��4ޑ@r�d��lf�@���Q9,����Y?�D�p10rZG���7≕���T��տ��ޘ�2Q�x�c�۔��©�崹�x����ғO�d*�rJȯ秇��/[QR ��>���wI~�MH����&ǳ�nH�\�i���5rrr�᱀睌�7��8����i�����Ȏ��vM!�׮�)���uEA�㳖�Zʞ�^n���JT��q���)���$�MQV��AXt�<�.A_^��ZŴ�1*o��?} 4�0���E�
�����������"
`U?��iy���p�2�Xҟ��J�,�C}?�r�=v���kS(O���\��������VCOX�?ݛ�?��ǻE_��j��T.[
]�[���Wn��\�Ɨ�$���궹_r��2�Ĭ���%[4�͐�����}�����~}^�s���>g2�A~E�%|�Ӿ��R4�9��xiYY���XcÇ"�����N�Èe��87(X���A����ʃF��Q�)���4S_�몞��Ehjh�Qғw	���k������2�A�h)�Qt������4!d[����͙7��e�h�����O0:�.��/	$�/���򤢮���ΠucQI	Y��ؿ�}(P�;_��zO��{8܄f�/��)�2�!�QX��Wj�3GO�0�yDP����m��ۋ��h���=���D��4HC%��_0�ʈ]��|�=�л�-��`~���.��9|�d��ɬ��	�p*C�R����'��e��)�a��ΪY;�*���O��g���ͭ���T�����TQ`S�h"���K�]5{��|�S��0�7���	�R;�1CɄ:\e7_�X>G�����d�!�ߋ)*s��3�[���1h��ò���k�7V�{,V���H@���g�X6v<��2GĮ�z�w����方���k=/�'��t�!tWP�I�D���<fq Rӫk�\��ȏaǊPR���gt��a���[r�����X�.���j�q99˸m���W����=_�m)��G��/B��yٖ�K9W�wQ���ΐ6f}ٵ�a������ah�yN� ����m1u��4@,�%TBV�r����-i?�=l�h≡�jR��6�g?�{�I�QG,�4�F&]����)1~*h���U�
i:���j��d�jarL��=������7��~
���Z�Y�J��{IR��7\�������Ǖ*��y�`��ۛ����Y��w3p$B���?#��y�����l5�e[��fl/�iQ3�x���9v�N�o3��s�g����K%�f|��FFV�����]{3��:\���+~���ڎ��`��xP)�"�����/�ދ���_�J؟�Z�%F?`���*~�T�3J'���G#mh��/*�IF����JF��#���]x�
��D�(*�9�1u�r,�}��s1(pf��!���Y��"�f9�;��c��A'zE����r�K�Z��λ���&���@HM7ي�y�섙�1�b���/ר�J�mi�09ض���Տ#Qw�a`QF����&,���)hq������Z�i(��^��H�������țg��Ʋ���9�t���M��?��\&�VZ�g{�� �w��Ⱥ5��*������}�2�k�w��m��%��iK0��5B�x��\���ngP��=�]����w��w�h�[��|��z�g�*�cF}kD�Us��omdU�����[G�굾R���to_3CJq5��x@H�5�Z�8��OJX����͊�.�����G�;�cc�X���	��Y��kN`�Y�P]���d� �#�,-}�L�]�1aG�����ggg��X
�^M�ظ�B���a��7^��_5\��$�Ȅ�k�Q�pl�y��h�,H%_O���ѡl��2�ݫ��ty�Pp?1Y+�Ŋl�^!�|+��k�-r��� �'6{w������;��q5G��WBF�v�(�@����1��D	����?�����݋��b�V�)zb��/�K�Bhd�{ �"�	�n^!��J˄>�C�V*o�n,�.�$D�"��g�*B��WC#>dl]d��F�W��������g�G㜃YVgW������W�~?ݳO~ܩ�si�Mia��֟�����T�Q�ϧ�ā�����ܤ�	�I�[�ֱ��ξ���ݿ�:�&\���i�͖�9EKt�ďbȰx'8;;[짌�uj�UB����/����M�����C��mP鏤�֋Vux���~77����?_�ĪJ7�(�*G�!�����Z$�=ё���/e�tf� �/��n%�?�/~}��孽�c'��B��������MOLn�q�FjUn͏6�;99-�M���s��C�,1M���K�ڝ�> ��+�Fڽq<6��le�7��%�ۜ�7��%3�q8X_O�S܏�4x���ε2��ULv��?���97]��8�+�����4ߎ<$����i���n�����(d_����pk���u�6ŉ�����C�¼���Y�N�=MǷ�����$=�x%��U+��W���l�%���7�!^X��}�d���H$ɤ�G���{�kjѳa�Y�47����n�;�aq�&i�ak���Hg+�����j�,�m��4텶,����w��G-���ҲK7��a\��uQ
՘�Y0=�#1JA�Wm,�t��������T>�ѭ#���&�'lA��N��������\U����,,�>��y���"�Zl<r���f��(Q�DqV�$�G��h�E�u�9�Jk5oD�����O6�s):�~�k�Fhsֆɜ�t�b����wL���z���"#�W!1���ڷ֬><9��o�j����nڼ����WSPyW��K�u/�������R}�������ѳ���+ ��S/�w@�s{�]����-~Ru�p��d��������Ͳ��%P����������7�B��`B������5�Jӛ	�PK   �i;Y/��<  �>  /   images/686a6ed9-be7d-4d85-81e9-18457125bd85.pngŻuT\O�9X�@H�B���k�@p��Kp�C`���A������:���o��{���r� g�������N�g)l�� [FZ\BЁ�О�<c���Jk:�@�;�/�x��$ �������k�a*zʤJ�~�0�Ϟ�Wɾu��
�eD���]���E�=��V�ڵbkq"��NX�w�k�B�"κ��hK�� $�O�����(�{J�>�Ss���S�ܼ�y�m6��&o,=�����C��E QPPԁ@������~�A dddB�0���뻂����T>�)>�������4J�j��EDD���P�"�����R���٧���h�gb`` �m�ܒ+ZL��$qZ��f20����N��|ɏ������Ĥs��z9�L����ཥX}�D�~Nm��K:�_��)�/���oŞ�I����RU�5������}p9ZX��<� 9n�[��9�׻��#>��I��7�ϑL�|3���5���I؉U�����#_cJ��������OC��24�Uȫ	�ʭ�d�́ď^�R�ǋ��kmmmD�$O|J�5H��w.�=�(֦�|4�7����h��Xc��-Ҝ�4���N�Z�wFƳ���K�K��7���q�q���j,X#ϐ�� �f=��q�&'�&Z�,MO�&�7ᅿW�x�v����g�M���t���_�4"��r*���d.."������.鎛^���o�?739h+3��sX(�	$�>���1V*��_�?��9o=	]���:�D����*��)�7F�7�������fh>H����ʮ�����A�������{k��9��g�[�R�JB���]�D�k�W���*F+�r����k��ם���ڱ]�4V�>��/����S�������_zm���-/��G�5��:R'.T��� ��(����ܛ������NS����n�h�����#�G��i��fĹY(ܰ�K��n=k^����ͻJ��y��z�L���z]LL���U�ec�r���0��WB�eڹ
����0����[��������܍��i�mU4�}ZvQ�p�\N�S������6�w�G��¯3��q�$�;��?ʈm�����,�uK�a7Z�m��1��<�-C��s�,�۲�!ͤ��F��u�L,܋�s6��`&���QK��7��9l��	(ł�|�ͺN�5���v=1تd5mXڤs�F��A)��>�5�b���ݵ2�̟�sۭywg(ׁ�Px��-�a�O2Ӗ��_�
�h�P\NVZ��;#2�4��܂��w�H�+L::��� W��5ij_A�R��W�`�؟>� ������Z"���m�`o�*x�"� �튰���n���?�(#�O�?���3^��U#`~��.]c���}�z�>U�,_%m)���~x��(����Lg���C6���J,BmI*ڛכ�)	t�惻#H �\-��a��=ܭ@̲V��o���?O�pbH��:	�jg���sX6����2��| K����x�,,���o���7�̦�B�M�j�|��T��(�5���C�?9��S��Pɥ���Ѱ�v&p����t����߰��z���q�pMN]���cN�)a�;��[��n+u��Q`1�3�r��.B}�S�xJ�_+cԳbƳ��u�O[��	%Z�tQ���"�s9�ό�˧��V�v���)����逳���c?n՝1�W�G�s?��3�I��4G��Q}�yL�JP4�_��V�+�+O����T��4�4.J��!E�(��1s��%��iW�@|iɓO��P!ᴚs<��NN�x��a'BM�$���6�L��)k:�+�zt��֩R3Sױ4_���*F2�VΜK��E��)l��f�~�3��w�)7�"����nZJ��w�x�� �C�h�����Y	�neY�n6�?���ip�@�Y�+Œ`�	�U�������x5}��=��Ql\�!��[7��;E�д���7-�C�ో��+��-�)a�!���
��$Τ�*Q��;�t| �֟�6OU^�Nq;Yُh���ٗe�bf�d�{���$N8���;4�0��2�����>�bu�k�1�\-Ο�A~��#ȩ��v��y�]��Z/�Y��@�3��k��h"���P�֊|n��Qx����WOΪ����^q$����sZ���y6�&ν�����մ�!��j�Yq\�%�K��޼�\|�cD-�+��vw���öв��w{ _Eǽ�㳘*~|�ԛŖ�q���]0�%���?=l��ܬ�g�X�_�i8�ny�\�{�Za�t�A�L��� �g�KCT��i������L��.8��X{���-�,���Uf���r�|4������h:�Maqu0�k����&a�����_�~i���D��GsF��">V�sۜ�P2X��/���G�"��Ⱥ��ϣ�]����v�����z�i[��&�T]����l=���l� =c�SC��'6ǝ�
:�r� �F2��)v}�Ú}|d��I'��U�ڱq��%���(vMﭐ�iY|��Fݑ^�@����v}���F��8�_\\��E�SL��VГ6̸]V���!FҶ>�\�ab���-��[��>�(K��Ak�G�����_sF	���^���9���.�C��O㊷C�ʎ��3,U�6�K@b���� �|{��ۮL3�i�^[���B*o����g������҆=0��}jri��Ã�tJl�\�¯ȡsW�b�����p��4�����Xyv�	��mȒ%���Mݦ�q�N��LE6:�O;pD�j��a�`Haۈ�?�� ��:�����P�['�%v��
��.I��CN�'��� ��_7����d�\N�ήcccGPy�67s���Q����3���1|�=��	ۧ �����k�=Q��� ]<�	��?�,��a����[Qc:÷��L�e�J���{�a�>���u��
����!T�"Dg����oyg�I� @�)+�L�pW���Y�ץ�����N���Vl�Z[w��S%H����ʱY���/��Lc��+���X��2����A0�MI�W������x觓@�r4V/���&鶈w��EoZ�/�X_��h�g괬��]4
d��XɅ��������/�['G=~�6z��i��6>�Ai��'W;?�n�b{5�д�{�-����a�S֍	|��CR:����*����Ĝ��W'�@�3Q�>��'���_���#���`�ٗ�����q<6Ly�_Hj�GN�����g��­��]�'����d	-��p}t�������'X���!R�Ao^!�u,���J|$����N��Y�Z4Ņ���iobvیb���T���VUeee���Lf�:5�(�x�я��]��d�N;�#R�H���g���w#����38)�j�e�@ ����Pg��|�ĥ��i_ӊN~U��ݟ�~�֛�B)*�u_xr�vm�XG�SR�_nomAW�H�ԝV��B8�w�AMVb};��'�x����$�c����X���(OF;<����3�Q�$$'ֈ��nZ�Y��������Ф��o�Y[��N|0,��v�C����뮋t�񣭣?�����WO泳�b�X���7����\-�0�ⱂ�"��-��$1}��7���_�T�_���,]ճч��S����<A��0a�����t��f�<&�G���Yi��̉v��j!綥�p�nG�=��r�on��E��8�4	˃0�����{OO�8t����}�u1bW7�wp�۬`}�D�E%�����Fr���9\�D�?E�W�|8���J��'�]��Z���D��o�ԇ\����-��'�I�5J�F��D5<��Rot%g?��& �Ҙ��jy�߷�L�l�ey�s�,����;Qäa�����`n��Et�lK��efY#K�C���ꀝ8f�!�-{�Wy���P��
@�NT�#	��_�Q�Q��J��%NO;��A։`�PS�͍O���G���B������\��wf\{u�ߓ��`�{R���4��>�}`�����|�t`i��*Na��:�jz�T�LM~;�Tr�	���qWn �u��x��E��ii��a�@)���71���W/�	�����������b�`H �T���¯���n?}|Áe��ᬟ� �\țKޙWV��rҥ���ם#�s�"�x�̾;JTfz�������?Џ����f*� }V�m�*SXX�|*��u�1�� ���[���e�6ozu���d��p�9�GZ�W�-��V��eL~��+�������A��Q����M�I�b�i¼.�-���k����Fr|�tjUd��Ǝ�\ga�������g�=mT���6h�\mq�����OR�����`�ͻ1zr��4'�N*�b0�ao��G/?�v���,ݦ9�K���_�9A�����s�1pY9��c����5�{,��;��x�)�ÿ�Y�j�g2M�N���g���)��`��ZO���<]żu�lPsYޢH΂����0}7����F��*�RJJJ�k��RW[�܊��ݵ�.�)u����A̬���}b'��#}�M������a 7.���U�u�+���~_dQ���\�!����Ձ2ь1AD�$6�}�C�C'���(d}�%@�Ej9xo�G�h��[}o�� �m)}k���"�N�=�{�{.��{��MYA�}�n�b V0=.vX}vF2�afљ8�>�\��i��d�}R�"�u7��(wUaԍ5��J3N�Ӗ��K���x�<U�"/�P
�����bw4��7����v����3-���
et��,�f�9��|���6[�n��Z���`>;6��Qŭ�T���ď�\�xKJ�������P�Η�%d�[�z�?&�����Փ��X���E����h9��kC ��K���X�q+��;用oz��~��L��� ��M���w5���r�\J}r�6�CZ]Z�EJْ����^�������-��uOuG��E�¹(.�{�5G��i2�������B6K��<jq�����U\��1� �����E�J�3�,��-�����Q.=���2�_��=M�ԙ}���Ҭ�!K"��~4��b.�}�S�O%�����J��f�����k_r[��F�=��1ul�'���5��c�m ��I�mW|���hք�Lޣ�7�}T%ͬ�VA 	���?�	�w\]�	�/|p;����[�s�HCqy|�Mժ���D���#(S:�g���T��H�N�Oi�Β{߬7:�@����/+���W�q�f��˄6�����7BZ��o�7J(�zo�p��w>SdZ�@�]H�؟�zW����[��d������m�-Y������p����Z{
=���;@��9���T�y@�|?���@��p�b���a�QuZ�B\\�?��������f�~�9�M��h���t�?ܞ�EKn �г�*!�Z��p��.�\�M�[o��K������u� EqyP�j�q�����Db�7 �;@����f�W�2/���r��#I�=��o�0*��B)X����1��������ȿ���\��#T��g�ޔA����|L��WLZ��I/��!�w%���GϾȫ=oĊ|�c8g�pHh:�~�j1��V�IS�-E�,XF3����g6�Rt�M���}55�t��W��V�]OVpx��u^�l|ўcLAlS�K�:]=}�MwZ�u�/��¾������@Y�x����A�j?��^������4U��(Ѭʻ���4*�#̃�0�H���$f�e	���iY�>�f
�O�g���=�f�a��/h�8c��VM*�F�:y��$soTj-ҿ�̛�����NƯ����έ=�f�U�G��RHa���KH�1S]�G���`�1��m����h�OԑR8$�[��fι���;$�e4��20;K��j�{��L	�K�o}�0�]iu��rҬ�w�KN=��R�9�08L֛n��Usa��j�v��|�8��ϧ{'�;T��U�a�,�q\:���ۺNA�� �%�t�Oc9�ر=���ɛ�o;�_�:/��ά�I~�8M�����1����������Uթ\�;��`�a{��ը;̜�v���8���zEH���Rr#�z��){9	������� �v���Gڐ#�J"�7cE��O����t���⏦:-��I�2_�,iN�� "Ů��'���w,���~��5S��ޏ�j�������<��,�jG�����L-�r��g=�,���V�U���#߁@��*�>UBO�BҮ��I��\9��~\��Ë}uF�)I;��R�y���y@w-�� ŽL1]�xw3�����XF܏����x�Q5R��5����	G��`�\�G��).:So��t�:X� �Hi�1��L�"&XD�ֲ&�cmu5���=�[�z
���͉G/b	����m!n����>3(���ygd���8��&Ἠ�/m�{܈S����t�������־F�H�d���հCl�+"��g&3]����������gJ�.vF�+#����ZLH��˃SӆN��~(�'΄$�Ж��p�/L�|���*!vF����h�m����:��a��\����n�.Խ�Ύ��@��8�����U5hY�نQ��X�MuB��(?z��T�EN�2���ed8�MO�6��J���cl��[��o��c���s� �X�\��2��K��P-^t<	������oU�v3�n*<�����i�ѩ�\p�nJ/��r)X`_���A c*E�ˉT g����uc����i�B>�I'R=��F��6��Ψ;�9]jlɇ����/ǀ�����+��w���dx�����QS	�ܗڒY�����Za���<oE��>�W���7��wL!��R�ֻ`1�ׁ~~~22�EG�oT�*a��4"�dl��K1ۃj�Es�`y��g\�y����*��{����z�*S�=����o/Ԋ� 	ԑ��WU�H�z�u����Ȍ�N��i���p��90p��Ow�_�m�7�f�	�k��nZ��xLw#�=�H���QG��O^�x�yY��/�/v*�r��7����[��yܞmBF�,���U^��w[S��[~8i�<,�������g� 7�j�K+dB���@;V$Eg���Hv�5{��@<�|��Vi�o}���%:�B�-z��0�(x�z�,����h��~����Ǵ^T�Q�V��z�bkyZ�apK&N[ȩ�b�Z-Ԛ�+[9Z�z9v~�F]o=��i��u5���R�b��%<�J�T|�YЇw���/�iw����J�X�gd'5떤z�@��/�:�Ջu�Ju��!|�
11�����
:��w�9)���A�Y0R4�V
?��+���&&!W���2z�T� �!P�ߍ-F��Ǟ���	J5��YA�����7u�R�������p��#C�����nߋ�R�֒pMl� Wv�V?�ǯ�m�x{�������AV�Y�1�@⑱�x��H��`��E��L�8VSK�9l��VtZ��2���{��mdbbr::�G;������ ��*@x�b�J����B���~h��c�jSP�ٗ�?��}h�o������9JW�0Ը�&2x�G7+��HH�p��hY:�cO��/8���X�J�1X��ctjZ������(��i#��!�}L?[�K����x����Y�`|QИ.��������_$�O䞘G�/�V�Q(h�n���k]�9,jk��z"����	
�z��9��u�������ׂ#36�k�O"�)��b�����=���M��R�XN��d��~�d���L����	}qc��MB`���+t�����媞7v�\6���#����"��|�7�Ā�^7��t� �����#2��mll�3�ת��������A�A ��;lOȨ�R�2�Y��X�yvVR3(���K��q(d=`U��E+����f�~!O�M0�"Q��1�6��K/�>��m�ì@��@#�w�,7ْ�t�i395QG,pOI�L���O
K�;����p�8ȍ��&��ƾs�D��z٧,K�ܼ�I�+�99ܜk.����K����-�4�%��&_�N��l����+Ё���w������&�XѱO�P*n�NI��Ⰵ�)����"��@P��MR`3��~��y�I�ʞp��+�zv<�M��X$��:2ֺ^TD����2�i�F9f��Y��(\'�� ��������&:�_��l��?�i���~���k�Ƣ;8�4U8�׹{%�ы�E��mXT#��#5��''��e-�~����g:Uu�~|ʎ�s����m���e�Y! ���P��8'�Z����2�=H2̚��I���D��ϖQ��#����Ֆt�*��|sE�U+���	-�w�h+	���)�����ClZT:~�bXw}4�ao�3%=Mk�|�׮#�B�G��]$�JQ1�z��w׳�W�Wp!++ˉ�/d��^;@k��җ�d)���+��1�d�a�3�U����d@6�H�X����b8KY�L��nWΜ]˱4_8��Ǽ�w(x���j��^�HS�U�{��<���׀&��6zbL�ala�1N�Ǵ������>5�j�8d*5�'ٮf�����`��&����Ҡ�d�e����3~��c��ߚ�U/x�aeZ�H'���I1b�ڼ�l<O>`�{��ߌ�����.�v�V3�
sQo��,�	u�Ni�������q���"Rɯ)H� ����}�X�J���sPb���)��&M���?�w.w�N���q�3�iv��Tr�n�%e���>������yr��eno}h�W���@���Tb^X�ᤀ���@�9�T^�5׆ 0���J�[*�\�}^q[������Ξ��i�o��ƚ\�$�Qd�����7� q	ry9��N_F _�m���KC�ݐ+���x5Z*�+s�?�Gȴ8y{Vݧu�ϳ���8m��"���l&�?�;�`�N�hf�U��z,��<���\޾̻�*�N�[+}��é9N}������WDK�vR�h���
C�f��Կ9��'�2&ECz��"G���)o��={f����m�1X3	u����IA�3��z%>]���/��IϽxt�M�	|{�Ȉ��|����k\q��J(T�}�!�He=�&���㝰m.����7wƣ��f�<+�&�e[Z0"��Sиq�-�Q�0��O�(4��^i�;C1U��;��uo1TӖx�o����IfP2"���bӭ����'�Qn��h�+bG�ˏ�Zf���{�\`��6́��.���ʒ���S�[�B��)�@~qԝ�jm.v�5��J������0����)VZ�C^�و�k,f�#$*�n&�ZܩȇʸJE~��Bi���.?��>��Y7��3g���fk�(YLe`�[������6����S\�NbSS����)�^6U6���\��V� �h�f׷^��T�-�3�G��=���-Y=;�h��`��У�z��N�����	�gK8�Y����j{�)�	���N����Q���M��:B��"Q�#��UV���,RW��|Q2-K�7��G��:��⁎n^h���-ڛ��?G��CD�Db�g�0ߺl�v�d.�~#������(
Ñ�O9��t�P�o����3)5��y�i�z�LP�Kє�����%���B`b��`�����x�~


�
�0���KǷ7��D�!-�]�Rd���k�4%���3|�z��X��0�M涞| 7|�7K>��QO7M!k�/+zD�!��͸�Ĵ	lԱ��4��Ԉ��ݪ�ɿȟ�^����Ї�����Q�p3������E��u\b�u�EƉ��fQ����2��b�C��rx��TB@��>ZcMv�8 ��sꪸ(�x�H����
�Z�\[��'����Ģ��_[����0O�I;x��]�m�+�;&@���U��.*�UWU� �ظ��,�(����k*<�;7+�u�� 0ֱ�|��L���$v�<y�o�
oC[YY99���G�?�54qlg�S\��»���!OZ';�9������⏲;( �/C��M��
_�����I���Vu~���QX�Q�]x���m��ӼN-�`u�I\�#vմ��K�z�hF'Eg�Tڛ-�$7�=����6��H�����G�r���{0DIGG��C���{�E�VaL	����ﶃv���I�I��r����5��8F-�_��6Q� Rs�6�ؐ[۽l*cY'2ddd\X(7h�5���EF;o���Hwd�/i<�.Cqn����*�]�\�uc=��-�L�],'�tw4;Qs��3�1��+�f�ǭ
�lI��A�KcXo�(��'��W��u�ෟ~�AA���ӰAO�+)QQ�x��@��]G�6�`4>MH��A|f�cr,���t����F��o*t](�zQ(d�:��*6E��O����3�A��"�J�qck+�N�`n%�}E7f��0&�e(�_D��{6�^8�M��Zќ�m�P�kKI��0�ԫ2�THښK��F m��՜������W8]�5jٌ���L*�7ka�Eh�qq�ڏ�H�e��%�B)�C�A�+�c��N�/����&�	?���0:�|�݆�U��G�ܦ@�HkՉf����b��*��j�9��K\�`���㰝}D�V�ȉm�Ǭ`]t�n���?n���K�w{��'��������g��f�v���$X�3N�E1.`�3�(�x$\�9OS�T9��Wg�t��� �b��\k0V$����4���)$��-.�)M����",�-ۊ��_��� ���9B3����2�{�O�����.hp�g/тz.����b�)+���]k��ߪ�\!,Ksͨ�&R�NH�~����t0c������-��(?iZ�9ȋt׮�e��j~JIb�mpxG�����Ũ4�de�L�a�๞�d�J���}5KZ���f�E�R)OL� �g�=3���5��Y�;�+TV��=��)Ն��{k.����^L.��j�M��3[?K`a��5�4ahc�֐�obGш_��$��6���4��(h;8���� ������z�tȎ��W�I)�d#���mTU� F\2�G�q�M�ŭ�--���:w?�P�����!�a
#��š+gݐ 
�����q�z��8Ԟ;�G�_����+���4��
���c���#R��ӵ?͕�`��k�f�p�F{�D�4]i�Oʘ���D!0۱Y��Y�|�mʊ�1�ʖ]4�)F�U.�Wk���߯��M�z�������I�VkŬ۠�`����1���!�2�2�Ц��C50 �Y/���Q�^���W1����֔W��A ���'c_�g���aȺ,�)m zzu���He��7:|%$ �8ƿZ�������ko9d�/�����������P ����:�?Cp��1��}e��Yg0W"�|�ps�����W/����}D���J�!�e �[2?�� �5556^���������e 2��8�[=#��*��7@�J9�UR�nFu���	�g=�H �஢��0$�t4j�j��h@���-��χ�A8=���܅ZYUe��l�:[�[�n�_�< �+m�sA���LA�h�#���N��':3`����"�J̀�����7�e�J�6R�:�F0�zq0b�K����<��:a/fgg�:B_�s屸���рQu�=���0����djcm������zx5#	��^}z� �PZ�͞����I����ľ���3�X���'�Fi�̦^J+ֆ�U�&)ئ>����ĕ0�G�Yk�UGVx�_�B��\�R_��3N��lqN���^����,/4	�
$#^��T�}Ij��*���<r�����������`S�g��*��O�2��5ric��І�^��ʛR��;5x!���V3,p�p~�H&��(DR|Py8]�7�uw�)�gQBk���|w����m�<ҹ�}(Y��׆��/*��H<����]��y�{�]o�Z��U��B�����#�-�P!p��^^����[$F]ᷴ^���S��=�������C��﷩[���Z�t0�O`R���=�=]?r�?��O�"��r��A��Ax=�wg�����gx'k��U$�x+�s���5��xQ��.9��s<S��A0����/��V0
�e���@����+�?A�t!a1j?��P�gN�����ٮ����]v�o���!%Uه���āW�n���,{��i[�o���n���$whq��%�3a+�z�a�)�ըK��p��:^`���m Q���/_O�����l�)P��7A��i5]���)}!�,j��E܇�� �}��n{��E��|�Z�`8|f0�t���$-�z�8���d �@��A��t�!�w P��p^ݶ��$�kF[l��R�QK��La8@�46�.�_�ԉ6e~���`|}��>"��ɪ�����oy�)oL��3�ާ	 [�ъ ����M�6��<�!����])���4�Xk�aҭ����'�<i%T|��U����3�!B>.��`�﯋[�iy����>�}�bw܇p��?�-��kv���a����*v�M{t�,U-Jx��f����b��qu�zs�u�:L���j�ǣ�jI��W&3�V��B��\Ӝ���䵄sI\T�G)���j�&w�dw�T����[Ï�|�v�L&�B_�	:�.��E�;��SKQ��`�V����2�[���:���5\/?Q+��@�E�T������f!i>��-k'��)=a�A�hc/���N.�8�vwY(vGM��U��hv�]7���������n~&��Y��`��yف��W��%f7���
�iBн?ES�?J�S�����y>X-$��7?�m���S���t@{��3c�h1]JZ������Pܟ8���֯i�v[=�M�Ԫ��W�=d��zwj�6�G��磅�s"sF�|�B�n���5����ױ�K�F@9��ok&�8�r�-�n�N���]4��W �xT���y|�]����N�cc�L����0�32|�a}KjY�՞��9R�A��I+��L���8�O땛�̠&�&EϦ�������F�Ӛ���j��})!��q-����0`��ݞ���*[~f�?��l�y<��dw�4x��n%�pZr���.%���G59��J�$�i�&���"Q�&&$/�`@��w\�rќ�5�ׇ/�A F�v3�ڹe�`���~�K<�gP�z<�v���A��I��`>����\���y�X�b�>�LGQ�����k��>Efr��h#;AR�+���[�&4�������$�\;���_2��bՋ�}�Vu�*;�uN��pl�fQJ�˳Q�gEg����׊��%3]mO��2�V� ���;y���;���c��>A=���ڿ���j"�;児�k���>	���dJ�l�?"V ���b�ʄ���s.����V�����������^�o�(���4֙����ѽ}�q�k���tV��ۦ]��D!e���w��o�E;mh���s�m	���,�����7�^K�_�O�qYt�yKT��|���B9��>��c�A�[��p{�:����_�
�}1*%��~_�'��k����b)�[݌�F�vyA��+~�3TY���&mr��T�������ɶ}��U>_�o����O�Iɝ�j��<TB�Զ�,9��H��g���
��k�i�|k䏛��7��Mڈ\y a68z��S��r�I��1�z(�g���1��ikQ� ���}��/�}HZ�tDo��E4�,�� ������hӯ�\��v��f�(U�k�Qv��\�K�f�^aX����'�X���d��e�Ok�<pE��Y���c���H�)]ٖo>��l�����p�1w�G��a��iha u�?5d��[{|U���~m�D˧ !T�|���,������װ�jBR��E���m����1l��S.�.�ot���|<V�r�t�ϗV��=Ü,�u�V=��ZF]H��c&�Cʅ8�\I�|µ��.Ap�dܷ�f-�����U�_
�e�W%���w��vX��=]�T.�ۖ�0o�
�8�%���介�85Kbu�~����~0��[�� En� ��Ge�Q�x+��2KjA]B�t�����t���T�$ǻ�{�|۵�]kY�ˮ�x)p�����ϰpf�j"m9}4[���H[�\�G(b�*8/�$YO�8%ɓ�"����^�=(������M����2�^-$~D��6��>�Ggϑy�q��u�x��b�pj���NT��mq1���F:�ND
��sD�h`��j�@ct�3���U+4�-���F���}Z����q�zF:�ۣ�vHX���?���_2;�L�imY�Nm�E=��:�@Io��=����&q^��i��a�pV��y��*l)��v!G��j�$��1V�_/�;�)�T�������m��nԯ�?͇|4X�SL}8�;,H5����~l��|��?�˒�6<���ik*��`�|��5���p2�q�L�[��UQ� 9<�v�{�L���ȗ �����a.R^^�\zz���d��t8��I��T(Z����}Wb-I Э��-O���n۩$��K^1WSQ�շ
i :���|�䘇�<y'sZM�}�jE& �n�&m9,�i&n���v��R+D��y*�:Y���֕�[`���]1�Yބ������4|��!��=��pa�J�rN�%*��Ia�޸h*ֶnN�QeH��웘�{	$�6��:l����N�{��/?>��)�k/�P�Gj/��m�ug)޾ڹ�ퟷ1��ˢ�N�u�g܆rW@q����Y��{>�Ai�Z��S�����AP�v�������n��'�N�ig<+���u�4�J�#Q���:d`��[E�����5�(ˀ�ɛ��m3R�}u!�$�a����>�N�ø�C���[����*��-C^������ķ��I����2��Id9t:��g���x�Y�,��i�S�Vv��j�[D�Ѧ�'�O!�?G�[��T;nѽ&W� G���#6��_�@��x�����KV��ؿ �d$�KE���PK   �i;Y5��s� � /   images/7b4f3c61-861a-43c5-a680-e3c3f7136b2c.png�eWL-� �	����;�:��-���{p�	�}pww�����ӫku��ԫ����Ցʊ�(��_�|A���P��������;�EH�����˗/���������_�|~�J��{���%�\�"y�Ls�

n�zt���2�h;"@��S������Ɨ$�F$ff��R�!�sr�WA���d#�%��k�����n1��G���uҘ�����S���qL��P�Z5���|������K��GlI�4'��F֗���?��y��z�,ll��C�H�b]�x5��妬��:P�!r���}6�����m��e�:o:���+5�<��c�#&iˤ�z��I�P�H s��s�l)�H2�Ғ06U1�cU����+{|�WJ��vm�.����ښٕ��ļh��I-j�^�����q��}�H���{�1Y���7��r.y7i��.���T���j��p�-�Y���R
W�H�ӻ�U%��)��#L�w>a�h��C��̳��p�HtSԨj+��Q�U6���	 ��	���a�ZC���7��v���w�/��`�eh[ܚ�{�K���O�M��S.��o�*%�.�\p�ѣ^��c�EW�Joݖ��S�磾�2=
��ɠ�!ow:$�� ͑+I R���bz���$�?�GI�Ѯ��[�³Y�t-�(L6Iӈ�l���"3���bQC�-��K�g������g�n\y۹���=�!:�>�F�4�)����cs��nm���PP}���ںF�P�]UL�T�_ȡU?�y�Z�]��a�+ź���}�����f^���N��Z��"0$O���W���\n��A�j�[?�l�U;$��&f���Ս7��k�5R��,ɸPC��7ؾ�.Ӊ\S'�IA���"���5�.�	�y��e��lϿ;��҄#�&	�O��|<k`_S�$;D|���^Ʌa߼[�����z�;�sd.�ʍlV��5���θs��Ŭ�	(�4/�1�����[ךȈ\]ee���*��6E�]{����nd�SO��&Re��&�˶�d<\4�U�W�3Ɏ>Q2-Ǟ���;�A�L;J�¬rN�g�6���{��H��_Jn{��;.�0Y@�;_�oR9�*r�a�r�
x=9h E)g�؇��X�]!�rkZ��c<��V9]�*�d�HH��o�z����:�>�4dMK�(��L��E!� �LΉš��8��%3��!L��,�>�'��7C���� �s�k���t�J+M�J����5J�.�$ӆ����4�I�g��7�%��&�\���cJG�7o�w�M���M����s�kd3=݅sӮ�_����K��@����F��y����kK�G�ó��.;a`��`�6�bM��:Y��������Xm�#��ۏ�F�-�p���D���Ǚz>/&�U�?��5����'��j��u����\C㒤�5�=m�{U>�Q�����)�%�L�;��dN6�.{��C�1�Ӣ\v��|.&�oÑy�� ��@!h-���js7�<�v�����P�l��3KBĿ*����� U�ϏgJ��Cz��1�%H��칷"u�j#��8�i�y�k(�7�;��a7�y�KC��Q��#hM���׳�t���ȯ?/:}��<��r�9o�\~�|��<9.�℠*'��kk!��04Q��'�^�a~�.W��jU�J�L��RFa��>�c�Z�5��Ol3�Q���\�Mz�$<��)P�O<���!f\�:v�%�d4S�4W:��\+mx��:�13�{ۭ��މ��T�x������ۛ���8�R\����&��q�Vh��WB� �}����v����:��\���sw�١g��G���!���6똃�����U<!CQO�Fw?�e�q�������}ˏd���;��1[K�6��w`�v���(��Q���nV�<|aT������
�3�@�����!�e�J�J�K��I��[�s?��?:sU<��H����VI��8`�"�M����J�V:��X��r-�E\S�n���qJ�����d������nxd�Qo<�c���������|u�j�GOO���9������d!�qgbZ%�DoX��b�6��!6�X
�=�
Uϳ�$�ά;fQ��FRG�Э������T+c�Ok�Յa��e�D�)����^������i��ein��5�+>D�)A�I�1��$Յ��:}&gaǵ ���(^���B�^���8S�����@���w��P�o�^��5d8�HA8�+��"�*��FH��V����H]�Ғ =�����w9�iY��~X[y<: �v0$�#�� &���9.����_���)(>�L|o�]:R?FGe;�v���sqpp`V,�������'���CdwE�~�|�g3^s�# �Ȑ�w3<�a�ne�z\m[���A�7%^�s��<v[�hֳ�CB���[iY�M���"U<��(P7QB,�1_`���g�`쇅��B�����>���4���[U�>�1:lIց�������'+F��~}�x�8YR���E�����Rc��X[^\��hni����ZX�^"�z��=�o;bCU�7{{�?/���������qA�6���?��)�V��T\\����u��:_�/KJ:���.f�C���j�7A}�g���,��xbR+�e�x��N�������{���0��&^���/��݀�P3�F����@�������f �v��Z�o�K]X��`0�N��p��eAf�K�FS|(�Y�~Z�:��+mX���m��v쥨���H�X�A�k�>b���-�M����US�����O�o�*���� �S�����k���񩬮��:��o�5=���M��ޖv?[朆_M��Z̕�S�����E���˩�����^-�(�]����ZG������3�.E�O�!�d�ڀ�r�JO�BNs�Ԭ�!f��\k�M���I2�H�VV���dA��66��R�e/���{bs%u����Q-�F@;��F��F��6��RS�Ě[�<��ME2t���E�#a��V8�0�BӜ[ߣ�*�X}h��>�y�/��w�9�O�?<���xU{�l��G��P�Z�s訲{|}7����[:��<ĢJШu��ɨ���J�#����Y>�w*�y��6�^eC��O�\�����@w��^i��ȁEǕ:����Q|]�����Gĥ[mj���oN*��Y��!now#���S~[a۾�.��f�Q�&&f>!i�iX��%��� u�����s�obb�1��X��:��4S�ڔ!�*�j�^�z91��<�%YH�9�Q棼���y��@O��l�cK�7�+�#K���&���|[���ΣU�5�ʇ��jm��)��?K�;|u�#*�m"
�J���x��@?��>�I�<���ȯ��������o�ht��{C�z�^�|y:%�j�X���
WF���=z�E���?V�;�z�z�R-)G��
9�n��mث���^���s}$k�D����/������Mq����K�Q2�|�`�L�M���9�Y:T2���#��w#ӄ����GB���ܳ�eC��j���'Ն#j��$`��3lƮ�����;� ��j�1t<l�k����ѕ����[]dy]��������*�d,T՝W���Օ.�����a����|��HMM�ΰ�i��r��
�HB��/Ѿ$�C�����D���N�vZ /���BD�������#Z4��
qȡ��W�N��k�M|������C�ǼZ�ݕ�Tr��Po��D:��,*����������"�Q"�*�b�Ey��o<���i~�X.��{�|t�a��ԯ[Z��BBah��Qol�*�ŀ{�q<;��cbrR$usoU�K�!۞i@o'U{���M�l3�l� ���
@�3[#$<�EF&
���Nn��D��k��#`e	�ٞ��7�kg�c,�{?z=J�{�(|X���lrDQ����Nݨ#���ȭR���_8���Ka���Z�Np�^	HK���lR�V�~������U�/�q�u�˹O� b�����
��"j�
ӘpW�r��Ev���~I'q���hz�B@���|���O���K�{�fn̿��2<��cd4~�g�Ϩ���+_�Z ������f��^���V�י�N����]�������z���}�.Tk͑�~z�»�C/-λA�� �k?}�{�����#�Ǧ���n-��s�m����6������L�o��R]���S���؈a5��c�.�&#ߋ�'1�oNo���wP�Z�"g������(),����ĒBGm��R�(�?�3���h�
*޼�z�xU��+�غ�z��r��;�ʈv��|lg@�L�: f`+��[7!��5\O�I�>�XH~��;���
��UA�(y����
X���^*���^^8>c�@�eC){�mz��r.��8�I����Ø�fLĬ+ˑ'}�rϞ7��MD4��:z�0����YKH���/H��<kjw�g��hR4�.	�};�OCgRf� ��hΥ0�*-mCRp���+��M^�B}���`c*��Z���E�j׍�uε�u��m��[���<[V)6"�>�5
fTW0����q�����AV�(Є������:|�Zyo>e�]T��%��u�(�ѓY�Y>oñ3N�c��Sy��Ԋ9[[� ����.K{���y_�5zdf�US$H-z�S����n~�EWs���tI�c����yړ�f��Μ�B�����t��{�jئ�0�ۭJ��f|\���=�ݹDv��f�e>*H�޾�	��O2{�ۉ�Y�E������-�pJ�͐�V����ϭС�!
��-�;|&i4��H�8�������5�t�wT�_�?1>��o{y��g�լ��2�&{xxy�`3�C�r��<�d'Yh���=��2�R���Jc'�ݳy^}�e7�o��c��0��1�~���y_J*_&�����֘�A����|���0	��Rk�V��8��/⠽����o��r�G����f?����gJL�K�G�U��\.��OF����B�W7���p�ǭ��)�>~��AySHFeVt�
�T��M)'vj�=�Y����h!3<Ԁ+��}ٜb��W3�'wv���^�V�>Oo���k]�u\=u���!L|໻A��p�􆆆��p��-n�
����˯mZsNc���Y	��Y[ƭD;^BQ?���)��@��)�*J����t�G����6}�	��Տ��C>ݏ��N����u�mNu���k1�,n<2�k�kaJ�xWBbu�\:�;��<��c��{	W��N��ݦ����Wi�C6�Q�W�i��<}��<[�'�������dH��{�SJY�<Nk�� ��y�����僽ZȂ��[�T�3�|�Q� ��h�V8]^��-vi2��b�|����P�'Nf�F�������!�W~�����r�7���wU���9Ţ�o]��9�	ʺ
�j��ș^;�����
ĸR�����d�N��Pkbw̊׺:}��.z�VY &�6t�{�Zz}�M�x"i�{Mn$Yq��������5ެ��ۣ�~M�<��Q0@�n�g66E�������p��$]�:}`���dJ�ǖi�
���Y"�{��[j�^�v?���\��jc��"�z8;��"!E2d����\�1���T��Χum�?C2��;���.�ԌJ�(�MxS��}=�p��v�i}�y����(h����s���Z�Y��ʴ9�
tpʭ7���-tn�R�ք����_�C����'&�,Z%��mfLވ3���||���5�y�̟=��ˌ���^����4�a϶��#���hge����[����/QǫL
㘤_�i}4'4���=T�"�����դ6(ĥ7��%eۥ-t�-�b��W�pI�W
��h�_�O��_l���9����.u����U��	m�)���B�}���d�Q(�pmlￖ��{��­�"fm֟�T�3�.�ҟ�}��n˲0���>�5I�����V���V���uuu��zJ�e�&77��v��x>�w5�^�w�w��]qӡf�ֿ|_�&�}퇚t��gyE�N�����dM�����i���{t��S����+S��ȕ�c��e� ��l�Z��ʻ��}�E�l#��^���)Oy�0��P�H����N�O��ϼ�U�D����Z�W�W�xm�O��c'VS*,p���,t���&+/�2�3�0ph��I����)��b+��$���PPTlz&��\][C�u�7?�ܥz�<>��K�ٍ۩��*z���t����x��v���ld�}fc���0�͌j���K�a7�"v��D�� E��
6�S�6b�~^����l����"47]&ZR�=�̦��Tz�U�1${�''��M����%�8�\BkwK����p[݋�z������qB����ج���S���Z}�I���5�Du���?�^	�8�ʣ99~}P�����8jĦ���-M���y��蝮�q����z��6X���G*2?H�)�Ӿu���U�k��tsf�_���՗=pOהM�ߜ�G���҄��/)j?���j�d�e��v�:wuO�W������!�)�8�s��Z[al�����6x�J�^"_bqnp@�Z��XM�jz@��p�W�oC��:������(�d�Gd+���9G��V*͠ȹa��>�X�lrM�$�dу��Z�4����޴վe�s1N/w�]��k�d���^�����>�h�}�M���%n�
)�7=itЕ/�yX�RzI]Kk��z�FU�h}����z�fLn�Q�>T��?|o��NKO�f�Ա��‖3�[6ll��/`��v5W��i7؄��&��(6V���i'M������C�m�������Pv7n���5c�����������53��X:�?Ŋ��M�W�-"�\c�i2��z�{�9U��O�<Y��u���x�׆g;k��F0o!7m�F*K�`D��K7r�[y�?���.�b#{6�mpb�Z��c;����S�I�m�029��RP,�k94d��Q|_,�DT�<ԓ�¢L��kn�����fl���ˋ�ܼ�^r����N'&&XC��#:��W��M	��x>�%��0�_Gk���ܼܟ��54�źv:��]��dx:Y[�:�n&�k�k�[�+���1�g;i���U��5ǻ�yyJҖ�Թ:::�]��c�J�o2Dιx���q)$$�-�g��ѥ���.R������.�?�ę/j�&HjVZ�9����Ƒ-���	\!�pG���7���p�C�/�<��f+�щת[�8����b
�W��������5V��y��d��n�bu����愂Me~ԝ���t�N%��3ݴPo�Օ��Z��^���Bn>������l���Q�l���7Ы���}���~7�����8��v+'�k��n���.�-�����,������XVf��Ѳ�/�;��|�K��Г�|!ʢ�����155Qp�*L�'&����������݃�ēJj8x�������WHp�mnjI��޲d�������8^@��kf�O�ѻL;F�Y�~�r�g(bτ޷T��K�fc�}��w�۶����9Œ�a�֡V��EL*��d�%Dބ�����[I�a>��3*+�H�X�py���.9��ѵݭ�h�c�|Y������\�Ħ���~�'H9�{'M�G�ť^i̖CFJ��(����`�e.jЕ�Сh��{�L����*�R�����0Z I.+ _$)���(�8�/z���e��U1���S`8p����ܭ\��[�m@8�T��:y߀���i�����6��Wd��Z�OI�\�m}a�<\o�}X���
��3��e�1Į��M����r�q#�y��ϑF8�<d���JJJ�rhϊV;A���-�KO�oNݎ�FF��8��a�u7�'�������dF��{TA+�����T4��3e�'���$� �(�3V�������%Xd
V�]|a��a9�8J���Y�- [�*����ȥM"E2[$c'��°��f�w[I=)M�skD��m�����m��X,�}?��WV"ߛv��;m��r�� �=}�7��B'`�!oܟ�,<,�����y��9� �)�*�-�p����Qj�R��0�k���)HYJ�&Y�CAIi���q�5�G,��K[�p�A��LnF�֗��kQ����f-��E��"{8eA�lO�Y���u�2��2u}{�>�Qm����]��so�����C!��H�:��y�.y�%!wu�ӑo�Q�"��a?�����UBCY�ƥC�-��6���kzt痘���=�~��T��W{�?����p�O�\������epT����m��vP�sm^�9X�2��G� �����ҧ�T���Ð%��&�7P��-p ��q��q���{���QxDt:M��w�z�QA��՜����N�4f�o/6�/k,�\ ��HeM_�-r"��
�*�R�D���a4hQ�Ż$�NSk"޾����M2{��>���f;v;�rJ'������>��� �A��6��3=^o��V`j���P)Favp0%�^6�Ta`O���.>���6ͬ��vr�Q篧����{���_�(��֜ߓ5N�� ���^�m͓��Z���k$�i;�S��~L�(iQ#'Ls�emy�iR}��{^D~ލ|N�?�>w�sԱ����t���c��<�ק&���2���u�6)�l�$�5Ͽ�Hk*������Us/�7��K�
��ף�o���+|��/�e����q؂��C���tES�L�4-��`?���̈��k�6�D���f?�}t ti7�kMq$�[�|�w����K�6bTn"w�?.4Y�Z1ֻ�4�{0�������/�u��tΡ��!D}\��O.��+��Q����P��m�����IWm�5���g���,|B,���,=X�5�z�g,%��#�_��o�??O]�.>?^�@B�hbz����K�s�����%��~�Oy�-�r�}�8����n�cb��'�xP���T]��ȫ@���pM�� �+����k�!(]��f�z�k����M��7ʶ�5���kFP;J8@�do����x�������`�lPUS��6���I@r��;�ޚ[I�ì�9�}9��E#{������kK�L�=,�E�&浕�������蹅��Ͻ�-7���Ѿ��٪�qP���F^��ڜ�����y�,�~��!,z`ۿ��<��y����+A�]:<<p���Pc���^�2|�ՖM����G�?|���p�ď�L0#	>����p����`�"�O���F
�`�11�V��~8�d�z�j�S)0���jK�]X$�ZZ��2���s����6�B�+*�lȢ�q�?\�2�D-��~��)(s��|�#X�~疃�K�ٰj=:25Q��(=���X�IEȎ��%��v�V�<΍��EK�o�ꏿ[���z�{HZ�4|ߋ�?ʍ���S�T�"�cq��&]�����P3g�߸���:���oG�v��{�cA,��y��J^�N��r*�2Ȥ�t?�X��zuS�_�C�
�kkk�RS߄X'�+�&w1u�]��1tL@��"ܲ�u@��>��x��B�w01�Q��E�'B7�nF���?���Y��p�&`>�q�Ӕ���e
��,I��҂�怛�Ė�%x=���0��4Βz�eK�N��(��:�x�^"z�E�s�n_��?oy��h��dZ�n-�� �2���tR&9�t�.��9�py��d�z:�|�'
�
�!5�JII1��Y组����#<�~y]��l�Z���,�t7����Z���ʂx���9߾y�q��1�Ώ���=��w|�E9x_kQ�D����P�#����-'C��>P�Κ�fo���(W��/��?wܼ����'j�Y���x��u|��1V�����Ҝ��>T�[��~:�}�xdy|C	��&F���sߞz)��|�N��[$哸��my81'8�?'��Ͽ�R���"����#�?gq0�+��)2��\����z��F��aonY��z͛���ʒ�^�^a4���ɜ(����Z�	 `����,Z�����͞��)�kO �/�N:�����5��:����>:::��j+�HP��S��%��Gvz����sz�{����b*���z���7�x�?"!BJg8�#ϒ=��z̉[�rM������i%v�L� ��Ϡ)������^��
����v�tQ�/��~7�J�=cjnk����������ʔw��v��}v= xq�/ d��q�=,�>��V�����	����q���wo���9MR�hۮUk^ع�SS�Q�&�9]�Ci7��v�K������C��)M!��`�/X���6�w`�篫���g���G��L1�b�A��ĊN��K�t�_=!�X�0q���4�/�X�O��5)E@G�K��<J*���DM9�"A9�'81�ǟ"����t��7u������A�g�LA:I~����,n�߀������o�F
�����`׳#��fk��͵5���z��@���h�����H��Q�T!ܻ���jw�^��
<*���d:�1.?�Kfmt+7b�?�`�%I��U򋪎6]FC��r�?�@o�)����=B�s��%�R-[��L�O5�ŹcXj.L#b����xY��&�`X�����ӵ3�PA#�/�Q����W����n��ا�_>x9�\��j��r�����)3��e�J� z,�����Zw�-�!�ej��z��3$Gq�0b�ߜQ�T�)���ZTt\�:T��|tG�e�Ri�[�KLsGG���ݒ���-�]���J�����o�9��L�'Y� �~�|�[_j��<9�2s�Q�f-�'�< �jw�Q������^���J�C�q��k�X}�'�����v������+���m���t�G}h���++�5��e�?qm���^;犻��z��}���62B��P	�#Q'_�'��i�V(�ض����ך�1�FBȡ-�����C�f���]�h� *�}i5_�H�h 4���n��!����(�N�m�\^���{w5��X�9�c,�N�ﱨ�e�����J	����Yf��c�h=�/�����K�5�B�V���G�>������/_���~�,kf�_�V����n�,Vfn#)���Ko��-=ʜּP��:
���k�YJ>-��V���¿WW7j��Ή��5���/F2*�z���B������?�v=B�k�0�>E���鵄rF�oz�[��`W�6���C��Cs�/����.���P|������!f���O-9��N��z��rOK����8hW_��d�I�|�V	�?\l�32ڛ��@����m��l�{�zX;�����N�7��=�7[B��M�������Q��Q���H\E��nKm��6��y$=���X��{�fӜ��6�A��jJx��^�&%"�ԝ�Ծq�'�V{����k��o�IM�
A�qzrB���i�~��Dj07�:	�E	־����U/����v��Z� ��{���kp����O�f[�;�7�q�횤U)���_�;��&�������5�&:
@b�������M��t��o��I)����x�n�W������~:������O��u_�]�H��]�Z�O��ᬐ��]�oAl#��aZMIP6�٠(3RO^μ���z�8eh�~Lv�q�d����b��6g�"đA�V3��?Y\�J��_�n�u&�*�*�PV�Ӊ�ͱOܤku���{g��iT6�e,���%�p�ml�U�αm�.�'o�vG&�^=��T�e�QU���J��8��x?��ᱫI�Y���#�o`j\`ҕkV~i?a�t	m3�>�7�2Cb$8ක|�d��\��!	�����Dd�c��+��*�yؕ�C�Z�G2S��6a�Q�֥���#��$Mwo�k$؞�w��&s���[I1	>��J�<�����%hhhA��c�R�-��-�K&��PI��ǲ���F�d��m���$�ƽo����mB��!*��Vz�݆���Za�,�|�)-w�]��̖�0��Kt`wL\Lw����3X�H�����-�+���L}�{`�æRDF���򨦌>J4Z?CgӖ�6]^ ��Y�����ѣ�%��a�BNL��jk��$죅������J�d^,���Y�舲�\�  ��r�z�e�dQ��Ri�Ÿ���i	d&����|7.L��i��'�����C��w��cb��;(�"s<�v)�:����~'�۫�8�i;�~"���Q�1K��Qr�`�H]��,>��%+�Y�w��Mg(	Hp��~�T��������PZ[��_���������T�$!kmy��+
�Sy��!��O���9��Er�R��2s�ҠM��q�6@�,?kqsW���������m'�F�݃e1%ʅ,-I�o�ؙ��~��qزgڰ�:>�<n��-ˤ�q�!n&fG�n�O�ly,-n���Y�V�f���/�X��%��Wwe�I�[��t��!v8�RQ�WR�b�+�-�r��#[!)�맨������߾��4W������iv��Q�N����c,��js �|Je����ۏ�/����n*$>��P���
xiǀ��LW�����8��)*S��|����)<[-V'�c!:]z;9&\;C�Ý'O@c�G�L����.���|����=ޓm{|�=�x"��6&=�h�L���f�A<�����ڮ{�,��ǜX��b[��	wO�hl��B�� ��j��A�,�P��6�'�n~����`��\���-u:�Y���][z�Q�Y7�G�s�.~%6����-ފV��qC;Ry"�!�p����K=�1P���~���"�"T�+,/�nOqq��tX۔߇����s��6���#ނ�`�T��L��ZeM�8r�9�?����)A�����I-�_���a#;�S��l��B���(��d;���#��0����_����~	��6l0W�����w��/�k��5��yyn\B��Lȳ�BE��Jr R(�U��ޞ�eS����G��`A(]	������0��#�3���)�%E1pn��2�v���!ա����DS�s�6q%�[�%�J'L@���8��cQ~Q[|��%Ҷ��k��.,:��z��S�Z��ؼ)e6�N�� ū�ʨ�v�SgZ�����C8{�H�	F�?�bZ;N��2#fN�d�n���&2��t2ɿ�f�������3�5��ߡe���@h'(4��(�q���Y^� �5��U�.r� q;T�׬� ��o$v������99��|���B�mx��	^�Α�/Rx=%��`Ǥ'�ծ�34�G*'����Q5���gHZ�,�SNLU���%i�0D�E_�r�ޏ���ښ�ںH�M��*I>ȸ���~a`�14B�K`VZ�v�Τ7�n9�!��Ӆh�?=��'u��$V�R:X�Ȟ>R��100�z�#�*�W=�Im���~]�j�|�q�G�����"��%��~<W~|�)�|@�3�QT���-�N	>t���\�hT�5} ~��K���Ag��6�F�1	R��yݬvy`��s}�D�Wz:9?/�����}Y�S]�$�����A,����C�uJ0���W�{������]%n~1n�'T�2�W-h1�(�h��㼚��ף5�W.�糺r�1�]%��W�0L�L!{�yy�7��o�#�k�jȅ�;�Ci��  �o�����U���91-fgc�f���� 4}Q4��{�ꗌ���W��v'�1Q����$0y�ɩ4 �� ��l�<)b�:�E�R�B,���QO;�rE^M
h��j(­C;�f���?��g�������CL	�k��P��Nh)�ԟ�����ou_�	���^h9���/�~��M���Н���Q^��,:�3�j�c)�_�Y؆ߍ���'������2�����<�V� ��F����Y�M"�(x�̱$��tȪ)�xq�1��"/L"�ʧgf:������j��H�vNс�9וP���B�*8��s*�L0z��V��Tqj���[�jkK�v�O�@�ky������_���py���u=�Ш���0���t�~��9<R�7��Wߛp>��?$z��Ⱦ���}f+�u������I]��yE�+�'ƅLpC���.���}Yœ��f樯�d% �Y;?O/����fR2Y�0ӿÀ}�3���I�M�. �w�It���������m����wv�T��zY�. ҟ�ww�":���e��G >�G�_Z��f�B�W���JN������h �2��k*.Wo�zJe��e�;�)���;�0����'��Ƕ~�=���x�����fՠR�
&(4�>��S�9{�ӫ�8�z,�Ԟ�y&�`(�:4ּ�S6�ЂA��L#(iދ3��Q��0��Xg�"�B�VD�WԯR�,+��ʣ!T���'���xE��Vi���ϱ-��� �q��A֚괌!���I�d�)�LP�:���F@��e�Q`����7�&��OqO��|g�l��m��^�����Ɩ+'�v!����1k����ա"/���vܮ�b����	�s[�t��v�%�qg���p���)��
�����]eWg��/�6�{�w1���n���w���f�1D-Fi&Ou/�J�s�=4�=�_�����W�(#�⺟q��k�^��KӡM�V�q��]qS
�{�->���[R��g2��y�Dw�M�� %�x�5���ܿLD�y$
��:ո;A㺘���9l����^�aҵM�7w.S�E8Y/�l~W]wsZ ����V+k��S�b��K򵤂%���R�q������KYI��sc5�$��3�V�?��z{��~!N� �閏ᅋ�8�/L�3�}�CDg>�S�53�-&bߚ��?t�%��&~��G���U�G�.�$EZ���
�&y�R���=��~W<29rj�؎��ܭ*��9�IPs-C&�3�s��0��v�����&Q5f쎷��_\��s�\���}������HF)^r�d��^%�˸���,�^U_����  �������,&���'���v�H�S��#ˍqhse��h���O�kԂ�0�چ�JN�M /�,B�b�^��Hχ���)��`,��L#�|<qύ�#�[~0����NJ-tUrF�"?�`��i��o5�h��t���Át�ny�M-y��$2w�7���ǐ�hc��}u�My:�I��o&Yӗ��iW��0�Rb�؊甖����}�(5����D»�����Σ�R�d�fQ_�q��l��p�)Q�I�n������)��IM�ƍ�jK�e�ã�4�_�2[m���V����Ţ̜��E�)�ߊ+�*huS�!I �;Y=H�ͩ577��8�&�}���O="u��@oR�x�E�2��3���܇���,v?�S�<����_���mlB�
J�R��څ �q�H�=���o��q�e�$�u�������}�Bp͚\4����B�o�w�jJ���h8��bj�g��?Y�<\ݮݑ]+�(����z9Z'��.�D�����j
h�د��ߟ�>�:���K��:!�o�F��NE��+�Y]Z�B�<Β\���el��$K�Lj�H/���l���hBȜH����jy5Xp�����c��3g�1#
��L�$}j0�7���O�	�����p�$��R����4����<��M#ؔn������	�*�,_Q�t
'��mg��v�,p�V[sD�y��`�Ww6;�n��k���:�a.a֩iH݈���M䍮�"	��ćP<�ej����;ԏ��X���%1}&	�Np�B	X��?
Z/W��%pK�� i����B.��U"�����z�/�N/8���ͳxji�fm���n�)�̶}<��O����K���LiR1���f���ˉ�(��u�@  P��J|�E+k�о ������̘�'��D;��]̅\I�OP��f������~h��+��%����a�]���G3E��f�A9x���c��gD=�����)Pap�:��T��˱�u"w7r5��.>�zX��Ǔ�ȖWr����J�wF=0�_��#�.Fb(���$�`H���M��CC� (@׿9�.JY\:#�j3=r�Q�R�đ�$��PXD�Ï1��M1�AhB�\�Jo�}��9�6j�\�ˁ&���M�>z��|�I�m@�0s�Ͳ��mh� ���Qv����e�4�F��Ç��>��W> 8<M_.�����3��koб?���ijK�i��f���@�?,��Ƃ��afCҢ\~����b:��3�����_d>J?������Ҡ)����hYh��ݝt���鳟}Y<�e����kׯ���>�)q�G��R���з���&����~��;JY!��e��N���_䩗��6������^�m[�s�p �{ߡwE{�o�T�7-������gW'�
���݇�m��f�dCkiM���J�]�_c�~RFX�r�F۟�3^��+���N��ذ�	C�k�5g�ڜ�?�f�0X�Uޔ�U�t�m =�j��	�.r%�C��z�?q�#.O��ia9�N�8�Q���oh4���4�PF)��0�w2Q�۷o�A! @��l�"1e9�Be�	����I�@F!+wC�P���eM	��4��vI��K	M�"[���>Bۃ���ѭ�N�-a��\Ђܪ��<���fh;�-�#-�x��#��'���;�Ar��M��lR�Iv��I_$s���P����:}.ʹ�����Y�o/���?�k ��4�?�����/Y{eP�%�Lk[��_zޢ�Ь�	����>�����/|�ܻ��wI��n#Dw�O@�߸q�������-%��zi���l�L+��(?Mt�C=D�N��}�3M�	�(�vJ�޽�9�r��{��491CW�6���f�J�ۅ�����~� �lyf��{�	��>��g�O.�mr�v\<{!�!���
=��ü����]8w�XK��}��xn�,�H<�k$�t�X�L`�S���_��Ҵ�.�F�u�iTebiQ�v��a�+I�Ɲ�V��7���Ԯ�+�2�=o���(wM�wk��MK�6�O�D�+S3��$S&B����U�+w=j�10 ���
0gYp^�����1/����hϞ�L�> ?�"1��k�>�\k����(�8q�v��E[6o�y�Yl���:�� $O[,���?Ӗ��;���Ё���������!���UK������iP<�ɐs���eE�Rs���I���X.Rc�+D��.���k��onX�Oi� ��q�-�A ��׍(���'�g�7u���=��g!��M�&'��LH?pϺ.vQ��Hq�9G����d,C=��ŵS���ۂ}���޵��"���Ïp��X�B\szj���s������gy�������z橧�_�:xp?��|a��:99��� ��fyvi��^9/�Βh�=�����|��ݳ���L:I����D!��"��.�gz��)������W�l�P<e2Q��>���[�P[G'M��μx˱x`�e"-������:]���)zT��E�x��0U�С����Qo����=?;���NqjM�S�x�~X��-�MsZc�yneY�E����'{�����`7������4(^��E[f(3�ZS�n��W$���N�Y ��fL�c�`FD�Ѳ���M�/��Ǹ��ǈ���VqO]J�渑b����1$��X+��vyx�[l�7�Imr�X������4��|j��D��0�	s}'��9���]R��,;VM��Huӣc�ֵk�x��8�Y����3r���ٹ L �%6[v�А�H�fzD޻B��WQ��K�L'w
���LضlwXeo�T#���-6#�b���tq_��MnbS)�`߾�|o�6nqc�f�>f�d�
�ox|�Րe�N Y�2xe�$���s�,�,�����!�e�v-pd<��h���-�{`?uu��4=N�!����"��g���N�
a�d��tғO>N�?:NC��8� 4M3.������[o��訫ݩ���$_���٩)�L}�aڴy@;I�{�.-�<���!~&0Co�����Lw��N/~�Y:q�C��x��_P��D�
�`���B���9�lvv�X2�[,.�������˂$�M��p�N�>A�])���={wqF�ǆ;��i�Fv1mݲ���9���,����gY���e�6n����t�����cpVE��/NLW,Š)�01�����Bp���y� ��׎e��f,�^!����d��%@�����B�����3B:��r>��\�G�-]Jdz���*L��n �}��3h�$�:��w���0R�=�M���Wc�KBk��J6G�Μ��Ӷ-[)-�DL��UZ:L�< � 	�d�5�c^1ȯw]���hW�7���fp���d021��[e>S��J,�Mcj��-N�TL���u�rZ�d&���K�n sNb��5x�8��f�%_���Vڹc7��k���=�|
�j�؏k �Y�`���CH���W�	�<��֤���<IA�H�þr'����߹��������$�g���ĵ��=�s����A�{{؄ͳ�DC���ifjZ�G<�݆c'��*4���6AV���*�a����Ɵ��SN�35=!C���b`�nd�۷�߷�z:;��)�����@\���XkG�QL<��� �m����z:}f\��E�����[Yx$#���l�&t�}|nn�>:q��?~��7�T�H����7�ᨍ	��,,�/𬁱��ط��_����"�;ڰЖԜ��ک�-#�L�?�z:�g]Ů��͘�}#�u43,�"��C:#�%�;<h���������	S�\~�V�>vbO��TI�ϼ�<r�X&���}||7z�����_��7v���SY;�y݃���^+����75nk���q�0m%M�i�^���F�:���3�A�K\��_:|��lVV�Aÿ
?���8�w씹+�ϊ�;\-X�q�s��I!8�)<��@�T�#��}�z�����_�@�e��6�Hw�?Mv��*��6�S���(_r7X��?�G/t?����W��A�����hthwʗ�3�AԯI�e +�|s�xf~�������7l�j��;;�d����J��؆��yW�Ҳ8��ZRI������嗩S������3�iK:�s~�G鷵���q�R�_r� d���Ӷlns��9#)�}����4/�3s�ʻ}���������0�	:e�q���ꐍ�(����Zf,�m�}<@&�gR�s(�t��e:�чt�����M�{h���~�.]$#^��~���xfxN�p����E;���	q��7o�(]c��.��x�~n��+���r�_`�HH���<�[a2��w^aK�Z��p���d��T�n�Ӿx�h�2����北������wx���o���vᕧ�׮]���q�m���9荺.���7�W�D3�ikwk�С�;��Wc�C-�VSּ��~;����
bP=��L{��k�˭b:�~sɝ@&�r�|��P��/�f������T���(x��>9'7"�M0�*9���&�ǐs�k��V(H3�$H�XH��9��!smCsb3�x��P\���utu�U�¾�)���3A����,��u]e���g�'wu2�\K�bv��fg\BE \�L9��$r��A�����/cY�#G��ޣ͛7r� ��u1��9�����@���,֞q,ҰB�C84�B랙]䅀�$�T���0Y���RfwnL�+,0]��0�9��P�����;����S��l6G}�K�pһb?�/�f����H&� ً��X�ei���4x��Z��Oс�{�s��2��y�!�7� �x�u:ᜨk�ӽB�1ۉw�'�iXxR��k�}O�8�A��2�9�]b8�,W�Sg*��ǎ����U��� Up��qq&��7�Y{:x������!r���su]N�+H�v��~Կ���G�>Ow��ƺ����{��%�,LW�j��J�&�;��N���N���ξ��Ƌ�\��`"Ӏ&�h������R�m��=83��Nv���i۞�>L|��	:�W�u�<h6$��V�ۖ)>�]UNM�Q/�O�7d�8�%
�LB�DР<��f��g���2���0  ��7�Q�������{�~�p�M��+kUcv ��I"���=iAho�`��>55K��޷�?�	�y�n��ב���*W��y��� <ᚘw��U'Z_���b�p"��Ņ)���9�3�!Ǽ�^Rh�r���tX�C�X|�sX2��օ�x�?���S�S�5�N!@A�˭��]MW\�g��8h�\�_�E��~�M�8p�m���ޞx�0�1�Z���'�]�JgN��\v���8HS|�[Z���8�Q}_�ͥE~x/�}B	&���y~a�ɼ��o����7��@�DH3{����o�A�r�ԇ����^�=���]�}r����R*�������G9������Zu�ƍ;Řq�1;�?��Z�)�%���R���ոi�uB�k��^��N��F�LN�X-	ӑJܯ��aP�YZ�i�]3:L�f�t��Hp��N��>�&t��sn1��K��M>�"ʖIlp�"�O����#���ZvL�12�II��$���Ay�D�R����UM�z���h�� ~p�ɷ�LmH�9�H�GbP�$ #�HF��7�n�3�
�'$���[K8�k��8��������j�,@��5Y��CցWiK%�ͧ&�y� ڙ�o$n���`2d
�0x�-/��Z��9�m�Nھs� ��(k�')�B����_��i��6t��X�#��uzn���eV!��h[�������]p��q��÷_��s�(�4�$!x`.z҉�@�c�2��8u��w�yQ����G�xZ�oyN���A �l��V����-<Q�3��p�LgZ�U��^fiya�	}hh�#��,u&[� ���-r�Z�W�M��(Ci�ᬶg��(��r_�9�@�z⽃F����m~~�ޡ�!���B�z�j�~�ϋ�}\)dT�,���w��HӻƝ�Z't�����)щ"n�|�Q��?�	T	N�)#�a
ǋ�]Z�6�� ��Q|��F2�+K�|`D�c�,���N90ë%[�O�`��>����UEK�t�z�[E�׆�D�s4���/9H����I��c�<�&�m�%NNu���Ƿ�B@^��Ξ�U�@>(���g>��B��6��<@��9�&y,���!�%+Aq��0��/�����eA�*�4�����r�7`��r���a5��~�gd>�_�)o�#�ѦhK�waV�1֭Gt7�A�`f�ќ�I�}�&&iC� [8��K_��o��M[idd�5�B>���T�BC�t��ѫ,x� �ےx�8������e~�)��>zXִ�������z�������w���ׯ�ǟ8�ˡb!���\�NԻU��qld���G�֎v�-�W���~Ϟ:-�e��T>A�H8411E�`��R����x��5w�>W�Lpp��ϴ]�x���N���+k�LZZA���b��͘3�}%Z�j�ac�A���v�r�~[|�WVr*�\ZZ�?99�S0Lw	���6��x�P̵C���V����P��j����� �:�c�����Ļ^2U���lәi��bp�W+	y`�P��5�kW�/�*S����0���\�9�c$۠�CC�h���+q4{�~�Y������L`�D66�Y],��i!����'X[<{�<}��9A<�G�5�{�GF��m��7�u�e��PÙL�f�t|��0@�{��G�^�o��1M�ח>�"ku�Q�A�\�y��� )h]�׮3)a�1"�+2�!�����>��g�L���#�§l�x~�̬V�!6����\��g�T�Mh��D��O��.	���\����'�`������.k]d<��4��ǋ� '9��=(���x�qgj�EF��G?dA����Ǣ�b��p]~�0��&���=�6�Ѓ>�/H!M=Ļo�M���o����#,H Q�?,#>x?-.e�v�}0ca�S'��J��fo�%d�S���/��=���������<O۶�7��/YN&3��t�l:O�{,��z�ޣ����pB��x�����[�������Z(H� ����/���y����{�>ڸi��4�K��ܹs�����V�&��/�k�#� �W����(�'VW�|�X��y�M�������� �<��wc�Mv��P�A�sI���#s,�)u��{�ҥK��<OkB�j��^y9����;;>1�B)#d��f�w�Y�(f:�T�CZŜ�wg,t<��*��͗BV���d��	ݦ��~��-l:T��F|q�����8�"��rկrY�/�p�t��$hnz�#�1ʌi)����V��z�J�V�JE ��u�	PL��碰S��W���B�{�駙d h�����GK�B�f_C0ߩHu�Y��rDemlLh� �g��9�*��/��O����vL��M��T�ݖK�b����@.�sJ�9�nH��$�H~�m9��0��@��L���8|�0�qU����	�G��5X��F[|��1�S^��C����;2l�I�$�*a���n���/�h|t��9>��ll��Lt0CH�z�6�f�fT��'�WO��B��K� ��Ewv���]�h׮t��-
��t����E���o�ҹ�ප�������̳����1�K�Z��{��w`?�H~rݺ�n������q/s�s��OR���<,�6���'�[@�;l�|��ǪV��c�@0K$bBH{�ܥs-v�5��'?غ����Yl�X���YP���MKb-wE%\k�wk��I��1�r�dח���4#U�M�j��7<`�;-N��]��d��ȫQ�y)PiN8��	�S�UUv9E�*�NY���{=^�-��kk;�Y%�Li�la�T�I'�e���'"�U���b0W��z؎9�X�ap�b8T�ul�5�E=��uL���J �f �z�>��8`������CCC�+�����%�%��18��؆z �>���}���Y��u��4h��T�ɉ1��wD��%�:q�u月}U��a.,,	��t�����>X�m�"�!x����qoHP�i��T����,_v���O����R6,�9�	˓��e�~�7���~g��hIh������x�qg�^�`���#�+���:4#��������u�p��gx�zX��O�Ȼ�=�{8=-[o ޑ�Ӱ�T{�~�F�̨��Y�:8�_9�?}��׬�}pp��?����V����a�5ğȱD�w张��g����zq�;�5M�W���g��n���s�nx����(TB7뙓�T�����1̒�b[wkVj S��q<^�`����R� ��d��/5oe\��Y���+ѭ8����$aG����񁘡�Ia����ꫯr�2��~�����,*�7�x����K�X���K%����cp;H��W^a�䨲ߩ硖�<s������z���������@��:��ˤ>���D1�"��s8q�8+g�@ ��0n<L�0"��z�-hiQ��7��ߴe3#��;)|��9^�g���Z��x^ _%$�>	�A�'N��{�@�Ǆ3�c�v��a�I���+�z�hs�l�՘c���W��@�rq�N*���}�7��5m�
ֆd:A�3�l�W�xg=|�����8uP�+x7��X����/��x�x��A�Ӵ� ��˿������/�`����>8��н��!d\]�����X��	�aXH�j+	�v�[�H:d�&o$���o���s��k9c�6&�$*9a���fĮr'(��i�KE�+"�F�cP� <�	��U�"�x��9��rQ�
�����i�d�Jpq7�	�  �Jk�ju2�Ff��1(����&�|}ED���)����0�iph?�V�T��1(��u��.� ū�9&r�����7Ed'����YANǎ�ө�z�+��1�)�4\a��Tr֦E���`��s���{N>�J�@�� c�-���"֞?�eQ�Sm��@ �S.!ՏY�q4a���&��g�oGYZ:�ϑt����M�7si����6�r�,.�>���P-&3�A�Qi���$�����Jun��,ʏ��bx���y9�\�+�X� ��PK��K����������7֚?�g?���/�A:��)���,��-�̿����&�;�5O�20Cj�>�jPxN�P�ͧ`5~#���5Ȥy�I~�4�������|<�>��p�:(]�WM��`�����I��"V�:��r����%tu]����^J�  ��C��7q�W�r���B����SV��ߺ����
N��:T=AR{�d�Se)��j;E� !�Oms��ν��9�=��o5%�b��*�O��[�C%n��=R���z�4
�ݛ���D������E��g㮸�n��/b����0�����}[�exU~7��]�b��ے�5���C�t��{�p��y�n�e���5���db�l�k~�o�S1ss�,p�\{�2#��]B���?<���w�޽@k o���֣����S�ē�=N�?�2��S���U��c�wx�=nD��'�5O�&����~��8/٭ƤE�2e��S�
Xʲ����ʴ�%�YT� �Ō9��^������� �ш}���f4En"u�����N21e�Ur�����c�*ܦ$Fiz�Y�*�Œ�H�%��`���A�*��Wv������6��;���NA���X��ɡh񌂢��)횯E2˙�>�k@i�JsW	j�}F{�Tp�f���Ш���$'��q�#�"E/��b��{-��`>��#AQ"�Md���9���*R%Ͽr�p;����e�jw���1k�5V�3��B��/�t��v򖓜)aK�x��0�N6C̥g-��{�y�e88#���C��;kp_u���aة?[�s�~�&�7:�*��y&* �q�+2����
�}``eW��n88=3����x/}���om�rp�� ^��-gΜ���{�'I�+O�ED^uvU���o�q5�8H� �rH�3+�C�][���A��H2�d���hH�F��� �����]�u�!�����#*2����*��`3+3##<<��]��{������xO��W;�Q�J��jz�l���(�c��"o����c��ּ@7�y���q,���D��O�؂�t#bn��!��F���!4����-i�b���OAcNhy�x侅�B��["1�̵�������jk~������)�[D��s�**]-mW��)b��ؾ����|��~�z�zN�H���Ӿ���?��JmA-ͫ�Q���u	��1���������mL��e)б��Q��	���݁��\!�z�s%��k�=����-Qa�N�랫���{6��(��z)8._*[Wz�~�+@�tHg^��E�V(��F,��:^X����c|�ZF���n���_�p�d(�@yEQ$p���Ά###G����g����w�}�>|��'�+n���_~��믿�?���枷�X�
'��=�1������g�~��y3h��u����f1)��׍H&��Pg�w~?N����;�[���R�cB�u��16�����ؽ�i;���J�@"C�k\Y�1r�s_�������W��"��6} ��G�|e�i�Qɩ�q�w���x�:ҥ@���x�X�M[H�P]�b�-|J�)XǡJs�d���5Н��f����B�Uh��)\����k)7�A�k��"��B��A�˖k�6Ϋ��X9�s.aIb,���o�O�˯&]'K����]�	P<�/\5���Ց�%��c��ر�a� ���sXϩ`F �|%�c\�9m.�`�|8$���=/?{!b��)��	a%(�e	�"q��/��]:�t/H�`���ੂ"��2k��w Y���{`fv��{����>����'#�����a?���Ϳ���������ٹ�G�~357�@�_�/����>3o@�֍SϘ��|:>�&c��*{M\^U�ğn[��X�4~�k���D+odcB^
�^�;�n�~l�mz㳔�{��b20�9>w�
Gf�)�O�� ��^A�W?���r4�hxh�8��#%�{ѽ��[�3(P�V���[Q|��t��a�o��ǩ�8��c�)��c���e\���>���V�n�{�^�tк����H�?�6Ah�c1J����w��l�|������������m'���נ/�}���}���<�����}�tw��c��O>��-s5|���CVh_�Ƅ�!���+ok^�(���+�1��U�w��Z���:�R
���&��1�$�����X�����b�(����^z��K$W�l��%_u±	���fZƅ'�U��wp�C	P�<�ƕg͑�X���=�����}�请 /�����R(V����r��~�x�,�\��3܊��gt�>���~�wƆלg���	�����Y�/��4�%�B��@�O��J��t�����J%3��[��_�?;s�ɱ�S�}���oߦ�7�<w�7����EZ�:�ٱ/����8u����o2���(�H;E��2�i�F{?���ߚ(��|�~&�<�z��Ukk^��T[ˬN_����_�v?���]t�j�h>
W]MJ�r������qL�]ufg�� 
r���"� *U�����% �6�F��}���p@�Z8�5
�)b���{�����jX���~׾�b���~1�J��n�EsJ��E!�j�3s���w.W��λԝ�M�
=�X�{�8���kx�ԋfs���;��f/�{va��/\���/�湉щ㓓�3۶U惠���:i,�`�+#g/]���W�����o�;�Cq���E�P�!��w ���z�|/�6�b�������@_������m3?��
8�n���Z[������L���9���ҜL�[Ȩ��v����ګ����*dW,x�>� �<?�yhؚ���ZPl>��1�|����}}ܚ_��=o��]�x�>��cφѝ=��s5�*-W�R����q-Xe�(�e�˓����w�0RO�J=/4pe�(���{���ekD�1��jX�!���g��^o2��ƍ����V��r�ya����X?l���ժ_��m8^:�����c##CӥZu�:Tm����A'���/lx��Oom,�_ػ���qqa[}�a�����7� �Դ�t��YΨ��D;
�d����&l�D<��ܔ76=F��3�/�]��ּ@O�+B�pu��u�9�.� KY����W�޷��6�RHG��A���|Cf�r�\�XT`Eg2���R��"�]�2�r�m45������+J��Hv�Z�̿x�h�
��" 
~��g��$�Z[�����+^�յ�n~!�
��f+uI1��
�=�� �W��
��%�ε��V�$�/��{�W[*�Ӗ����}����e�A`"ek��yM������I���pm��#�r�izz�a�U7F�B�R������mְY�q`�s�( C�vs��h�k������Vhxt���g���V��@�C��ҨA��L� Q��*'�W�T��0	օ�*�5/��$d��(�^m�˽��1���%��Ǩ���T͢�sp/=��c?�"GLd-p���(N�#4�L��[�;�p(v,>�� ����׵c�׃u���\k����"�J�q��'űF
r 9�����}]M�V�/yem��-.,�?
L�\����4�;�}Q�ܾg \���)O�=C�PO����Yx��=�݊/<�������[�Z\ 0c�w�KnΪ@�z���:ȇ攘G~ΈEr"�B��P�7lf�*����ŲMQex�p#���:
��4G�>���'�p���a��f�f����,s-�U���
�X�K�~�!;n����M�S��V[�=�]-�"��~�^C��.:�߄U�����F�/���t��GX�#�l5�R(SQtB�d,J�Q��->�{�����-ss��F�u��,s����O96	�Z �H[4eK��,�n9��g�%(�Ů����km��D���
y�跄����H����B&~	G�-�5��V��Jp�J�
�� ���oͮ�}~�t��
��e�[���ECZ[��q�j��㙙i�(�&ȉI!���G�ƀ#���뇲_��YQ�� �3��H�.^�1��,��9�r��c�}N�|���r�#�	u�[^C�º�}5ښ�1W	��
��B�b^� ��	ؕ��?���[�v/e*K~Oٚ�h[�޷�m%�~rLݸ���z�~��c;���ǎӳ�}�>|���F�u����6Z���0���<r�9�Yԕ��$`T+C��Y�J!ǻ�vz�޽��20�
@�Zc�����+R��u�v�㍢�Q��p1^b0�����3�a�-���~>���C��矣��p���9�j�.� m�l��%�k�s�5��ynq�~ b�k��,�A[/A�;�n���(uCa�Cy��j5���
/��IP�7J>���A�*H�1t߱�'{]w�%�NVH���=�.=�����b������Yan��f��?"�Ct��}�	���p�π�q||�3b��k3b���%s�rEjգn9��\C��a�@K#>����+��<{1��~�BKJ$�r�K���)�e��D�"{$�g�֩�.��D o>m5;�}�ښ���(+q����s5k�.,*��&��[������\vդ�E+�А䦣��F	�p�J�=o�]e�W�Z��"�eÉ�[�M��r�ER����ctA)sJ �Ŗ���W��=�~a�~�YKC��[�˙_��#r�E$��]F�2D�x	'�/�rʋ^�Iz`�#&�.�d�!��W���|�w�����u���'^��^n���N�R5�i:�*E,��b�xw�;c �nxX��"�+4:<���� �tW.�ԑ���[Xl8�>�k5�"�醳�.��eY:T�N�`�py͑�$J0��_�о]���U��H�y����lV���H�J��lڴ��~H�?�<��!l}^p4�� �~�w2�.5,Z���[��%���4���M��6�ϱ�q>��� %,��b�.J�d����K^n��F��s�^�p�����I?S�3��8�w��I�ެ��@Ϭ(�\�����X��R�-]K��* 9ϋ����ϋp�}�|���i������0�^�~�׾�+�����Ҙ�'!
XzL�}F$�y�4 f��]j�;4{e�	ֲ���󪻼k��`>p!�n�Q�
 WZ���O�=#�,e�L��U�0�%K��gU����} ��u}5��@�su�tϻe�u��e��yl���D�7,�	��Ѝ�z��g9�ֶ�^��[o��y���d!Z�����W_�:��:����w��C�[�hq}���o(Yʁ.��K�J,���o����m?,às���.��l�hy�<"E ��p �s��+�C�Z��lv�oc� I��|�� l�8*r��+��n�[	�~������<1E���\	�����^��-���*�E�C��?��:�
� V|�4F���=���m������Ba�>��=p1�#�߀l Jϥ�2~�����9.3�aeb�J�k Уvr���f�U5՜���ȇ������_��&_����1mu�KL��kkϞ=,́l���j�������$-j�M`rr���>�Yg��XrN�n�7hnV*5��K]�>0�ר]�{4/��6T�.��~�+r��Y����k��b���՚�Gؘ|��0�}l���azm�	��Uq�y�
������t5�
�"Z+�i��U��D���vZVT��z����+�{){������9��1�L4Z����>I	jb�S��o7;iY�� �z6TV��<%��4�O=+�����H�����Ps�ܺu�Jm��RtJ���}��%�|�p��DiG LO�>��V�� .t�׿���ӷ��m��+�}~n��|�uz�w�0����ohh��� �R�5�D��E��6�f��AiYl��ە�ŋ�rܠ�u��9�X��h�/�~y�����0���;V��"zC+|EXbi���������.��
�$XB"�<_��!�����c�A�/�y|p��;�YF�c���nКױ�7�?_�1�����gM"TH�2�Z��P�V���H�#K
e�%,���8�T�K׺�d���=(E��}�V��J<��u��j�5/�M�A�B��z�%�Ox]~�O�..䮭�͟Y���������v�����o�[����&�#Ko��`�#�1b5a/��o�� x x���q�+5���\|��o�˵��~����7�~�$���Z��kZa�wl�_�RK&���UK:��Sņ3!�M�
O�/�-��&
X�W�0�]����{R.{6U��y�W����[�>�Oz���`e���h��v�N��B�h����λ ���>���������>/���6l�Ϋ�� ͸�h�Ԫ�,w:Z�(�q<�<p��0��;k@JS��7.�kA�VyjI���	��{+-���"�O�/X��W��y�n4LW=����V�zYjy+�\cQa.v�Z8@�V�=��C?����]���2��Hffz�$�5�o�q#���P�Q���q�f�Egϝ��6�"UDK�j_T���{L������^�����M7���]ܻ���:��K�څW�@������ޫ߿D���rMj���s�:q���Ӿ�bUY��W�v^�Ð��}̿c��$pnWɼ��+>H��;��Yk��(3~��'�2����EqN��g��׆�^ξ��]��/��珿��C�oa�	��=oBjh�C.:39���d=9�l�=���h�R�w�yH�ܸ]-�aк�ϙ��I�.�W��y�n�y�L�8?Y��l9@�"+�?�_�Y�gz���	}%�hK|߾}��C1B�:#��@ÿ��+4}�
��Zcmh7�|39r��#UC�g h�����L���kc��o����~fa��Q�7���r�n�&8������o�ǚ��c�^�E���7G���J��aK��-W+"�BA���dHSpi�@N1ׯ��=��;P�e�]�Ԭ�T��E�,��u�4RO�"_E���+��uy�Қ�hS�7�}�O�p�ss]>>�r,ͪJ�K�,�*����Wj`�<�޸���cI�u�g�R��c-�.,~�Da�U�P��2�[��0N��[��� �ւ��,�-ϓ�����T,����3���2�����&Hb�ad�i�¶V�y_o�W)U��!�S��H�4t�g,sB�#�)gBm��g���Ņ,�/"����))�J���s�Z�z����z%l���u�]��Em���V=^a��o��5�Hx��!�� 
ǃ��w�u�Q���7=H)>��S����9 ��{	(���c�+�ߞ` ���ϋܣE��g�,�$��a� ����馛h߁�T&�as�`D�/6D��x�� �*<z������$�������Kbu�7a��7��x�:�&�%�lڡn�P p�n"(yP� �,תF1h��Ȩ�y��ȑ��	K��0s��0�İ2`���X�,�ϳrA�� 􅜈��������Z�|��<�J�eӏj��r��.�Ө�.4mמÜW�W:?{ͳ���|0�/.x�5R�����|�'&���p�9�����r[/o��+~M~N{r�\��mEm��8cۮ64s���^n9� )��+����,@03!��4X�`���/~��Y6ZXia��-mHQ{�����f��A	�R��ʈ��'���]�\�8�s���-��3��N��$�l��U	������=
�޷�*�!�	L��/;Z����6�RX�L[�T�Fj�u\�1x~d�
gg猐�i��XP?�i|Y�3�P(87��;����o�;�}W���<iwb�Ԇ��>�\����8��M��4�B���i���(,� �p����.��  b@��+���?�K/��(4\r����Ņ��sa G󙺇�I�R0�X��ye��vci}���myr���'��A�C�B=�n���Ӑ^�����������ܥ�@����Ujk^�Ǒ%1\�+}%ଢ��s��}�����X֯��;:6�eT�~�i:z�(o̒�&�s�� �3��Gٲ���ԯ�AX���H����S8
Ҋ��{�A�z�sz.E�(Kv'�"��+��O~B�F�e�J&�����4�.��珉��H�[�e���]����1��:F�RO �B(?�������6�k��hZn}���{�^��x��-�hՅ�x�$`8s��N��ݭH�:�g$�!r"��ةz}����+sA�[��V�T}q��(���u�`#�2�Ȝ��8�x���(M]*#׹m������?J!��l�A��zZ��	+�[�����-�%+2��A�;w�?�AQK�O���c��V�zY�r]Z2�2H�}�ښ襤d�nV����_����u\�s5�%��r���d� ؆GF��
�"�1�5�a�C���γ���n�b.ö����ƫ�j��v�����
���J���{����+��.W��>c@���?x.���	�8',�j���N@�C��ݬ��=2J�a���"��X����l�2�y㡛��h,^3��9��8p��h�x�r�'��P n4�m޲���r����q�'��c�}��i�c숆80���h!<�KԪ7��np���''7Ҿ�h¼�I��{4?���s�?��#��R��G7�`i��/hzͭ����Z��^���A1xiE��/���-�س}P&���w�/Y����
�Ռ�J���kk^���yP�J&R�K���F��A� �I���ք{�c�6��8,/Nc�������3*~tTܬ@���mNk�0�2;�=��۔��h�ſ�E7hq�������8�,&MՁЁ Ra���&��Fp5���ǟ�s�<K3�Wh���m���Q�U˕(��<i�^��N�]�j�ivz�u�.]���N���s�n�$Ei3W�0.
�K���磞���>�q|v������3g��瞥�>8J7l�̡Xa Eb@�����w���D���d���Z0}�gno(�6B�s�O>�}������Bo��U8��_.Wl�Dbc�!�3��d^��
^��.�����z5������&�r_� KȢ_����RTk��>�+��Ӓ�|��v�m�tƐz@���`���j\v���j�Y@o�\�4	\�LǱX��L#�#�u�vz�l�`��K�3W.2��۴�9zv�*LK�s�o,G���:���ϳ��'a hu�P���0�X�@��\����y�~��3�z�����<J5#�kH8����j�댜G�p�E(d�-yQ�ֶ�P}b�#�֗.����}��͆�T�����#�g*�@qZ�j�Q  X�3�|h1b^R�$4�����^y�^x�y�����o<�1|	͔ؓ��+J���:�<�f��G099�׀�1?7KG͹�7
��w�K�&�k��շ����#�r.Fꯓ~ϯF����v>j� ��+h
	��Z&�����~�� �"��u�!�x��aX�pr��9����8~�.�W��}�������H�U��X�~�K��IZ�wf����`�k*6\��'�&��G�'�|�]����������/�+fC�tq�	l"jR�d,�N�~�9c��H���T�����*ca�5��
Ǥ�xR|���Xe΃ �+��ȅ��(�A�� ����	ڻw/�<y�>��S��@�a�`ec|/ٚ��'�Y��]���C.Q׸a�V#$K�%�����ô��j]c�W��D?�u��+�Ȃ�*)���q��=?�����O��_|��}�w��[�Ӟ}{�6T�ӧ/��]2J�6;s���^��g.0���MC1�w����q�Go��.�ŧ�~L��~�������:�>K�#� x�ɬm���SNճ�(i���z�A��W��{}/Or�½��Ⱦ�u���g��n�v�䫼G���u���:�'�ּ@CT��c�A��VJ�#�:�βΣ���^q��.1
6���!�J�J��l����Ty�|��64\��n:H<pm�0�1L��u
a!�����L1@J��+Ua4K�TX�dܘ�.�����X���e� H���VS�-E���1NR��t(����}�Q�c��D��N=0�mj�0�ju��?F�����X���)�j��1cz��I���f��6R3B��+��}�%@�@��}��bA�xP�A	���,���x�C�` ���[�2<B�/\2B�I�##Rh�7�0�ܯ�c]�	�)le י' q���j�H�J��:w���Y3ob�����޻����۽���ry�� (+PBP}o|l#��#:q�$5��{.1b~n�E��8��NP;�����{ &<ǀH!�Y4��� ��t�+آ?���$C#�R�Z�V���"��ru�y���{-���p���� ��^rE}`k���^��p獝U/k���k>K�(.�k��������e�"$�<�϶Gl0	ؚ+��mk~�8�}�J1��*nѫ�m?�킌(�0X�&\�|��'m4�Z�2i6��~��rMcM1?t���t�tJ�4fʽ�=>'w�T���A����)	TJZ��q�7<��fQ�X�@,��#Ǳ �·cI:�}�\����qe(}bշ�r�p�_�eA���2H.!	�![��� "��_��~��Oӱ'i��S�k�f��7@��ܯXo��&{a"��]�>�t��Ė[]</���ቜbx^�����ԙ�������<��Ξ?Gw��(ц�1ڼy3\̕ru�zx�N|~�����ã��ٳg	�7�R�.Μ�1k�%��չ�e�8��l����
4o��s+�P^��\$���u/b�z��|�E���'.�Q)j��[�S�f^A���E����=�wV�]���z[���z��YD���|u�ɼ_Br���~*5�ֹf�i��FX�����.^4�_z�~��0�.�$Nh�C�1xy���R4�y��ω�h�;�틗�������m��W�-'����o�踹����0����������E 7��,�*��־�����6�w�N;vns���G�,f�2���K?��?���!z��?���R���"�!�2�K��V���.�Gb����Q8l�晃n������ҥ�ݷ�q K�y���}�b2��* ��6�(�Hnۺ�v�Ȏ���<wΝ?�1x�è$it]����[��I~/��G�{$��+����爼�����j�b��}e����b�Z��WT�ͯ�k�����ƫ���r}Η]Xo_a[�=)��Q��_��-��^�wI��r������]���p	�#G�����E�uX麹�&��`T�]�,�Ӓ+�zaV�������Ac�Ks�E����z��/�tw��=�]��U8b�f�ʣ�d�V�q��"���v!�Q'`5ĕa���k5[�|������~���t�=��2u��y���9m�u��g`��1x�bou$L`�$����Jɡ��g9�q^tu�"VE)���}���'��7���v�R��� �ZԷ���Fi�N�c#��g��(������{"�^�B	+U8R�EB: �A-��@]k]�1��V�>#���K_�T ��ͯEPt�A
A�p�*��Y��O���:�1/�\��oE���5��W��rg�h�ψz�6 �m�t䡋�g�õ��9GO��R<:0�|&��K��B�H�@Jz���@�Wx��b�&��#�݀��jw���+����sU��-�1������_�9�	I,�Xp��w����ZGS�Km��IU�T0X��PݖB�ډ#H##���wǂY���-���� �nfFױP3��m����˕�jQ��:!%3 � l�޷� ������)8H��-��֟�.wCPl�r�������Z��m�63a��t��e�f�4���kuZT+	W<B
�_&�~o����Y3��̕�F)8ESǹ�CX��	K�@�ま�����36�T����
�@���UX2��9����~�y�y��y/P����{Y����>��wʶ�\���ů����z��^��}5B��t��d��1N�H��0\cdmi "m�����ܯ���Ra>���F80K�+2���������/��L����=�x`���<1��@�i��]�A��EE���X�G�-w>^�}�S&�8:��lN�+ ��o���ǧp#U@_�V�Z�ʇn+�a@�\X�����Hk�{�a�r5:�[y(J�j���p��\�V�>$9��Wpx��Y�C(��3o���\
@�Y7?�ny[�9�2&���s��b�/��������)mݺ���svDy�xl�)�\�%)��ah4X��ɩFI�J�{����GQ}A���b4[m�ք��V��FI�L������e.�%�U�Y>�ܯ�K�Wܼ���?�^�ͻ�gx&�����'�u=�-s�o�����C~[��t�~���R�y��.�!�޾��z�'F����"ɹ"m��8�������~����ʐ͏fH\��G`Mڶ�?唱L�!�rU�R  =u���o��{�#�!^r�#�t��. ��Py���A��ռt�-���_�nC���ƭ;�V"�j����C���X�UHR��}�k�k}��}LЂ�MP�F�J�v�.rѵ�7��~��=���i�,����,�����aaX2Br�i�$q���N�m�;p��|}�F�Fu�8() �A�����*�{��wxm&F'y�u���a���"	�`�LN�a>��grr��������ݶ����!s� �@�c�-J�>EEe�z^���Ak��0�����~+r__k�g���:Ot�O@+Nc�i��ZR�x�������-�.{�]�ۗ�ּ@O��֖�e�_��/0��� ��-��,��p��ь���NR@\�ظK��E��ֶ��S�|LE�5��|� s�K?�&��q(�����D�����,s}�8��ŝ4Ϯ��~LR=z��R��� ����
�y\�Á�-��6����,�st�	�BU��z�� ?�W]������U0|�͆���!ER��Ǳ`u������'��E�Q�o��m4:2*�����Ӵ�-� �i�s��8��*Ր�gΞ�:�CC�\�c4<6N�F�)GL}�i�@/q�Y�k�����=*W
��ծ�^J���o��J���1�M��w?���6/��.yŖ�w��R�}w��A��Y�(w��6�?���:���D� ��p����h�\�l�a��EX��l��z3a�е��nҵ@��
��bChv��brh;(D\lB���\e�)U�H,w
<HP�|N��cJy�C�բ"��	J�&�涖���zS����@=��w,�*Ȣ�}�Q�bׂ6���zZ'��^���K�/r��w��{��޴i3��1�\ִ�fw�B��4��]��ǂ���hñ�f���qk�ކ�ָ�he�-��v��ʑ���*mܸٜGʽ��Q�0��_��M�&8lwʴ{�.��y�8p��������M2w�t,.ԩn�7�k7m��gsyFpPf�pH�2ەx>��ȴ��H��D�$��fe�,�B��bB\������"+;�}Aѳ�c9����{���b��V���6�7�1�!�+���ޱ�JR��ƪ����s'X<^��ye��8�Ȅ�5�2%FA�_Ά������@�_��¡5ӊ��Fe�g�Ū݃ϝ��Yr�]����u��M'� $^sf�+�j,��Ek3bV~�<$�U7�|T��G��2�9-���ZU�	#|ڭ��;:g�*���o����B7o	���w���t+�^��am:刲��e�U��4���Ӷm�8�qn��!�6nd48,Mл�����4EMk���C0���F�����A�Xp>���͚��>���s�����6N0=����{���<���m�R-��Uo,ҧ�~±Z � Ȃ+�^	��g�̅���ŏ,Q`������=7V�E��������}�mPs��?�>o��-�~��=�Bp9��k�>�$/���%~�7z�fX�JJ/�{Q�������iI�:�d$�b2��=����F���*���@�}(��5і,"�;�ٶxQj1v�W�l=�p�T���\j��jY��MY���q<�6C�p}� JP:�lp��vV*5#l�i�t$Vw�k�-�bz5+Q��+�K��M�%-�Z�n��+�x����{��Z� W.1C�Ʃ)�仺M*M��Q��6���p(�R���䒟×�1��  �F��RG?���G���Up��1���M�ھ2}���Pg*Xu�a�7�m�:���*lbm
v@c����m����kW�r3�Fd\b쪴�sbv�sC��DVs�ޠ�d����F7����YU3� zý�6x||��Ŝ�]C'j]��t�N��l?9���
�^֯
��\t������{Y�������~�y�Z����N���<:���@^�������_U	�'����{&��SR���R��9�J:�C="�@����5�z�z[��u�K4\�~	��M	�]sT��n����v[\-L�2�ԥAł�2��a1\�t,C�仡�;GjW�*n���>פ�C#c[�B �s�6B�#5j�e=��4�P�������F��.��1���F�+�&�-��c�+��d��Jj(�Z�c���qס��oF.�M0RU�P�En�77�X�ڴ�-���>g�V�zp���^5JR� �!��\h�ر�랕ܶ �ʰz��C�s��ص�X߸�����W��������nyl�����q�߱O?�l�z�+�
�.z����������Q�0�Rٵ�V:�C=�Y��>�о��<��o�5������^�g�t����w����+������?���/l9ђ��*�����+\�=M]��<�׼�8M����D�멄X�k]��F�Zt��M����W�������-<�7 QL�4$#�r46>����[�؈�҃`�"��0aӢ6�w��[�w7l��.�+�s��o;t4*��B?~�84.رwm��d���?w�N�9E�r�]�s��?���\�Ԝ��p�p!X!T�\��iR/���gflc�ڊ���.Y�g6 %��=MLL�^� ��F�ՙ�\�����/,FX�[?}��\l}G����{�@DϦ̘�������hr�ԛ���9���-8�r�1�
��J�8>�A �6Y��~��9���x%����Ξf��7l��a�fC@w#c�.���Ho�6ߟ;{��><\�T���N��/N��1�
�O�<2}�8��*$�RȔ��toq*�cJ��!�N�������ϲ-ra�[?���|�\��;�?_X��q�*V�6��7�B�_7���<~Ճ��w^��y�U�z��0�}盲�Q��L��S�*
�.��j_�n���X�&�Uu��.8JD�EZ h�����[j���n��6GeK��v��9�6,Dl�/�'���$cq�������u��U�а��/.�b��ǹ�?X�|�V����RZw�-�i��G����:[6L�����X��O>��~��g齷���2��Uq%+(�H�����x�qU��y�8�Z����0�5���ڹ�)Ro��F�зK\�
c����~��m|���q��������G��@�B\:C3˛X�������������(���i�R��͛�q(r����K�2U�	hп};����Y%��F�GŶ��y�>=m�Z�&��Y��98 ����Hd �w�wTr��ޫ��dp�H��������a�>���k�@�+�Sd�Y�����N׋���V�(�-�^�r�k�� y8$�9�H��-��h��O\"Z�|2^���k�}�m��
�ƙ��d����ſ��`���L��@�P �����4>6�Ѥ����"G������F*#f3�EaK��O�\�4,0�!�"8�9<���r��L����6n�;6��Єo���[[��Vg����yH��F���F�� ��4��J
���Z���%(��d��	���V��?�0NB'�a��ٽ��=��� 6F�5�C���F�[�F���	�c߾���|��sP|�S^Ҏ�R�Q�J}�^
l�Bl]�A�Bw�vs&�^po��]ڳs'�C���A�v�V�idx\�K�y��t���ϯ"�FP���<( �=�VFjC����KS�t����
�Q:����,ʝb�O�&}U�"�-��c�^���G9�3��:6����.��UQ��}A����gx�PCA�!~�I��"�D������Y����&�kLt�P�o\T�� >ے�_�Xo_Y[��2-��^/j��nk�$y�i�I�d+u�AnS����:p� m�4���ec��e�T���@[[�sH9Ψ$iq��JH�66�:W �Z���%#��n��Q��e��"~,)M �I�ߏ�t!<�ie*鯠�[�D����~`ɶ�W{�7)k���߂D�j�+��[TU�<�Ĺ�u�+j�����#�5�	��Ic�B�r�R�ĺ:�p0�k��6W�B)��"���o=��5���~��r���N�
��]dSl4T���ͨ/J.�Ʃ�462����a��̞�6e�2$ᄊQ�Zm��C��@��	{$�(ti��_ٜ�'.��Az��7���L��B���*F~��>���q�~/�؝;	����r/�r�,'���u���Y�~�|�wޚF��^�� QP����c>v-��]�g�U1r�6�b9����M��Nh�SEJ�M�`h������kc���n	�� ��4��SBY*�u��
m�t6�a��X�pq�i]ἁ�+~9JA^���R�Y�粱IW��$KP��h��T5�fj|�-!^����/�󹰁'qK�uZ�qN%Ma�����?��w���2�q�d5c�5[4�Zئ�����.x�`����lm�7��.]����p�H.t)B/�4+56c�87�¼m����m��/�J��y��u�N�!}!tƍ��@��������5�=�8[�$���b�+�q��9O^�$p�f "��0�`q��y���>�1R�z���q��1x�j�ʼ �+..��C&Pz�����q��.��'��)�2�K��u��ss�.�Ѳ`<V��s�-ޣ0/�����C�0J�=j�	����yi؀��̳*Uknd#7BׯJ�T�^!�8��a
�RW{��E��[�EkMB.��.g�JJ&�t�[�"�䣘�(Q�"�d�O�?��
<���^x���ꈄ�n�-t�?�A1sH�Q`.�sQ!����[�<N�.ؽ{7�s�=t��C�rh�s��ʎh�b�v�^ �'���$����W�(��π)|��qܺd��l(`L�f�^�2O�;Eǎ��'Ϙ�s�F���<]���Ð"KJÈ����ڰ���ښ��M[+�g}��ϸ�|����c�_q ��fϠ#>_"�0�����׿�5ǵyÌ�^tAb~xx�Ņ��5�_�s���P��	4�W���J���g���j�=�̾Pe�7�`S� �E�.o%������ڴ��[��� �V��*8�\���c���!�o���"[��j��we��g���5�qap\}��o��^�F�!&�	D�K���7oLR�QG��v(x@�c�q�,����,W/2��ƍZݹ����X�����J���~�q��9�^=j�	M�Zz��s��G�x��ٺ�v������>�����r
h�6�5�֊��Ɓ�v%T#��.��E������-�A��@w�0��(�k1*�����M(��V�"��V�	+!�k����'�qb��5��N:�W�CVA�qǳR�1T�)c�86��+���rn���9��tyf�>?~�^}�mz���iv��q��Q�QI��=���u�|�ښ����$E��zSӲZ?K�_�/��G��A�t�˻�O�R�~����'�HzbѺ)HV��԰��BC�]�~?T0���M}C�@��/jI�w�d�@�5�q�_oׂ�������N���N׹
яf~#�� ���}�y��㣈��E]�o��}��1�^�}�IԢ�R	!Hq_L�b�W�\	j�m��P��m�nֶwo}`3�$����;X��8� ���<+f�Dh�G���	�B?��'���!�����F�q��?ρ��HH$�n��;?�`���.{X��i4����V7ʧ��\b�o�Z�%WYI������С*I�
)=6p]����ֵ���s�g�=F���?oz��9(!4��k,�Ӟ��� �*��-K/�q�$�u�:�o�Q��<jZ�N���9�煬uY���f�P��.�]�%M3a�0�U�b�Z���2ݵq���
�<q����H�z�y<"���i���.�W��y��h��|W�ۢ�G�:�\�-�Z���
�j�X�\}�
t-���I��T�[����S������A�W0�o�Ԯ�s7C�!���[nq�[l:�\�6�W��<?��=[)v4��s����_u]��=s活G�w�uU�ak�l\������� �����c��0�>6���kD�ҧ�B�ٱ%���{����x�9 O� <b�lX&��qN���˙~��EC($<p��<��XW~̖--!�Ksja�����R��__���r�ǚ֥|��Ԙo�s5K����0c��0����qN+��Ԓ/�=�b���Z�1Y�9��XOT̼
��|Ay.Wj|DӺ�
ʄb��o0u1�<����E�լ���4Eo�0gp�Uh�LI<I[�l��[��Rê0!�����;���c�R�S��E��+ɺ0_���zR��ٵ�kU�\�*(�?� W����V��e��dAE���Kr��e�7*�����ڱ�W�0┯����8���6�J �UG<�@��u9^�+�E���N��\��N�_,��ˌ�}�1-u���Z�:/�
vu3�ΌR�xs�B�X��B�^y�4Ɔ�^
uI���U�J���-��&xU�|�D�M7w�`�Z��\��Ї��J�
�(Je5!��9�O~Vj�#$�I���
��Yo��y�&02�U��0T��,E�o P��]d�Vv�z=;���.i}R�Lj�b�χ� �~�\ʕ�u�@�0{�X���n��#E����>{~�p����!<ޞ��wTA &$��i|�ߞ$���W�h���$p�w���k��a'2s�MO���
x�>��c�t�ܯ�Q�筴���Q��
��-\"Ї�Gi˖Mti�6���ؽ�6L�}�2̤Q�8�4UU�JhG�a(ڋ�$X��ּ@��r���K�\�^�}W�{_(��Z>~%^�[�����J#��#�u�	�V��>�����E�3i�M���|�i�8 `���4���V��7���퟿��*еy~����qF��	��d�W�&�ezk���K ��!�}���+���V�r�+~ ��5q�E�+6A�ɏᇴ��y�8/�ɠ@�
��1	߀Σn)tό�Z�<Wߝ)ղ�x��p�wN��$�����jVa #�E�U5���Ҿ����j��_FH{���]��{F�����zD�R�;?oR�B]���
F9��_|�@���4$I��>�;�
��'�l�;��4j�=x� .�|�裣�.	��fX�7��������}���=��l�����.�u�X/H�-�5`��Zb�A�^�yGP@�����	� ��Uik^���(�i�$�+���jE��"���>��t1�fc��4������AFxK$���BL�\�E9*���˗ln���C�e�u��`��{��e`�� ��տ�h��b�l��y�����=�@0���b&Ya�	�$Q���*��Q%R�����}������]�C�n�1�䓏= �mٸ��p�k��
D�ܒ�9���h���5�.E���\Ө�Z��у��|�o��:9r���	d>ʣ�2�
�a[b�-��s����6w�l�q���_8��!��5ޛ�E��X���#v�#v�Z��g����b7�\ˍ�g�EuIb��_+��g։S0�>�<��_IR�3�d,t_0��W�?Xp[�T	.e�_����1��d���,G�}�ܓ{�GϹ�P�K�ـ,�����G1!̻O>��kt��Ta. ��<ZJjz���0>�ר�/��b�(�!�?? Y�=AT��	c�[�I�v��(j�--#�����뭠�y�N�J=�{?A��\<��g�u��2���}t�V��-���K:��B������9���VS"����:��ĺ�ڄ����tm>6v�!���n�XΓw:��� B�S�l^c�
��Ǯ($�o*���+����L;v����K3��/��C<P]�I2̮N��k?�0����?��i��a"��?��?pj�ƢC���@�#��R�|w{�,������/�Kf���8E�N��^x��ܫ��u!
�bн���̂�N@`p���� ��� �ܵ�^~��/��/�g;܀��ZXK�0��h,�%_	%����,'V(�3�g�ݟ����g7�#�$mKw���]R�M�ctb����)YVz9w@R��K/2�]�c��%�x��kS����+?:����-荂;�ft���?�?�	�7`)4S�϶ �����|!��E{���i5�B��'TG6Pmd�*CU�bM-Τp���)�Qȯ���W��y�n&_h��@݃:YSwnq쮨�TP�I�c~\��Zs
"sn� v.k%��7��q1�7'�*[9b�<�Ķ"��7�BȚ1�7��@�]fs%(�kxZhV&,8X�~�&�� �-�8Y��7z�E�s?�`�ňk��s�oߵ�>��]�<��8����b������B�b���[���g�q�;��!�O]�. a2�:�(�[�lv���Ŕ���������Hr�co�����d���}����3���?f��w��ʿ��=UV5a���� Qƶ7�瞣7�|�J����t���#!X��u��\�n�FO>��s�rMt�L#f�
X�o߹��}�UHT�����Q(N���ٳ�-���Ez���\nnǢd�G���;�%k�)bzSKPr�%}��z��8��Z�*4���$�C�U0cSb��cؗk�G͈Ǆ�jePBEM3�]�[$B��(xb�(ߓo�V8���X�e�]�!����%f��رnPm�*��ԓ�!<ds��g �C��V2�ԍ�����������Ի N'����V��Y����8��M�4�	�+�	{�N�>@`��`�FS[J�QS-�<,ss�ad��S]Nq��hhN�@l���j�5/й�t�"-�Z���{z�ZyĶ�6�Ө��l�|t��Z�J@��A�c�j�V{~C-Ypr��
{�7�w�����&ĕ�&'٭a��B����[�w�H�ꊾ�co�&fcpr?!oD86l��z���O�m��Z��'}N�����5;���(2��N���1�OB.6�eT5MN����8����;w2Y�G?�?�XҾ�GD��<�$��KU�H(����Q⍿T�AȿU� ��q]�Y����I����'���i7���G}L?���hמ�<FPb^y�M��*�h56�#�`V�es��(�}�c�l|:w��<������12<j�Ν���%J%BQ���wNx.��0� QN�%�7�J���yg�39��RHȳ^A�+�!��:D>�(��Y<a��F 44�����*
�;.���}>���(��`��yE�Z�4�0(�6t�}���y��g]F��3o�m>����FI������mܴ��!R�2'�͂��Ug�y�,,p�}�m��DV��r�:C��_d��8o�7��\�*��]�_$�@O�š�y^��c;m���7�}����q�R��q� ��R�5!�MV,�O| a��Q�%�P��l uk!��s.Bl@q7-QZM��I ��vŚ�&$�ɚ���-97���S��c�{�1�y���#��e-Z0�1 D����ߞ���r��7la����-�-p^�꺉��t�87MB�ӹs̽��{��}YX��=����z�q������m�{J,�Pb���t��a�ꫯ�;��g���A<D:p�B��Ul�x(z6��ÊXb��3���/�\�Y�ġ��S�0 ��b7�Ii<Y��>c|�ٿ��c� �э-��Y��o�LV3'[ (�g~���jtd�]�ж?s��ms� ����O�{!<H�#F�3бZ�ys�%F��bWh�\G	\��^$�D8
��y�@�X�7r���O"��hW���:*���.je�ñ��07�Hӗ�p�Hב#��m�����ԋ
��{�ۏr��;�A�bXo�t{��F	�+}��}(�`�q��m�� g�����y�u��Jm�t����򐴴�JZ�����w��o���H��a���U��A_5e���u�:˅��94n�[˖B(��`r������@��������\�O-�vե����9�٣�Ll~�����|�y����*j:�	���3�DD��j�
�S|l���>�(3�1���}��,���������7U���u��F	%s�]��ء�};}f2FM�����.w��)���) ,a�����˟ܴю�lğ��	\c���?���c�<�G	��g�����2���-�PKq���
 KJ��<aA#kM��wC1
f��n�!<��e q}��2�Q�x m�t�����m5?#3!hݛ3V���0�8+�Z�@��%��a���2�jnnZ�ڒ9KI窌)�E���_��@(�N����ub��(
9B7-�n"� �m�#A���'x���`~1#�-У�n�lI��.��������}��t$n{x�;FI�a��	�0A�n���t:��q��A��v����W�}:p��䄵���o���T��T�y���U�k��~�
 0��� �����z^�J��$�s'�0���p���7� ���5��,��o<t���#�]԰��m�ty��x,��6�k��̤��[����2	�Q�q^�6��>�}$r߻�t}o�tT�/*��N�"��Eѱ��`$U�RW#
��~��LW���/�Ə9h�W��w�u��;��hcX��E��[d�6.k��mpl6f�n��%�+���b�e�TG�~5?�_���S����H����SO=��e����@��xk��#�i|t��o\����8uly�1NN!���^�<�J�̽ar�R��{����g�g�	���[��r |�����u�7�ۀ��R�B�Ԇy,����w�c� ��M�"V�`�j�,��@��o�C�v�c�N��o�G�N^0s|��c~���D	�-۶ҭ��L���r���#U����yԬ����;o�+;e�-�[p">�c�N�t��c}��q:s��x��q��H�0�@���f�@�U�����4�+Tf/[^����R�Q�(}�C�1��>;s�N|q�N?ƞ$���渻%:��3�?��0_���zanT�"]�N7o{|�9z~��7<���i���L�m>XN���R��x��Ȫ�DZ���!F
k��;���qb��X���O�heRޠ��
���nآ�>Sb4���Z5�a�BA �^��"[SA�筳�MR�3��������1T��A�6C�b-t��*xO,�%���c'����m۶�����o��x`��Jq8�ҼjZ-m���B�ǚ��)+냧�9�=<���/��0Ê�5,�B��������B^� ��ǸK��<���y�4d��*!�B��RŲ̤Al�*,pQ9UJ�j�;��\��_���UQ��~@w��MV���w\T澉��Do��&'�X�@�Cq��|xLZuV֞x�1z����{��g�����y�~�+:}��(ֶ���p�����⻴qb��/+�y��$��D�"1��;o�m���_]
�nh��t뭷ӿ������G̽ч~BO��7t����2}�(��X�{gd�no�e��bF�u�g��T�ͯ}Ms�SeQ���6L^'X�^B�(� R@������ 0��O4]0;~��>к@_���z -��|�n�R��{	��F���z����'k)���B�_m|�w�qB�����l���I5��	>[=
<\tX���Ҥ��W���_-9�X:�44u��ح�\��u�y�Yw����s���!�b��Q��x���1B����`�k�1��Z��_�87_�N�j��s�	V��x�;q��IF�C�a#���F�����9֬ա��=<�+3s�7��q��|�s�ò̩���+�|F͑ge�����͏�أ���d2����ݳg����,�F}�Ν9�hup�3R�Tr���te�­�JnP �T+ClAJ�������,�<=�x�$}��~��ª|πL(#���esٵ�Ιf�C[�o����7�t��y�x���p	͸�~�0���ߧo�[�\`�oݶ���'htl�����V��%��́�o��-�r)��@y�1cO��%��,6��H��� �iP�X���y+����-=��c4T7��Ҷ���3��禶�[o�A�O�kC�!�S�PP�+�$Is",�8��~c��𞬕�Q^O�3���5h�^8u��ٹ^K� �u.r�y�z�m�ښ�L�����o	P�	r�m����?�����Va���k.�.Zl����욇{�����L���+ȡD4j�7��J�ٰ���k��Ɩ�Z�j9j26#�G^jr�Wæ�j;tt��v�����/$6�QpJQ
�b����#�ˀ��KS��Z���n߹���S����+DP>|LCbs��ޅE�s����ޣ���o��6+GH�C�V�0��|!��7���0�����u���\./{b/o��b3(Wg�x8�׽p�2}d,9Ks\	��d��(�s@�"x������PNpmx]����U0�8�9�P*E�;p�Az��o�����x�MZ�1J@��p����@VQjcu�-�u���5��A:�� [���Ĩ
�V��X�cl��v�a���H�Wf�83g���M����q� ��t�`�7���~׌��_����Μ=e�-,6�7��4��NQ2Ϟ�\��������3x��?�'�~d,�WG�p�}�ҿ�w?�C�ns^5}��r+�����-b�)7 �xl��A�z)ý>��8xD��qJsյV��ƥ����H�������ɝP�P�Y2k�]��z�
BL�
��Ely�V)q��P@�ߩ{)(���UcV��O�='�"E^+�1bA�<a��vy�R-	U�0�n\]�	�ga�B�,X���cS�*T�X�.6 ı�mÒ��J�
�
���O�'qh�fG��ė�m�IQ7��e�w! ɖXlK�\� $AZK̼^]2HX̀ZƬH ��R0U�ٲ��*Ooj$�M��m�i���f�K���],��x��������O�	�]1�Ĺ��|v��#n���b���h���F(^`������^�l�\���R����.�M�A�?���_���;hfn����C�_��c��# � �Zd+k	69峳V���:|�6�;q�������K/�k�ըA�T�U�,ā��%����%/�������I���"����{��[o������bK�R\x%
E�ˌ���7���q��[���΍o��CՊ���\#qS($|�����˝�g+v�"�*9O�*�~��A�\s���iz��Y9j���TI��@��E�:���ʹ}�.&䉨i��]��=E�}�a�ڰ�(}-�O�"˥!�����G��5�?���N������_��?��FjU&Tٶ}��.G
J\���7�a2 �c}q�>��(��^��x]3�y��������o�u<</�6�E'�ƍ�p�(DO��h�~���S��H�cÙ��V������=�+gZ�u���W|)J��X5IC7�.��B�ǭ�̉ k�
�������{����: zbNՓ�0����n�mb�]���z;l��^��-�"m�oy�����m��.`a�]�"p(�J�8ӗ||=�d-������.�R�" ,�0}i�7�PA$�2H��tSĴ�T�/��T� 0H����(��֣�?���Yr�AQF�&Hy
S�˰`��s2�S������mێ�<��^�4m��ev-� 5sFS��f#�%�w�wl��l���o������8����W7G��`��C~�j��t���4;?ǩc�ێ�'v, ��#��`|{�9��0S[�8���������:R�pJ<2M�(��O?��Q�?x���<{�In@���7("x_5��K��0	(�m#(`�>��w�P�왓@����Vb�ĺ���<��.VK�#�Y���(0/Oӿ������̜���Pl��]���?��8 ��O<Iǎ}n��
����}��Ǎ0����g4`) EF)��BQ{�[�de��\�I�2u��1�!m�( �#���ؖK5��ӫ��Ί<_�R�V��s����<n���@A�9}�$[�[��`,�����?+?n�<��ܳ.��=a^<�	�?t=O�Dh �L��|�*N��?G�o�+b_�܅���.��#N��a���9�����Hw�J_����r�/��zm4����&�K;�-,�ը9�R���J�@Y��U��c�q�����Յ��W�$���u��"��8Z)(3{Y��]l�:�y���#��-+��Xܸ�q[����aڹs;[��N��>CS�? #�5�)L�l�8��W"0�WL2��窞��޽��XXi.=3�
�S��$l�K6�W^z��&&9v
������z��}|,1��a�KJW��{AXذq����crC��Z�6o^7S���1�;v���!�
���aV4>9*!��S�qiq���}���w�e �����o��C(|����J"��ˑ{>8ni�Á����A�k�^�	� Wm�h}��5�Cq
����MT�m�
�>'O�fw���1��[���x��x�M�{�f#��=�y�[n=d�����}�d�`X��5��t��)����&��M7�G��\�����c�1�v�\�2�<�1����lR�!�c�F[k21������ʲ��}���������v���������>Kfn<��C���(�(���h��E�b�h��AP�L�j_��8��)�3Y�g��z�~�� 4�YC�DC�9����a��	5eOq.��v���hk^�3"�z��T7R��H~ҫ0W�X��Eͷ���Fʃ���K��,g!�`X�����q�&�閛inz��7l4����˝�i�F� 8l��)����(G���)�����m<�	X�g�\&�&\��k.�n�O��(�X���K�����'�ޟ��ט��V�+W��E˦oiIT�K�hm��p?��Oi��/��07o,�yڶu�sϜ>ɮv�0��Q���8v�z�g-�W�3u-�K��#���,1��+�Jn����x饗�\�wx.^8G7l�J�O�'�?�(nM��VcE� ���(� +G�M��v�s���
,�"����a+dX 50(�h���8?�t���4:�[��G���ۍ�����ct�]�h��)��L�N#�_��@cFA���'�T��2��b}��՟��o��Gi�6Bqc�B�����Q�Z�D�a�y���I"=P!�����t���<Bv)�:F�����l�� �1f~�����%1�b���gO�_�xN�B�.lu>=��U�gM�{f|�8�5��P�n�����s���Xp�|7g���~l]��B[�}P,��ȝ'#���}z?��oͫ�P
-�X�d]v>ǒ���eo�f��v6p9P���~�`6(lX��]�/.p:�а�tl�
O Y��Z!,n<-����;l�> ��F�1l�\2�ai\�F��Y�7�*���Ѫ����M66��?�ͭc��?�9m�+�S�oô8�V��L��T�#NYA���(\B�B]v�^���+R����+�̪�h�n�LP�9���}��~�K�yr�
~f>Ul�,����t��2U��m���J�׉-_92 ��pIX���x�c�p��B@D���bmCQ`%�,����PV��.� �\�Fs�����ZV�Ӓg���il�TfW7�����^��r����5�X7'��ۻޘ�q��1����&]Y�������'��Q���ض��"�$�s���Wu�c=T�#���l��&�/ z��p�(�7M��吟!�r#�C��o�+��x�P�\�e�Y��a0F���z�i�,H�R��Wi�Z�:�
#��+o��դDXBE�*�˼��s��tރ�*`�]�1��v�^�Ie�$����W��y����N���|��`/`6�o�?� ���ŕ�&�����
U*r�a]�ܻ�����;���Y7�4�j��֞�0���U��F���pl� sA�c�C�d.f�����U��h�LS�4.��;Ȣp�d)K�n@�t�[�K0	�Y�t�GSN�2��ސ��%��6�@
N��b�̹�%[��1�[�8���0��c��r3np�<O�;T�9��� ���P+��aO��L��([���2J�xP�*0M�����|S-U�8�ke@�T��M��2JVz$�����#gӚ"���se�ZZ>KD���ز��<B��o����E� ��!�ҔJz� u܇�C�"�Wd�cь�bQX9vĬ�vS�Z�:��M����cQ��M�� ���hԙK��g�	E�c�aޛ���6�I��4Jd����%A��ˬ;^ݮ}N��t�� ��J��U~1l�ng�4��Qo�U��wJ��PT�d��@�ƠT)�D��U�ۗ�ּ@��^_mϏ��
�B9���ϣ��%�5-�ݱ e00���rD���px�5�-&l ����SN���X649Ҵ�*TZX��σ�]�����{�gI��N�df-o�}G;@BH�HQ�%R�p$J�=���#�p������;<��P
I�)qEP�(� )���F/�}y���Z2��w�=7O�ʪ�^�	<���WU�ܼ����x���q<��sZ6�"k�� �as����#�ma�NKQ����=I�k��^x�I���,�_o���qr�(�.�.��Os�;>|��!�Bx`��s~A�ֽ_\��:!�������`.�*�j�ʈ4�O��\�+�x-6�V�A�I+T����*m_כ0��ݽ��PL�-(��[�IuzJ�I� H�\ufjj���6�kB�����2���#�,,N���Y�<է-6��ٿ�J|E����z�5���JW�^�`�[4
f�䁖R�,��C�\[�sj�i��/=f���)˥Dj�\�V�	}�쏜��X��Ah�\U>ȎT�c<�T\9eRxWV�+�%��>`���l����c.g9�
��� X0r_�m����,�D!�ո[����UZ�] $/�"s&��aX\�������4��wFM�|y_�L���,	A��q��sE�Z��w��p���?���~7Iߝ9��QMwa���ϗ�,��ڤ5�7���	�M�]����_c�u��k[b^z|��d�߶g�e�)���V[��k��c�1Ĩ�8JTk&[mG߭&�L�����1���\����V�|iy0ٕ��)�`Z6O/01�T���󕫗��C�E0��)0tl�;ﺋMvo�����x/1�V����`vO�Jh�LWZd��&<�����̀(��gJ��[����8�ؽo/=��C�}h��Z��}�vƚ1յ����Y�@�>���'�!�)�9��9#�*A��;���71�WC|�RR!p�f�p��w���E(C���~���l:���cnU�DZ�l��]���x�Z����M'O��@,4p�$��0��7�����pj��uk�~�8�ܹ3t��S��К�֦������-X�֙�B�����X�9�t�.]8O���R�'��A(�����=#&��L�-����@����Ъ0Cy�.��;���w����9A��' _�H�.]��A��c�Y�C{�J!��e��KR��6r�MS4��n/��(��j�h�'d����`]����a�Z�`�K���P��N=h�(֒��޽{��8~8||�ҥ��Zr�]��w'ir K��$ieN *���c;,.&}��DױI�;LPH^���:�_��=�
�S`zlj������	���+��+K�B��@�!Ùk�(���J�N�i��R�Z��=�����qBӎ .�آ��S�
�˲�,��U�öܯ5�t�����[n�.�^q7lvml{�N��[�,|��+�S�G����t5ٳ������aèI�Z��%Vߔ�� �br�F�*S�/~Y8s<�r�xk�Z1���\uYS���O480A�k��f�`Zؐ`������w��|�믽B�+7$b��r`�����|#�B�C�Z������<���+����� Hd�1?��6\)�Z��Z@!��?�C:v�#b2��x��f��(l��W��]�� �_Q� ނ���t���gY�L�*cA�����Oh�b��o	D�"B�I4��#g��࿤��Y������Ax㵑��%w-.��
�S ��\�)��(�:��� �4��\�c���e ����-1�1��0���W��=ē�t>�Y�~����c;�! TH䐃�v�X��Zn.��%���N�����Kܼ:aĭa��]w��|�wŭ��wZ3c �3�A��,� x1(���Nh ��|8���!�9��[������o��|�fg���s;���/�}�i�]�q)[�s����4Yu]�r3�v_�+�5,J���yǳ@ =���b� �E����*��[�Gm�G��[�U�r@*D�p?0t�;w�}N�J���o�*��Z�%�Q�w)�ֿ���=
x%�c���5���[�c��EuN��%J�k�3�bW$�,����0�~�wۙŘ��v�UT���8��y��\>���q[ts�r���-����	k�<�1m�3t��r�nT�?Y��	�SҬ6��a�h���ٗ�p뽬�.���eŨ|D����R������X��SJ��z*�߼PS� �0��@��h40Dlj0s�P����عT*4�t�Ǿk�w4�ͶI����Ě���m���;�C�oa��@tT��{�O\��"4������U{���T���R�Hyq�%&[����,�];���}�
��u����~>c,8��+��0益�^Mr�+���P���{�>�9��l}x������a��"�{������|�i��sk�a����ӂ�"|��}������<�.��ګN�[qs��v�1'`9��������m�|��s�_�נ���B��fG�8��9��u�0���_[��_=NW/�g� i%|L�YA�F�d���J����@P�Bu:�J���	�e��B*%b�kLHp=��9�l�	L��s�QKy�z�Z�^鋮? 騫O,X�
ܳ*���������T��-�qVՑϔ׎oj�h�g��Ɩ�X��ߛ�7k�m|���K����
�������O�9�Q,�ۇ��'e9��l�To"�ܕ����T3Z� D��\�������1�y]��T[���A|����5�DSeX�_�{򻏰F�.?���8��~_|�M�%-%=����f߹$�#�g�Oc+'o�1<�b캟G�)��,*�Џ���!�fx�p=��3� �޶��?��q���¼��{���0�����16����g,��`�l�eg��a�A!B�MUVb�^��t�g��8d���ǡ�OQ���3�/e��֘P�և^��"9+k}�z�\J�(=��&W �������[��^�u�m�Y��w֊��~��5O�?��63Мc���.�n�Bwsѝ�f+���Wt�����4�-o�idbrƘ!���yZH��� �TxT��:*��o�MQ2"�H��K��U'8t��5���V�����/.�
�u�Nx��u^����Uv��ɺY�(H��A$���&��T^O���}�h�2w@��`%��,��yJ�����֩b,�T�[/y�V���G"DW@hVXT�(
��nӅ��u���Ҙ��M4~#�c����wI��6͸���kι����W�^���|c��}HzZ�̷����[So��Z-K��UR��U�����V�Ƶ�>���&k�2b���:,,;6x%��L]m��M��A�晙�O`&;��%��mjfh���kĦ�2�	}��ƎM���g������`$�6�u��п���ӛ��N�����r� @H�|Mkf��SR6vP��X�&w�|���P&Ъ�̛,>�-i�o;�j�iׅ&��i��]�.�diЂ,C�T�y}m���Ew 硨���$I?J�B�����'�%1�dV��l�5�>Č�J�N{��l���_z�_0�á�o�^ڱs��GqV��e��z`���O�yv 4�A��D�&w]�3���sw�〺^�iD̆�&�~�+�v�;m��FI�LJ=�6[AXprڿc�(��?XӦ������ $��·r�W/���X"Ы�R���J��Ǻ��� ��n�p����j�1zo��������uc�д/m����1�I
UJ&��$Z_M׈��8Z����1lK+�5;Fz=��竀�͟;�~޳٬�Cϒ���>�f���ɋ�\�Z��\�yj�	~C�a��Q�Ʊ���Se��ۢ�y|e�0�����ėi=�'h� �!�bUZW@�}p.6ҙ�G�c7�}�G��I�ˁߵ�q&C�g+aGmf�{Q�[��h�����<��>a�����E���Y�LR�rBC��g�V���*G{���jm��rg_�c��Ƨ�i�gO?�Aq�G��R������렶x����d��X�b���q=H"Naj�̜����˟����Ғ0��y6����^����ӏ�>6��T�f���/��*̯`Á���Z�T��D��J�o���+�R��`r�X�cn%tp�^�w���i�(Ltc����8g���w�_>KW/_q���֗�hݍA�<fr�i�m�R�Rܘ!������>t`�ǌ;'�Y�@�U�Чi0\c`�)�>��>�`�x�N 4W��e^��� s��s�܎92�R:瘻ڱ�`׶�w��%�&g�K�q�.U����[a��eο��033S��Kɷ���1i�5���⥭Q7�
.�}��r<��yj�l���I���׮+l�]�]��(��#�5�����k����xf��n��ʍ��m{�����b:��2n�yYi�UY�t�gnQ�b����~5-�b�>���8�k�3x����p$��_����j�!��$�>�2�2*x?v�%Q�i�k��%n�=��K��[���\6��9?;� �E��D�`��E�N����<�� ���[��0�@[^����?Ϛ.*����$�%qU.��?Uݲ^M�d����p���}��_g^�wNφ��]��ŧ�!(N��b���4AX]�"�B��F3k1�f��b�;�Y�6�bm�����65;E�c�\�F �����w��;��i��o�5=��S\����|ܼc�zm�;z72D��S��.qʁmnO��-!Э��F;�ܯ�p4dm�ƍ��.H�RD(�}N�*��e5�kf�������r/�:�~�҅P)s w
bX�_/B=�O��=�����!�͓�i��eؚ�fᠭE)I5�#�͏�\���=��DS[SØ�0�M�2��~����s�̮&Z[Vc�0 X��h�q}gY��g%��hoo[����p8�Ԧ���(�x�<��j�qP�2��R����AHL�e�8]��D}��a�A2Ն��\ee�eB=V�T<�McY����O��$�Ėѫ��*�
=��R�I+��x:qjO&�x)ÒD�o�7�;��m����ԛLY�n��D��kX�%�H��n��Q��_�ͩ � �Ϲمp}0��v��"(��|j���Ř����ҔR˼��'�2,<lj����j��`��p�I���3����7����na���>f��f)�����,,�,�/�S�a�'Y�D^-��͸}"F��f��-�������o,���ԝ�fP��%-�mM3
��ˋt��iz湟���!#����"(/>�<�;��^�-:u�8%�Tp� �ES/_�S'��?�s]8�����j���F�;�+���!�Ԕߵ����˜�(z$c�{V��Nw��,��'?�{z�7hm}���4�5G�;���?�n�gG���ז<C���cm�&,�iXO��R�����h�uZ�������b}�m*Kc�dd�JbBa�ku��ut��-՞��C���o�Uцf���z�u���c�q���c��1}HӤ�7��W�z������&ڶg�05$f�c�h#��	Zf��M�+��Ԣxi��`��r]e�4�Qebl@ݐ��ZV��޿���O�Az��ʆ�(T0	��q}�� f���d���Q��/-����CR��o�\#�#��f�(cӮ>_�&�"z�jn[���j��E�~�;�����	�d���Lߋ����8�8�wZ��R
-OR<A��&���~h֐Z��U�f!��X-
[K+�o��]�����k;X}��
$�^�D��
g6��2�;'��3�]��w.���𜗾2Xs�[7OD S1je��̺�{�+��ȍ�0����9j�t�w�s	XZ�x�C��	I�EeJ�|�m��?�S�^��S'ߥ����L�i�K��Y�s�ݳ��o�5���x�K��D���\�z��LW�3T��ghu�����+��S�ҷ��]��Ϟ��7��N��>3��9GN h�8I�^�6���y<
��Jf�{2��N���t|�`m�5ݓ EP��^�z�+�� e�RU�Kkn��4�Y�x�>,���2�ţ4xO�O�_+a���T{پO�ԫkdD�����y�]��%*e���&�ZJ�5MR���,t[����,����{�k�'���zq͑�܈?��اM���ЧJ��jV�̒�����D��w�R�VH��y:5���'6#+P��w=��%�8�#flJ��K���S��)�i�nǙ�yS�U:	c>�	���q�i�s��4/��YC�Y@�Bۇo���8������yO���Ap���Y6�x��n.��1�%醅:T���>�,��° ��k7�?�jdо�Y+RY�O1C�z�{�F�4��%��n�����w\�%m9��-���ʊ�O�7�Lh�<�E!L1Y6�D���Ӧ���>�V�f�}�'�"&�da��n��-�ZL�{v�bA��|e���n�|�U�)GP%��Y���Ar*+ߞj�^�˃�jB�m��B		�ϲ/vBn,/����Y���ziY�|��9_�㉀ѡd�sNC��XI#u�pїD��.���z�r]��U�1�S:w��.���q<4bd�@����X0z�i�D�Ҡ�#�R��+(�����:�������k�נ���.���a�����<|6o�$E���D]u<^3�U����F.��W���E챎9�V���{<�ӀZ,���ȳ��:��f�M@W;���vZSK��c�$o6���H%k�tk1u�"G[Xx��<��{R{Ox��q�k~�8�0�)�wY�	t���*d��&��"�lH���\m9�|�r8�=�0�����o 7���g�W������.��eS�h�m�3t4�í���W�շ:rMoB��&������x߱9�^/�K�D�K��-��Y���홡��sW��R����ꇕ{�>�����]�4�ҼW���mV�S�z�xO��,����&�ڱ
d�	���Ƨ}�-���^L��b��x(�A�aa����:��y�̜���e]@AJ^�f�xmZ�����}�ZLG��S�[�t�����أ�>Jw�}w�5�I�F��B�u�Ux`^۝v��8��+b,�!��)L�k���� ����ƛQ�Y87���u�LFܘ[n,� Z�z�&am)�קTֵ�E��������Q\h%#ڛ�깕�h�T�2�!�_$�F���,_�i9�СK酺fx��i�K� (��6v��Z�3�>�򍠭k�9�\�#w���Ϲ5�y䉬a}j��q�<�<j#��H�J5�}\O�����թ��fY�Nw�J�$�eٚq�ͺc��S�<)���@pH�~�OL�Qc�]����R�u�Zn����r1����^ד6w�Q��wC��K?��h80+K���o��u�}��T.�����6��Zu���ҟߒ�$�C������}��}�k��������=�����ÇWi�m�3�5
`*h�o�~��K�A`桽�dυ0�>=��g�P�R�g+�2yմGM���f:��
Fu�e�����S�
����T�X����/ 35?�&�Q��Z����O<G�x�pL\�{9�[��A3����H�V-xK�\��n�=�/6�r1u�V��Q"c�*Y���e�%���� ���5q�r��=J�9)R��l��S�	��v�nf�����@�TR�:�u��"\�}.e�7��Q�:��7��B�3������d�E51���b\G����AQ��>��'@x���5��y��(�鄞���+X"/�$ռ���\��E`(�4�+��8% h�������C��h˾��y�<���}����������jy]h\8�.	[��7��?Q�i�{�fmV��A7�|�o���X9ĺP���V_e�Efa�M�K#�.8�\����}�T�r���4�`�~Ckb&V�UMH�WӪվ�i�O���'��^�1r������{4=w�@VR�J���-MM���S�3�ʹ�m�5YU������~j<��@\x�����j�LĦ�*m�k���ۗY����B@�B�.c�WLQ����R����G~ d)0$�"q ����"o>�7�7{�<��*�/G?�]��a�O��׭f�"I�J3Xh� ���8�_03���,tK����Hh;�����V��~��n����U�#��~~R����.q*��֪p
�D�m�V��굔���h�~����Cje�(��CI^��N@F����<��%�t.�A��a��3�۷�>z�ݜ�733}�1�W�\��Ͷ[�{ƷC/��ц��s�1X��F�k�F���j�D'1�����js��G�S֙�=�����ʑqDE}���ʰ������b1EgJK�:
�Q����m��5b"7�@�����,��#G��#�M�;w�5=)�� �̗�"%�&i�
*���}?�B�h�0�tA����ud�	�}�9� 9,+��s�D��&�/h�6[2hU��T�~�>�Ļ��L�3�0�;haaN� :�A����	:��Uc��)fP�~�e�;wF#7���Xͽ�%I����_�n�"���Vl�V�7UTQ�N}�> U����"dj��+$� ��j�h�MB�M譎�� J�]���5�V!0����yH�CF�&CU���3A��������v{���g�ӛ?�I��%ZH� pЀ�Ҁ!D��ZQ�◽Gl���ǎ��B�S�6���k��V� s�eX���z�X]G+�5�7<�e���sg��x
��/��v�΃|W�(�ί�h$����r�U+	fy����n@_�;&q���o�cm�MSl�������<�v�<��)�@��r)g�8#ݵ4i����[��3�������BB�Wrc�/����\}�y��ziRYxd���_�l��6�c��F����V�ƴIV�&RSK<�sm�;݋�?�f1�X��0�3��{0�1�񓮱��@�ȁ/�P�v��g�f��#���~��v����9�F[�kP��,lM��	�[*��nY��������d��2�x9��G6+�b�k�P뛜�����4�&��>[4XQ���x���C���iC[�<߿����Ga���231��!�����¤�V�n�ds{eb�J/�?V�VטT�h&hi��๘QO�0�=q��q#�Q�+P%�/f�q�C�3�^^]]�\�>}�s�a~�|��`^d�6����,U}��C	w5V�,�3���;�5�~�mLq�z��<}�Ar�f�9�2�Z��X�|e�D���/<G.��}�!���M�EO���J�����R��l��7�2o���l�x�_1#�LK�d�I�����"�b\�~�� ��-.r���ln���f�]�~�9+��#�|���ɤ������D0�Q���ѻܺ�+h��O�K��b�;���ǭ�����m�Ч����m҂A�@�5 �jfW�D Q��c�ܶ���}Qf����$_�B伢��y^MW[i��7������
���|�����mu-,�r��Q2�KԻ���#�0��|�;<�`�K �<��ct�]w�	s?e�)�y����� hH�Au:�!Xsd��U����`x��U��%����S]Ny:�����=z�W�Y���~�eUQ_�A�:���Q� \y��WӾ�����7ޠ�/���#��W���(�����m�}�B���(f��VQִ��2���qV,�{M�s���ǵ���^���b��
hӾ�i�ŋ�.o��s��A;c�z��ĥQ	�:�z���E�(Æ�(�d;ũ+/�q���4U��td��^�n��h۞�k�&M�,��y��� ���e�j�9U�j�F�f���&��'5�N�5CE �gQs-~�gS���O�G���RT�`���L^���X�yآQju�Q�ce���Y���1SS"k~��Y׉��]�s6�}��p8l���G< ��|�-��B��`��ڙ�T��u�qMh��;��:ԏS��h!{�'��r���,��Q�����i�Ao�	���K�/���"��_��:��)]q�s��]�Vv��Y���@=s�<#�A@�h}�\�`��  ��IDATpZ<��;����&��2��@���/q�����]qE�+�"��v(�Q�n��}R����j.ۤ��Y�&�k���������>^˓��� �I&���-|+��+$��(�u^GX�X�81?+7�s�Y,��~r�M]�]jeQskT(�#���2
�^�u�k�Σ�hխ�u����&�\kCh���k���i۞���̈5X�j�&9�U��K5rhU`�Z ޱ ���n��`�1�>����z�Z�&���׌��pf��+�G�K7��5�6~�x��K|��5�I��)7!M��4RyzR&��g5������8U���c$.Tز���o����eRA�N{H\�@X���~��F����p���H��a�UJ�'nj9X�Tؼ����	����+|�}��K7�cM���KAs�<4n�Hhu;!�Y	6����{C<�h����?�qz���x�/��?��>��g�Nך��+���:R�H���5.��h���"0��쭭��i��.#�4h����E�mD���ip�fiV~}���������hV��bV�ڳ��n�`ݡ�o�]4r���	�+��\�t���v+۶g��t�� 2��a�z" E���� �����:��{虹~F��j�T?�Y�ku,%�z=݌�FU��Z��7qr���vЌ�B~p�_�f�3�$�Vs޹�����L�s��� �@	����	�ռd<
��e!x9!!Lۻo�������VVE���FOs���
������:bB6���w=���Y��sჾp����s}�{H��x��%���t?��X�|��HM�d� �xrоA8?���i�.��8���������a������S'��J��s l��kw���E@0f��9r�c.p�_��_X��e<�����#�e$u�˭ľ�m	�[�ڭ��{ꗢ�h9а�V���P2�*)���ZE�7\E�O��5�n9=O����]%�E����V�3�a�͍I����6W��X�s�Hpss���J�Gy�15U�7I�v����a�*�6i�b~��-�رcLA,�|�8�"���'����x�*l7K0�RmG#�5�ަ��
 V@���X2�u0{י�V�K��Y1٭�"�g��b���U^|=l_�@ ���=���:��s,���4ͥ�e.!���1?�\���aU�<�2��0�9������m�ֈu|�EHK�(y.Ae�h�2iQX�hP#_���u&z�n'0kN���`�k(�}��s�s��Z��X�����!�\�r9������r{w�%�#y����`��57=�������Q�
\%�\�����&:04&}�m�f�����1]�L���(��>�-� n���X��y�:���"zX�/#�:�U�gu]k_�D@���[K5t���\}`�@���K�[��U>���%/��|�����ڶg谵�w�FUD%�M`"`�X��n��f��]z�ET��&�o�el�\�a�?���T�Nͼ���Yӻ���݋�۠_�a�2Z$�F}�
3�z��M%�W����K�����"��R���U�	�Ͼ��.�8����⺀�5���˳���g�c?��`�A�u�OM�֜�sc���IʜH��)�Z�{��qriZ���r��})Th_(��u�u0,�"^�Nl%`B1ĠI�v��=�����),�����$3��"�m\B.Hp�(�u�l�4�
\pgP%PƂXm^��-*�����x������k���4o�ǠH�������R.V��j��J��`�I�W�7�%A�VV��ʕK�3k8W��y��p���}pݢ�Z�u}I>f���ҺaQE�s�`I�{���ҖT�C�ͬ����/��Z%Y4�ռ��m�3��ڮ�O��3��v��w3q�#�W-]}�jbO�:�3&&7c���e�B��e����(�	f�1i{�O�XE>�����4=�J��clh5�H��͗V��ߌXAl������i'-��dE�!����-|Xz���'�y��2�Ũ�G�� ���)R�@���k+lW�K�����B*a�=sF�~� ��Wu
_�}�F�R�+{k^� Gd�̭#D�3Z\ZO�\[�S��{nn��/-�╫^�M�rRTJ�Z��D�I�}+����حW[{c��ܓaq#@�Jc���`���eJ1g��=�L�������:%X�B����l�}X��[��}��ׯi�Mce� ��`�¯����~�F'i�y�4@3O��^�f�D���[��������9:��� ��4�%/�ԭQݚ��b}�7���h#��5�kژZ4��G�X�h��'�G}��ls�5
[�����l����:&���c0i���P#�Ȇ� y�#xԡ~���SO�h��}��J`\�׵�R��)Gӱ`������mM��A�Ϲ^�|\@AK�������KU��K.�8(/	�\&UD�������y__��㮂Eo���*P(1UA�/8��3縀A?8���ʿ��.��b� �ޛ���<^As3��Z��k�淚�eK�`-e�[�6�/G���T��f����	{������a��8��t]j�
�m_����W�Z����w`�zO��^(b�c�E�������OX'�w�����}�hl�J�}���H��}1���m��Y��8m`�A�u�(3s|^rq�1s���3]��i�Vs�j�hM��5�~��1h�-�=G7~c��rUB,4� �dX�;��ݜj%Pf�}b��o�l��ij��E[l���}t.���0t"�*�������t������-:u��f��xΰ_�Д>%4��h�MP䃠�XL=~�7`ߺ�UU��񭷎Ӌ��J��^�0�(�"�\I�iUk�>o~a��u���ɟ�3?�9��*V,���B�M��UD;�;�A��
��zS���G��%4|*Z���Ɗg>]	p��x��4��i��ü?�������s��Y�
�f��_�����?�^�|�^��6�(���{M�Քz����U��a(}�<Wb�i�֥�~�揤�,䙪�P�����k�;EYw��H+nnP�~}e��2T;��ej%y�A[�.�?j}�@<y]wֵ���ձ������E�����G�������o��m��O��:�j\��=�0��	#��=h��+������4J\�p�&*Ek�5�q|l�o21+A��� �"�H�m~�y����Տ��FU�-n�!�Ti623��YI�S�N�Z�g�r���g�g=X'�
%��q��ߴ�^��F��BZX�R�Ba��B&�Ou�0�Øտ���<'~}_d�s�=f���&��7�x�Ο���t+]^yXg�ʜXD�	ڞoc����[��B����=�Myx$�l�	7R�Ж�F�����HA���"�����U!�+�p��W	eR��i�;�
��AACG�nLr�g�Qz�g���/M0��1�q��� �BP�������%�%r�w�ʌ��� |ҧ�N���gffiiu���!�(�������L�3<Bou��׽\��v.���ˬyv�Gu�9b}u:S��%�����U�X믱��T�cv��\���'��p�	�u2�W�1m�s�ܽ��i�ֹ 
�B`�)ݞB0%�2%Zi�!{Y�4Tj�3ZHs*��\�4�@G&O�|`�O�b�"?HE�&R@�]�B��uB*J �x�$>}�ς���H��m�^���v�m�3t�eWV����;�o�ی;ļ�$�^���9��C���bo�Ĳ�1�������1Asj�g-�c)[ˁ=>�5�s�j�ѳ��hͻW��i�N���(̗����5;�em�ͱ���O�L��;̳ �k�k>�6�M ��,��h%=��=,��Yp}�v����W�Yה4��L$�a��{��j9^p-Fע�Jc�G|�b�����Zⵆ��E4�Mf�T�K�d:��﹩iPh��A2��1ܡc��1��ɀ�ڈ2�Xq�23��`G������Ǩgg��g�[�YG#V�}.���߻sg!81���湲��Чlt�g��	���{i����e>����N�hS�����:��y9�����9a��� ̣ω����к�7���}P8Z��^�u�]7�/�5Vq��ú��Uv���ٹP׋*B2�	�A�gL�v��
d(��;���ΈST�_���������CӘO5
y�� � e�&l�"G��O��>s]�r�:�>*m[���u����mW��ժ4u�
�e�%��1���}ffh���\}M"ե+���ط��S3y�U��=�b�����+�%c�� o� ϴϔ��`����	4�"w%I%p�1EU׼Ƭ)���z ��c];B�
z������xQ��[є	f�J�?��Ҿ���{��XZa�bzz��?,/r������}�������_Aɱ�'�>z�|�Qz����Y+�m����W_�_~���%�L���u�
�0����5ڱ{=��'��Cp}��.���tꔻ�[������E2%��z�%�M���sX���Ě4ed3<t��N���u��ٙy_aO��F[][8���0�j�u���ĕ\�ִ����%�����V�t����?���`�J0[>xѠ �p$�;����ߺIԬ�LբhYF��c��uR��e�h귶�1�����d�����c�4Zg�΢�q���~7\k�1��Q>�9�q��60n�q�8M}�����1�?�������>��!�P�G|�&��>K<L#�g��ۿ�&>����4�wS{�L^��f-(����+_��~I�wO�w��=���(����BK����G���{:p�.:}��o�뿥7_y�v�Oӑ;���ſ�_{�St��Qڵ���m�\�}��ګo����{�t��Y'48�
�c��c��/�&}��_��N���8&����kcu����x�~���?��?���<G!���й�6���Cq��4Ւ_J��B�dE�X���$�?�Yh���.��;��*���#.EΔ�V�T�驥@s�u&�&'%&�m���>�25y*�A����i~�����qA��F��l[��I#��D����γ�Y����T���nR@�>VF����p���Xph����y\S��f
M����1,��0yKhT����u���e�O�_�9�����ImV|[߯�²�g�L�z�D����!eԦK"h%^@��<i��Ms�e���#;B_��ߢ�|��"T���OJחo��Z��Ĉ������{�����ݎ���l�W����?H����>���iva����n!�~h�:��0>pt���ߥ��NQgz���^�o����_�N��I}�
����0���B��p�0M��pa�_<�t+ܐ��:���X��\��.�y���	^��Σ:4՝��R��L[K�6�8!�7�jIXk�j� m��Q��'�!�VfLҺ�Z�y]©�%�͘6o��ܶ?C��2s�D"n�co��q�V*�KM�֌m���w��2�\Ƶ���Rfma��a�-3��FmD����3g����X�B���sb|���s�ln��:��C�{+�`��n��K�S�m��X ���B���x$��W�US+S1���Q�?�[�0/v��	���i�)�>A�BY�G��08b�w�=E��n��^ «p4@����&@�����*}��_��xa�F�%0�o\�Fӭ�f��iϾ#n��؝w�׿�/ -@��o��=s����=�أNPع@��9e���\>O;w�_�O���'>�If�@|;��l�ga3�r�`�jNG�,�h�v�=�/�LM���A��W=ȋ ���ү����F3$&���a�e\5(���$���Ɔ�5f�-eT�v{�۶g�p��.T�ۑ�Ơ,�2�������@k�L��<x�����IL�Ik�Mk�k�js��o�g�20�w�9;��j�%Uľ��61�@܋�z|Ϡ��	~����ϊ��75+��s"��k�Ic���1u�c�>���j�H�h��uR���|�����z�z|,@d�y��d���ye&�����1�a���n5�rP`5�%UL��fC���A�Y�e`HkPU�5?#�za��Yk�S�~�����;�y�#��z9�����w��/S7��C�_�����aڱ����(������/?K�<x�>�OQ�i�Q9�<=�����3?��+i��iw�G��~�J'��޹�1�=���C�N��\*�f��
�0���gE-��X��.����!��G	tL=#�Cl��$m�:�$o�E�>V�R��LQD;������b�`E�Lc��HqP��,`��v��9"��su�i����c�v�HG|M��5'���m�yb�b���h��Ģ��몖>������ƚy^Og��e��_��I����h��c��~T���u���G}���b�zS��}��8��������1�@t=�b���#s�`���~J�Z�ʁߟ���4���j{�A�3���=��t((�5H��C����Un���_���o�+/��N�Q�_���E����������XZts��;�fߙa��s/�H�g�emg�[���������W����c�s�k��Ae�e�>��W�+���-�"'�
&S�Ap�������eZ�fuȸ�X;W���}�U��Z�2v���u�$U��'b!W��Z�����2@��}��*��N9�V��4@�f�K�.1�&k��o�9�T�l���V�E<��XejJ�:m���2e�{��Hq�P�E)c�x�6�E�۪ɿ�&�Vme�q ����"ϫ��c4B�	 |�>�OꐋVMF��[L� �g��,�i7��,�^�ro���_˱'�k5v��p�KE���pV�˦<�4zf?o�:�
Z���$�	(}̪.�ˣ�`��RU�W}L'��X8�t�f�0��9&�ʫ~���KFC�5��p��W��K��t^w�����d,&9�ȹ���yǐ_}�5��vBSn\!���K�����{�����/�roͭmњ��f�ĩ���Lg�\`����f�����GO���g���ct��"-���t�����k�2����lIXXpB�ZU�`��-/P;R�Y�{�v`L���E"AAs��Sw�I�!��,���jukŢt�e�b�nz�&4�S:a������m�3t�X
���Hsѕ)¿��e�|��F�Aj�m^0&�q�Þ3Me~#fO�AzTQ���X�� D�[�2���#u��՞'�u��Z�=�Y�3�q��F�ʹ��7i��������Y&���6��M�o����o����9`@�)�̂$���wQQλ���6;-H���s1+�a�ǣ�f��!���mye�^|�:}���NX�wp?��ѧ�cƗ/^�˗�9F�p��e�^w��Ӛc�Ǐ�MW.^��M�3����bk\�T�6e�Z��d(sR�5Q]/|A}V˺�;�%��JOc�Y�jZW�C�d P�p�})��<&$u��YY���A�m��	.�$�5��ʡ��q�;�:Udk6��r� 9��mM�e����������+hJpc̛9�o���p�$&%�Ϙ�J��V����˒1�����Zf�猻�F�I��f��{�O,����
�Q�DT�pe��\0<��&�0���kT�~���b5�y�Y2�\
�6�Բe�XS`���V^��mnf��/^�
�;�����Lϑe�>��^�x޽��������T%+YcL3��!��\!B7�>�6K�A��P�Vn����@����(��H������k�ty��L0�U8��������!�A�9�}��X�x<��R�W�V�V.�l�-�+��$e���T^�
iu�$��U
]���Ӡ��|y#�'�C��t:����d�އVVёM/��68%��"M�ÿ/�k�N�gE�ra�Z�׮��Νe=����4Bm_|+_�S���1Q=w�u�B��}��e���
�VMT v�`1qP���kXR'�i�Ե���j���O^PPF�ߋY�*��9�6��?���[i8���1�?1�V2���@�&���{�}�����ᜨ_�V�����c��97���	�k:?>��ra�U}����[mո�m����'�Ѥ���i'Q�&B-�T��`�{yO���$^ffj�U��3�����,)ciZ0Ll.aҖ�Z)��sm ���~�V�_���A?h���rMzG��F!����T(	�
�0n>0�Y�LE�,��E�����=�A����t� ���h��=�^�)�EɋuP��q�x���K�'l&O����XZZ�gy��`�MR��w�=�1��y'��T�>C]\��W��B�?긹���R�H�6���"�.]:;]$��l;a��$E�
�f�([8Ͻ�AJ]_�{�v]��t�2w�^�$I��Z�*:����B'pE����õ�ױ�8���KIW����n�\�")�_��S蚉�T�O�5�BA�~ʋ���;�Ν{���/���wn3�i�3tV��*@� &IJL\j�fƎ��I�0B�Q���7�&1?����X�S"6�rj5�M���@��{o�r`�g��ro�~��L~TR��ZK	g�R?�<��c�ll����s�1�pt��"�M�#I�s!j}�����%$��wR����Gy�A���7j����(�C����g�~^�vM�FI� L�� �8��e���ӌ�F߻L�V®���&>dx[�u�{�y6��.A�s`$�ǀ���v5��̠��.�:A�ÞT䛚r��;`���q-�Z� Ӵ��6�ᦘZ8��D�7�3֐K�t�a�z;�@��$��yO{M��y4�N��fn9h\�Wq �(�q�	A@��&��~��7���.]�t|zf����a2�����P�cf%��n�ˌڱ4� 2g�M���@��Z%��f�am�2���wf�A�!�{1��� 9���2UM���a�pj�bKL��t�2l�#��ol���s�cy���������r���x�����~��ol��>]Q5],>���8�I��[Qj:7f�u�]����W�V�}��F`�6P���j��w�g<X���ҳ�����4VM�pܽ�����{E�ު�4��>��l����{[db���m�ִ/��.[m
���=�9�g�B���F��{��(?�&�¹�R�B�<Lw�y�0��0[��/]�@�ϟg@���L7i�N�ʹ=rۡ�3~���������6u�-�zmZ�Z�M�%X���ސ�ɀ����p��R^4��\�&��ম?�`ݐtLX�0.6EQ��
������k����jڛ����7�����\�2��u��:����@�bI�.���|�	��Z]ּ5��R�q�l��l������(O3@����^�u����sE���K@���&d��ؕ�7���ܫ�^3��`��Ɯ�^v�>�5������ÂW����Y��4n��qX�m���M�2��XI7>��sU`��)�t�|<�!#M��n�M&��1(��g�>M�����Q&���Ԭ�D5����cƏ��V�z XI1���c���>��k¤o��kZ�
{UИ����|�K�I��Μ}�����{��'�H��k�Z&/��@���m��eZ��:�E�cä�~v����M�p�g�k�S])g
�����~�9>k|-Tx��Ls4;�����Kʔ�8a�+R��Lv��K��I�ӺB;#�i�xf�+�����Hy�t=z��9�ޏ�9+�#�U�m�� �BW�}�\<�1Z�%¤�y�]��
�X����ؒ?�~�>��˘��w���Č �qI#:+�r�|,��H��^Ci����}�0h�v����4,L,D-=�J@!�=�����Qd1mM�\9f�lV#��8�4)��j�1�Խ���6���O�?t#Pi�5�[����m���_ô\T�f67�c}���9э?�������hM�Z*�Ɓ�7�?��H��
��Ki�����H�!��d�N�-�)����Y?Lӎٶ�=��������D.�����o�׾�_�����w���o�E�_������Y�f��n�kTx��G|�Cz���O~���z��襗^���u�gh�yjc�&��S�:�v'=�����r��g�,�<y�1�k����3��.��5_��0�c hϧ�U�>�,D8e���,��	�E� �Ņ]��,�Q����5C��S��1Y�4K�S閘�E�B7n��B���ʴQb��,Ww��ޗ��݀M��$k�#�"id���>�_]����Ǽق��|g�c-�q����)��._���/v�3���)��<�4�ėD��*��^p������G�˒���GjK�a������}��9�?+c��R�Y*�MW5��ڄ�R��Ls���l�Omm��'}N�U͞H�1p����>�g�:�����p�)��N����x@��
_;��m& � � �e�Q�=��ק�y�65B�ZqߋZ!�q-)�����*˰���X�FC0GoRx�[�C����UEHm��E)�	��U��b��0��@8H�(�s��ݲ����+4+�_;i�����6ɸ�5�̚3���9`+UA++�������{�q:��9����;�M��k�>:v�N���iye�f�0��+�П��?���Oҁ����Eڿ�����o����г�|N�T��{��g>C�G�5=�����4[`��:s��P:]����d�����i��H�<�Z��Î�����/�7��w��~m��>ѩ��r�Zfp`\�`�%����+��p�E�Z�6c��f9��N�f�fz���d/���\�\������K� � L�if�-�]�#�h,	=S&�ZL����D�G��o(��8Xk�h�j�NR��Q!�V%5�{}������9�,"K��u��� D#d��[��y��_;6��p_��r`��z+�F��Q1vk��,�c�w�_wچ�m�й%im���YM�O�J�Q	�J�c/ߠ��k�2/b��E�'{���Ϛk������ �`�ġ��Ϧ���x���N�۩e���hrM�,���N1�d����fZ��n��߭��f�D,�W&ō тń95�;�7�<Z�ž�a��� ��W�O`���z�M���z�q�������ǧ?=#���S�����5IiSۭ�z����o9��u����|��y�$�q�]��>p�G�_��'��z�����+��~��:z��ӧO����ٹz�����{iz�C�!����:u�.^���=��C��w/��S&��YX��9�Эip+y��" "@�F�u���)5L��D���z��&��AI@����V�����9�vgTsmh#�o�b��xY�0@I
�T�5ȴ<�(V�0M��!�*���ɢ(0��,	�?~�����q5vM��Ѫi���x��w��)�z�A�00t�L%�/�O�7����]��lԶ�ԹS�=F�7l,F��٤��Et�7���B���{\�p�
�[SS���'-V˘y�ɛ��Ǣ���Ob�7�?޸Ŧ��r��z�o!�si���BH��b��5�[����zL�H^w���ߋ�>��|���r�+j�իW���e��_�5��O~�kz�Vn,���`3O?�4�����g�}�}�X�7�]�g~�4=�����Ҽ{�s�G�.���s�u{r�1�F�;�� ��/�?��?�w��z�7i}����������s�J���#�<̂7��`�FjƼ��Ӌ/=O���ϙ�wQp��ٲ /��J�x��q,���6�^�&2��8!6�%�R�P�QS�ZjfM��B{���S&�y�ު�� fĥ��.���#P���+y�x��mI�h9�~[YNj�/�4��7��ks�Mݭ� .:��_y���������N6�C�00tR��ض��7�jk��4����]ms�D)O��H����HL*MڪH[4��[S[ Hh!�X*�]
��L�6�%��ć6篊��k�l[�f�٨$=��xX�S	�1����k[���?�����=�� ��m�c���}F��&(����IG����u�������������>�K�*�9�C����<�{��d�Y�vt[�{�N6K�|����y����o�/~� �����p�|�I������ŀ]�� y�g?�?��?g�9΁�:k�>}OX�-�竨ii�W�S����"���3�^{�j�<�=� 7v�ۉFM�Ui��^(S�F+t;���7���|oY���Ё]ߴ�b�~g?� 1��$�[�4�%}W{<��l�o��>z���a-p�$�m��wcmyy�G��ʍ黛y�m��K4$�R��'�����"h"�1�q�5i��^��͵���`�S�;��{,~�O��{�$E��}Fqd��������`��D���T�&�����>�Zi2Y��ٖ%��m�C?�1e������5�m\�7� &�D|1����n�"��Ks���.X ���U�"�w7��U8u������iIa0�W^y�:�s����������iqq��f�"�1_<-���}�N�>A_�җ�`��+W�����|�"[�|���_~�e�sGT�Jq��W��o�=n,^e�`��]��k׮:�?��b��3g�я��1��
�(/���L�&��	�:3����1(F�&It�)(�\S�ӥT�A��/�8��i�8!C�r<�E�f1��\���]�l���u� Hc]��~Ű�ݻ�s��Y�P��
;4J��/����sD�5�1K
s� ��_�LB��C76����s����c>;��	�6n��E���ϋ�܋�ط�����N@<���.�&ڶg�D��V��*�$�I�����7��Ǐ�l�lE;�2�
���u8���o\�����hc�m�sY�*u��`�Y������Q�a��\ڪ�TO�66�n��[����IRw�Fk���`_k�v6��ܜ��AH���R�?�V��<e�r]�T���l�y���������aR~뭷h�T,��mz�^��~��)_sZ��hav�&�_]���ff� Z-���l�q�S'N2��я~R�V{�"��,��*]��Ⱦa���#����R��ڊf�lj���V}������8G���
W1�w�;��%>F'	�[U��r��^5]m����'�"�d>�L��0��Kp\�EBa�i��WQ����

-U5U�,S��J�����<E%wN*��Tķ��u����!E�-��q����ܻ�'����1� ����]:�8�R���k�܈ro-e�ֲ�b�}��je}�s�ʬȳ2s�L���fY���w��CVLO��,�d����<��ܹs�������z);����q��+iҚ��J��m��3�O5�Q���zۡ_U���n�VK�����}�Đ�A���~���F�r�@6�c $v�_�MX�0�a���86��iJ���&�7}nz��i��d�ls�o�6:�4��M�iNǅ��h�5�?�LTF��V;���{�����z�/��=}L���6�ѯp�u����`�f<����2������g�Z˙	kpl�1��ʐ���8Z&��'O����p47J.#�j�#5��>`\����M�-����ZP��rX�\7"� ݌�̤�P;����%�"}*ZQJa�����3�z�Rz/�:��e��҉�d�T�xM^p�m�\�k^�|�N;�ˠ��H�l�����c8�C����h����ue�---�����ɬ���f�3`r�q?���Y�=0���Y�$0T�gY
���~w�,s��_��б �J�;M�a�������9&����-�u|��� �n~��N��V7�]h��SS �3l��Ҽ�s�K�{�BK?P4ȠŽ�m�3t�b8,c�,�I�c��L�vӦSs�ڻ�UV��<H����A�o��aC��,6_o�� �����=N��ǒ�8K�΋����Q��f���{�SӺ�6(�V\�#M��{D�څ�@+�]��_ׄj���I5�M�@[���u[�-�Z�3`.]�P�Ww�`��>qTXC�T�>36Pف��֜`У�S�6��XHd�=q���

�Q�Zb�]_�?g��EQE�ǁp���͊���<dQ�@4}6�����ùG�S���9!������3�e�c�������<{��]�v��ÇO:t�Xص����ֵ�|j`�uPHsr/�j�A;� 䇭m{�����v�T�W,�k�n���J��'����?�QY��}7���5�Q栄��9��/�̤΂��5�D�@:��M�H%���H(�3����`w:�<���D�L���+K�(���	�����q��F ���hl���
v�0U�����g���{�uҋ�X{x��Y5B�GX�Q�K�rXAM��c��,ќZRv�iJ�/8p� �+�IWͳ�.1�K7VXD��B�5L���:�sYR��N���q]qDhS}�,#��S=�8��{iv��G��}�O�MM����h=9����3��`a�Y��` H�� g�W0u1��<ʀOi-��%�[�N�FtB��$�������s�ft?��U�W�ln��h�q�W�[ļ�<>g`,��R���*F��f��x�|\+ 3�����G.φ�"� 4zaa�G�zj���St���m�3t4�t�hp�j�z�y�n�o5q2�w��IcC@Bf(JGdT"��:�'Y&�����_��F}e�˶�߯s��2��G���f�&K�8�@�@����"'��l��%�{��5ϋ�=V�e����*_f�M��O?�����w_���z$.%�`��!M0�g��ҿ��g��H0���>�����9���%��~�֙���V�Q�n|��=.wBh��#k�Z�I�N�5�J�h�<7�7�ۮ�n�EX!M3i�b�kVA��o����<;���՟Y�	�E&��_�
�Vh~ys��G�|y/T����#ǡ4A��Ek	c���.# ����;����^�D����>ݛ����K"��Y�.���Ԛ��7��1Z�E��	R3^ʜff�ai@�%l�y��~4�9�l�h&1�FD�*�����Q��e�fW����Ŗ�qMY�0��~�bP&�|?�)u&�es1���oVRI�%����r��Z�I�����Gy��94s�fT��uo�,s��(J�@(¡
�`�z��92��_a��o�&�Bȼ`����E��!�Y���{m՘k����ڲ�� �]J�L�N��T�H�Z�i9�2H8G�_/��X;���M��g�`�&���<ޏI��j}5�ku����S�>qR��jt4�0
C]�����"#�:��-6ĺ��Z;s�+�ݩ+�V6鷃���s�:��APn�[�>�Z�!�մO�����y'�������n�����Xc�p��r��v��E{���>cS��\6���!j7NW�uƖ��>��e0�\=V0���jr��P@���u$~���1f�z�
?e�|�k�������$ռ��,�AQ�zn���:�T!�t����oh���'賟�4�s߽�ܹ؈[�X?h��	�(4&5�BXTf%�VN�ܳ�>��'X(@zכo�E?�����W_e�tMb�:Ufo4�z�2�V�Ri�\���$�5�Y���C��-�Z�����B�w��夲��$�k�5��,��8��5���$�=[��b��=��>��X�����P�ѱ�-�M�G#�(��ۮ0k���������:D&@�Z�b��D�����|�СC���K��ض��[<	����8�jǎy&f�XYYD2NjbT�ġ�8�F���֤I�Q����k@�Y{|媤���V���͍��J�i�i�U�W|��|���u���fC����������x~��fU���4	�lmZc��%�T1���2}��24}W-�i�l��4f�s�Q�����~�>�ħX;<�
}��✕�%a<�rY7��jW�,(��iU���@e�<�ܵ���C�҉'�?�����x�
���*6�}�~>%�k���Hi�I ��m2p�x�Ad��sf�X-��@�yN���cUĒ�]1$���CN���V&�Y�A>:i�����=�ڼZnJ��c�J��O<͂�l�IM�A��Ț��Pm],,v�Ջ��5ZD�'I�Ni�s��2�*�m��^��5�0M�x��QwV�ڠ>�|�Ӷ��O�m{��[�Z���L��2����H�h.�Ǚ\c_S�ߡsfr�[��H�Q�u��fFϩ0>�o�0b��d�ި��}�5�kǌ�Z&Ɒ����[s�ϩ�2s&���Ф�B�^�j����%� �G�	c.t�l|����(�e�5�n4_=σy~䑇��_�������;�����R+f�L��{bŁ���_�ur��w�s3X
\;�\u�Z�2h8�+��Gd+ ������ؽ`���y��Y4�j��~+�$-3 0�L��Իe��&5�16IZw���i2�#���V���q�'��P�4A[��v���_������M;��+>��俋��غP��qѵ��O�̪�w��5
s�Z��M������/������}(:d[e��N��`�F�%e�Z9H�:���(�&2n�q���[~��
yz�j���Jp�Y�3΂����r��U0�T�j�Ӈ/]��-ҜsQ����3󒲝e>O�b�M�>��֘f����ʛ���P�z�
�8]�IG����l�7]s6EH���Z��|�������k �>|�>���W����O~���qmi
� L���y��9f�gΟc�hK :�#p|��4<�����Bt�Ǹl���߿ۙrkO����;�����7������C�O�ڗ
-q�ᯂ��y�q��ʺ@����+'�+ւA٦�U�3cឳ��m{���Y �+s2�fP�@
�g���V���>�a����5'$�n�Tk��㊦�u�BP�U8��q�Q�_��D�q)��'Bd&Y1i�$�N�I+�p ��[H�7���I��鶆���m��݂)y�%U�%�������i֦�j�Vz�&j�O�J��ީ�^E����2�#t�Vhg��[����a��Z�߰��k��)l��M0We�JtF��:~>��q�2�Z�kԴ��`긆M�S�s ��sRu����2��ch���:@N.Ɯ�I:m���ɼhjd�i8v�� G@��-/�҉����3lrn� ���勗��P5�(�I�4AJ� 1Q���_�2����G>c]�$����4O��s����p�;^jUY[[�������4����`��y�
��@L0�?����y����{��_wBf��z���aH�$uAY�{�'0L&�PF�a���������#��=8U�Z�YRYU0f:/�^W��e'�.��sp�x̦�DR��2J�-�)��[�he�S.�Q�+ҕ���1P��j˕pҪќ��t/I��[Q	)p?��C�Sx����ZX��.�K���Um�n��}(����lݗ�c����N;Y����q��fY:��$M�����F�닽��w�V>l�BU���{�&5���R7��` ��S�tA�0�BQ0�l̹ТR�1��C��$��e�Z@$枫��}�B�0�6)���2�97�#X)�Y9�J_���q�K_Iq�d��WC�jG����6�p��T�8ij���f�L=K9*&�/�g_fl�9�7��1� @a��;�)��]wZ���uZ]����D�F��0XG�x����k�1��W�z��f!l���Ю_~�e��w�C�����+�����y�eF�?t?}���NG�����]�n�h�;�yƵ��=:s�v��]{��G���P�+�B�{�iD��Sf��3�4�	��Kޓ���k����1������S_v���_���^�F ��Ք
ꈷ:?>�d��I�<*���g�����@	�བ�#V@'0p��F1�%@X�Ã���p�j:�Y�z�JX'�B�(�ÈO ���6vq���=C�>�25V�B�R�������_�\W�؍��4�M{���0��tC�G<3�P��R�/::���?�Us��_4{��.g9;tc5ˡ�!�0���h�v�]���E����w_���̪�k�T�N��̌x���{��ߍ������;=	�=�>4�s��HkF��5n���Ƅ��
>�<����Ax�V�.�Ēu/���/�b�����Y�8&e�%8�K+Ktk���:L366רխ��ZDp_x�}I�Ȯv~��Ǟ��Ea��eӡ)>��h@:��rt?���hM�QH9o�l��Q��~��JǹiLƜ:ӟ�gه�6��ձ�2�5�)/���('p~�l� վS�ͩ�g����צ˭��==_���gS�^���3'�T�߰x��q`���,Ƅ���~���ħ>�Z)���\lDR���Q��y�T��Ϥk5��i��;͊�Ms���Y��#rQϓ��w�~:��Y�p����I̸��&�v��ɂ�`ǚ����f�`�k�5��K��1��V@���G\������w̚��@������,��7ݞ��5Mq)_0��af��/>K��g?��7hsu�h�f2�V����	?[�������h�^�n �j�xA`�t��V.=�昚+�B�8�-A ��,�mЛ�q_qF�����[g&Hbr�T��B�^�4Eb"�+�Z�M\�!�C�X`A��u t)��U ۦQa�*C����{(ǁ�����v�e�<4�A��{i������>��<�s�<�k�!�8�-�Ǟ�Cڃ{Ǘ�!�*C���c�¦2�2�X�u]quom�X����o�[� U���A��⹃8#`��K�͉�S��눇��^���2�v�A�����W������l�|Sn@�Q�������Y��oX�5B���뜚f��D�ﳆ�w0L�����Z�!�@W㠴��h��� �Hq��̌
�F�@��-�c����yԜUZ	1ƍ{C�9r���qu/ea41��n�.ް�\�\�X0��X벦`^i&�Ԧ��gϲڴf|6ݛ�a՘���{���D���+k�jV̖
�n��~��Uu_j0��T�]?�F43��F�34F�De��˾,���0�5�X�`�b$9��Ħ�%��-�<+����@"�U8����y�ŖW7�o��aM����iG��(m`�\�܎��GG���pt�
��
��"::��Hlɲiz�P��\J5C�1����H��3t4T���'"~��߳�	+��cWk�o]���'	b*I�^�=�ǖ���}��/^��G��"Ǆu�����h���KcQ_��x�3^��̋�}� �͏��j��}x�U^O���=�Y�Щ��[����J\�	�O?�CJˤ2rk�n6���t��eFUc�7��L����*���?�	��׾F�hL��a��汰�y={���2�OC����a�P�p�&�|�u.�y���4g�}�h�0�CX��b}#.6̛]K��[l��cbm��A\�a����ԧ?�%@a������7�<M׮]?{X�|�!�o> r]"+�/g`(�sx"�ic����q�>#�.��ĭ�O�WX	 .0��1
�dl�%n�8lP��īd����{�>*�9̆�	B#'q��^�2S����Lu..;W5�_� Mv�;��	�8�-�]���V��.V�Ҽ��]Ka��������v�i;��Y��O���v��d��8�u�ǧ&ijs�	�^���L�a�k�i��W1�aD��|��2cmФ����n�*��\Jl �E~s��k$��;�}2���������Ad8�ܾd,!{��E�R_Y�T�^(Sv��x�3ߊ/�䗉Ԓ��^�M����
����93�O慚�B��e��F�ǚP�d����vHt Z8�읋��������?����S�8B{�{�G"c���֏�B�+Oi��u{�ӟ�3��G?���ڿg�z�A��!��˄�Hjaw��0��;�q3�O�s�\j�TN�>M?�я��G�~F��zk���Ao,�䒤����d��9��1Mo��(XS%~����U��w������9A�V͜K�6 2���4UM�
��Io�x�w:����L���)��h�Z�B�7qz��-�,���E���"�)m�3� }���t6ے���S�&9�k�5o-��H���bZ�c��8b��lC�����z�X]�4���������~��Ǟ�����_�\�be���c-�B���ڂ8�$��/Z����x���Z[yCVmP_PM��joڿJ�]�1Q@��aC�ehUq_�Z�hB*�L҂&�k�QP��WkIÚ��ru~������73bn�V{�[����[�3���o�9� ��GE�IE�g�s#�?�s�A4�l t��X�}}^/]�D�����?��=��N�8�DN�}7�Z ��<��T��{1�P�_}�a�L���^bfu��a:z�?~�����f�0�+R�z��?�aʉ���5↛�.ɘ��ﾛ50wX�-g��=�;vSq$�D�s
�����'i���o��� ����k�Z� {a0�vʀ1z�
�����3���s���'[<|]��m�dE���q�fz�5U�)���¸tlR@E��ĵ��vR@����묗3o��Ky�~����tϻ�w���9�Q�_�}�A�z��z���@c���2�3�]�~G�Ǟ��A�e"��f�P@[@�a�ц����bЌ9"���!G1���1��`��؊�IwyZ�����}�<��W?1���R�����M�y�0���n�QF.��ߡ�5��^a�Ώ-�[�lP��T[+B������ǉY���y<��1᱄���"?wD�wlIK���No��3|�t�������c4>6F���]�rՕ�:� hr�0�#�Ȅ�K7he��D�G�ێ�fyHy��ANM�o-��hf�sff�٤��	NQR�=�fy\S�WmПK�
���zb�-W�#bf���`M�o�����ZvT�L�, ���/���W(�͘S��N{� ?m>@}`Mjd�%p��M�g]~���է[�����j֏��ms���������~ApTw�`��y*v��A[��RyV�I 9��BH�([�x�&x�����޷��m�u!�R7L_��<�-�{����|{�B�o���+��s�:]���EWs����(q@����H-�ݶC�Y�.�|�9�Rq�]�D�p����5�y��_�JћU&�*����$�5^-k��c̣AMU%=���ߍk��_�|f�V�l���Sv�5uM|Q8f���L0�E���W���� j\���ss�����Jt���+v:�=4�����3�<Â�ɓ'��'��'�x���>�1�{�}|��>K��կ؟�k¼�uĸ�0�Hգ�t'��������CebZ�q��4����a���'AkL�{R�?��azjZ� +��U?~j-�`�@S�Y�s��ԏ������L�����,���[q��5�L�nМXQDKǳ���1�7��8���� ���?I&	[� �b���9��V�uI&)��?˪��i�3��(
��Eȹqc����[k�eFև��y�� s��w>����R�=��]EF�YYW���1�ʈ���ge�]֩\_G��g�"����li��@�z����fw��j{�nV`_�<e���)yo�\��a]�G�����&r��,X���cQ�I6���[5�aLܗ��k�Z��&�Ժ�83��!F+"l�bF���+�>�ٺ��_���Ȍ�L6�i5sD�y�Ɠ	����^�L�A/���5Z�X �4G�ɾhrW��a���w+��tn��8�w��s���iY�@P�Z�cL<����fr�˿��/�7����C�p��7ܠɃ��D�htD��3P� 4��.-�F��<.��F�Ӣ�LJp�䏈k�&r:�}�L���⺋�k�һX�x�����Ao��&��<� ��:k��f���b�gΜa�s���
��"	$�8����3�tk>r��Ta=K��Tކ��*�Jٵ���зOtߩ0���7��MNY���{B�k�ޠ������<k��y���Y�����u�=���b�ܥ[79f��:ׅ#���8N_���S�9A/��:����Z���~�{�:x`�MO�e'6�C��+�Ӎk7�_?'q
FH@�@�h�:��@��ڕ2"j�AYy��<ֺ� Fcc��(��5�+�Q�ؼxL*¼8�_���k?ǎg�VSbT2�n'r�8�R(��m��w�y�z����������3VXKR�g6��Gt'4u4�I��զ
9�K�汖�Pw��ӝ�I��a�]E�i6�Xs\��;}&i����T\�����fb������7A�+�N-���̬�~�s�F݃�/����I 3Y��p�O3��P�Ax����� ����
)(�g�gֽ�����򗿤_����4��GӴH\Ly�5k`b�V�A�o'_�kh�}#UN-�f̱�o���3,����l���x0s���A����~5B�Hۚo5���{��׋��,���
n��E�ˊ��ʭj-�:N���6��9���������8xQ6앍v��y�a3'�t�������t��%>��ɻ�;��S�D������������ӧFk�C4?;NO=���������?����Kz���O��O��c,t� �t>>bL�O�ᬟ�����w��~���3s�4�q�7m�{"�����������{�V�o��~j�Z[�?_HR�s:�b(�����x��Uy�C�s���N��=C7�h�a��F���js?��Ӫ��Qe*�\���Ç�Ѻڱф�����(J���0f9L���*Jb.�8��06SЦ!\5�h#V�y㜩i�	� �"h�sY@���#�����kk�l���V<!���=�='�C'r�@��	4[�u^d�+�dj��3�}�0wB����N���o���bMZ*��Z�5�j��`�_}��%��e[eJ����e?4��2!t
����ե��p� ��zY��4%0u�[���.��wh�P��;�6����<�a�0+�ZS�f��{��� ��]�L�����2� ��5^�������Z�ܤ2.f���)�y����|��?`��ꊋU�s̾��2���K���l����`��i��=��'�ə:����7��;�����Y�l��F(��I�o�'��f.�ON3�@F# pf@l�����5����o۬�>��?���غf�I�ARL�9�2���ya��Jfþ��,@`��f��w���3f��',���J�~t%&����]Y��<��H�-���0�M�����N��=C7�9Y��fd�d,jl$Deb=��#��jG�=
s�UЗr�<ZYC��8�VŬ���hey��n0D��z������{&e�P޿��؆	�^�d/���dV��Ә�B+VZ���Ō[����{�58�IW������gSf-fMvm��s<)�j
�*Aʤ0�Xj"�xѺݎ��e*|AVM������Z��
����f�0�e�9ZS���[<v���q�| c�x�:�}`�ul�s:L�<����!�qc��cf����m�Y ���Ah@&c2A!ձ����㷫�Tj�Ukr�����[����}�I��7�f��hw���-'c(�3O�ufZ_���"s��Y�������s�>x?}�[���6��^��:\aFP@ -[06%s��i���`3]@vD@$,j�h�+��	mf]�����6-.��u֏nW�t/E{k�
�X݊�uK�Е�;G ��J�2���X�#k׿>��~b� ���=*{-)���4�5ҳ�+ �{������=COŉ��,1[W���|�f�Qh��Y��P���\P�rA��T��i(ڪ|��iz��S.VS��$� �MY���%g�Z9��T�rc�1k�$�ǆ^����֊Fi=�i&�Zڲ0�2�c���[2Fi�HԄ���� ��X��oB?�o���؀+&l`�#��u��'yV�
Ʃf!��q�@���!�K+�A[B^�f�7`�)�W*���W��W���@$cB��v�����6�������> ������B�z�ag�a���8���� ���ò)�c�)j��s� ��c�*8��/��]1: ncw{��b�e��<f���rX����_|�E��Ț:�cܤO~���+_}�h��97�{��r�FDc�3�٪q,r����{����6��"){b^�9��T���t���7�=G�<�+f�Wd�����}��f�p�˽��O_��W�g����dOd4,�ObRh,��t�eȪ�J
k�Yb2�j���jU`�2�~��(�M��l�5�E�V7�_���y)y�7��.x���C�펴�=C���?zY{� ,zSM����0��U��ŋS�"*������ϣ�����L%-9cmI�"*p�nJ?g�|� P���B���ܷ� ?�Nϥ���3�Ի�c��|8���-)fUn
�ܲ��d.�GM�vl �=C�� a�y����5~�0w����_��G�� ��!�q��a=!Z��k��6�
�8_PcB�r����>�cAX!$�=��l��U	� �	�fƆ���/�:��u��3�f��Z��G#k�5e^���5����Te|TXO����	��Wc��?��]���*䩺O ��a&�
 ����z�W%�XQ�ξ}��̳���O�{l��aR�l�&�1��3����jN�׿�uz��w�/��������pMT��5n�3�v6��7�1c��Ɓ��i������i��~�>ۈ���l�>��s< �b-[e������� �?��ͷW�]-�x�*~�@X�#�帜��~��XrQr�Z��5����H��3�'N�7o��E���ڪ2��{xan^X��B�pĩk�6��F���)�MSy���`!i�����[xI�VW3�F�&I�1t_���H
2����z�0HRm)�Ǔl���o~� ��|| �QtZ��9��V��؊��M��.z^��S	4��b�����I-|����ij|�}�g�:;�/}�t�0u<�K���7�ԩS|Tr;|�C���ҍ���~0�WH��tce���w��[GHR#���O�k^�q&=ӥ����>�Y��#�O�*s-w���Y�l鱖"}!
߭�P*셌S���#L�T�N]$U��{m�|l�3h�=�I¥����
A������/9ƴ�H-jw{���~�N��:�۷�Μ~��6���i�qo��U��[�����o��7:�ګ/�u�����z�uu?s���&�{�M�d}V._��c�����Ϲ���ڌ���gf�[�;)� 4�n�Ҽ�
��e��)"k��Y��4�Cj�Լs����x��TAO�T�@�yV��1s��E�}3i�D �.�G�>���Z°��#�V�
rPS[m���`sno[|M�.�?y�\C�H�9z[�nݼ�o�p�	���ZX�q4��V�:X�E}R(���v��j0'��B�)��w�Jݍ#�p�G�Y�z͎=
j����[��-���m�y�<o����\��7�\o\��ǀ�!lҖQU�3�+�'os3�={�G;/�\t� 	�
L�/_�0�FC߽@.��� M5I���oX!��A�Y $�3
�UR���uϚ�g?�C�c����rF(]_]���q~�o�9-eB�y� 4Mz��9�Q��P�c����0�F�����ү�o���.T�rP!*�k)'�YRCA�{/�_pu4�M���Tn��G3'7o���25�-kM����f])Yh֊�ڒ���%�8θ��>k�Ȋ������tk�]C?����Ɩ���1V�77ש�6�1E!%3���al��Wg��/Ѿ�Mߑ+����8P���Ȃ"�LY�P�k,]�a�i�h{.s�5�~�5j�q:E��7Q r 4*��X �C�#q�V�4�<0bub���{�4�A�������������Ѝ�h�W���F�jWfas&|^��,�^R4A�|���M�1;�4��� D�+hML�;+���T�-#ȕ���v��ncc���8�|?E�>Z�n�%�����f�4�5P7�f�a��(l�U-����t��@�#�X8B�{RM����`�H�	�=bBb҃I��]c[��θ����􌅝HH.jᐳ�t(���}��P�ZU�iH�̱ȣ�0�ƴ��AKK7y�'���ב��Y�m�*0kC�m�czf�0�c���0�� }꓿��gk�P��|�h|�{�0��0$*"ջ=�Ŵ-c1�)Q1֎�c�)����3����P�cz�j���K�����P ���w�����~�N�8�Dל���b.���-c4Rh��:�&����<m�V�\�G���P[[�V����ތ.�ϏAC�f5�"���@s�C[y��se3��9�@����۰�a15�3__[�g�a�3�z����_��f�<o�a �X�q��,����F��7C6�MZYޤKW��}�ZGf��z���r�^��s������WJӚ���9Q"�o�:��������a��M�6���0$��1���u�Z���d(ȓ1�dF�q�C8�;~����Ǒr\4�>0�EJ�6"�d�jE�*UI��+3ys|������a��R�E`��Y$=�T��Z�D.�J���[�� �t�1�L4�a�Q�tܵ`aA*v#�a�s��^��Q>a�뚟z�3��=C77�������2)��|w�5s���*]�y��C��� ����g·���8�ת}!��g�
ʀ��c�k�fת{�N�U��S�l�͌sf��>�.]�M�����R]�0aE��<� �P+��IW�. �@����GCHkB��A:r�k�Y����� ���g4 ��o��~��|�G7���\8�5�X+X�c��d��>w�vJ`Z������1�l{:x� =���L�q�kRfwv~Gp�ٷW�#~r,�b��>���q�����Y���9g��D4<~Fa�J��4�����YFe�_Nu��y#���8��J&~[ �ll$l�v(w(�Z�������ҧ��� �ӆa�s�E�I��^�r��Iʕ0بOHU�3g������g�[F���W��%�o1-�PP���������y^u�h�Q��9��\k(�a�]�ȭ5�V�kotC��n�wZ��pf뭗������My���`Ծո���V���{J�~58�iݖ�1t�;R�4_��˷��8��m搥W��G°�7���5#��al>7�ݠ�I½�-��V�)��l��GtQ�������4�v��^�1J� �Y5�����a	(�>�Q��MS|N�4�� 5c������ ˢ@�Qa��>!�(� �oaA�|�����7�T3s�גw�s��e⅓*��ͱ�=���,�.,\[6�^8w��F�<}���W�m��~�:Z��0
�2��	�(&�Z,6�:6�H�Sn��l�ٸL��Ĳ�5�L�vQ]σPͰ���Mr=���6we� �a�#F�id;3ʨ�g���"̅6��ۍ���y��.�=��	&ZN�B����j��`�^]7���<~���½�Ɍs|��e�Z�] (�Xᔷ7X�?}�M�H���$9�[)|g1~ �(^3k�[��d�#�y_1����6iߡ��c������]���9�Q�`abzv���!(˨���x�n�,Qs�ſ��?k�y1F�ft��FX11�$� �}���B�fסAi�{X����A�)k�/�%YR`z�D`��.^8O=� �I~V�FpA�����|�3��sX�qv�k��Nǎ�O>� �FE�!�ܧf�Hn���`bk����"f� �R��K��
ݝ.�Q����<_?b.(�́�^�)�8��$ʱ��
�yYaŷ�7���#N��E���@�B���
��C\_	MM	4/�5��왇�:}�ߎ������g���\�[�Ʒj4�L��TщY������;*s���,��z`i{�8��E�=a��lU�W��`�!L�&O�#&�����O-�rY$���/|εr|=���g�J$R�ͳ���~�w�L�3���9��V{nG0t��a�KZ�v���|�t)�"����)碗�����#�c҈{�Lj }P_����k��J����ݦ�-%�غ�J��=՚8�'�U
/U�z�1
Q��Ȩ9��?�'Ie��R����%-3zQM�ȡ�th�v��߽��P���̑�3��,�|P*�����g���i&���`�ow�/��4�O�&��{������K��AaPA��lL� �4��9jf����Y��U_��[K,"�y������כx��{��
��6v-B�9�#���Cȑ�:�i(��^�Þ��ُ��
g�tzle-�0�ccW���
\+�Ξ=� :Ms��s7�}�}ToM��3G���/�,����?|h�w� ��ޢ�ﾗs�	�p�k���q��yTl��zƸ�>��0=6��9�Ef�J�jL��B٭�Įk��Z�8�5������j�c/�a����=�ٿ��.���;�ē �R3�T�P�6?�B]Pa��.A��}��� ��T˚��f�[>M)Җb��0���R���x�T~���v����-b�g��NYJӡ���ڧ~���-so@�:l>O����q��8�C��#z&�YYSS�P[�Qӑ?��Pɺ�y�7OU��,�t�|MyСպ��"��u�E��^_�_@�S���/d�}p�xj���Nt�0�T��V���������E�n+V�J�s�s�j?y�h%e[����8���	f���'鳟��۳�������@����F�4�� ���;�������&	V{b��n����h�R�J�M�f�\D�",�A��w8`s����W���'C@Y]�2���Ij ׄ��P�;��ި7>9ɹ�+�K�1p�h����DIc-�鰏7�2�q_�-�j�������o��i>��S. ��~g���A��4���U�m +,w;J��O�z��r�,\`l�����A��?���t��~:<�3| 	��:M&w���p6L�$Td���6�'��[��ʌ����3�s|o�v����8�̫3�����p��=!t�2�,Gh��$hzI�q+s/��h̲�@݊��疫)��}W ��7�S��kjpq�����o�/�y�JS$�;�S�����ʮ�T���{���ہT3\w�%�Y���|�̬}F��?F��޿>/�n� d�fn���h��:��O�}mY9�0��Gx��[���aBB�����K\ڿ���P-.�CO+�Y�n�@5`�8�l�Po�?�a��ΚZ��E%o��ˀ6����[Xd��m�h��x���Uߣ�xI��f[R�j��0f��'�6v�0�>�����=0tA�<+*����m0�%�<d�c�#���u����}���RC<R͜�gV<3�`��I���	�
�o��L�,h���6���&���$�͢`"�k�X�� ��	�܁]�Yw����6e���9�k�_�ϙ#ăχ�%���5����Q(�5H��˳�0_#h�5֢cG����G������,G��}�挊r`��i���j�x����}S-��>g��0ڄ�^�V��MԘ����s�����������f����!t����,u���J�W3Pxn|tE�ɲU�����Ӭ��+���2i���u�Q��ܰfuF��A`��fˑ5�����j*?Se�>�,�4�!�n��ǔ߫��ߔ�Ӛ��C���6��(Ac+�A�������H����Qx�ʕ-�vC��(<:䡖[yQ���5�7X�U������v���}W4���h�`e��M-���j�I?qhS�A뱛��td�I��S��"���hĔ�߻u�Qq�F<CkRي��a����;��1��^7��W���ش�Z�;��ݞ�G��W��{=�h�i�459mΟ�f�ť6a��+Ŷ�r��C]J̑Y Q��|N!S�DҴ7̺��z�׬��>5n�Ā�	��� <��u�l:Wa�tfB Z�`b���-3�]7�-�!{�
���G|R�����,DxO(w/ca�&sߍ"���Qf雂O�!�D���E�����i����< �������+���?�˙���8��?x���}�[�c|\2�-��$��\�ҥ��x��~�تk��/�Y��ΰuc~~?5�u��#п��B�O?l.�A{f������^i��
��l'���+ps�Q�v�sCt�L=��f(m� ��8-̃Wl��X���	2,�'���|�v���J�̭�oYO����*��T�t�����nY�e-�j��vA����ӷ|��Ͼ�V%�H��`l�^���	���Ҫ����#z"X�i��Ѷ��J~'=_�QI��f&�X�����U�s�%2�@U�JB�����v44��U��AP�[Y���˟�|�VY�?6�'g�UrU����"m�9���d-R�@@�NR-io x��i�k4�~�� '���
����g"�L�h�@[��S!0P1��4>B4ƌ0��|!�KX��a0u��gs�A�e4�"����F��֖WTg��4��rs�^�[j�YC��13�^�Z�S4b���1L��5cH��tO��cL�p�B��s�ϡϰ��~jf��8�=���u5�x̳	)%a���^��ù����!���Gf�) x�u3/F(ZZߤ����7�2�X��Vu�a��E*�ӫ��JǏ�=���ך-Έ�=�s! �,�2��˿���>C�����.���o$�u�)]�z��>s�7�;E�D8 ,��̴�	�a10����{T��fС�YW���(�HSy���g�L�l��ǛӁ*Kg�ҁ�
��~�/��QZz�w�U�@�4Ϳ>��t�I� Q5e��	���Ϭ�n'��_5߼j>wi��#�Y�YU�?`�J��	͏X�����I{��3J����1�|���h�e5�"�e>��)��{,/5=�V\�N͘����.Ei$t�T����LvZ+[�k`}S�>�t3��M�n�9��,�hm\t�ٰ9�5�����a���n,\���A�Q�L{lR|�3�3\c�m����o��rrr��,�-�fw��@k;z�h�HaB����kL�S���,<n����c-� 6����W����n���5:h��t�A�6WC�	��e�0��9��5N'N��&g�=6Z`G�5��ъ��%Z�S��c$ ��1���h�0�F�Z�溵X֛�r}ޡ� kq�}���(˘�s�J~����PL��^����
�Ħ�����n/�?��k�����4`��7��R�0C8{�ԛ������t�>��#G�ȂY2Ө�Lb��]w�M���Ϛy����f�3�����5ͳ@�Uh�͸EY7c��Z<�� Ը�����?�'jo�q�&r��kG� \q������������b�n� pi��ǲ�׷@a_�����Y�C�UT����p-e��ˤ2�J�[SW0K\}��Z)���Ԩ+�w��*�}X�]��4�w/Ҡ@QŰ�j~~��6��	`Vi���ǆ���N�;���7��'1�߆�X�趣)ng�(��&��͎lRP�c*�珋�@�]8�K�h6��Z����&CW��~b��i�w�彤���*$��}>;	�8�I&�3H'b�l�/h�@A���'/6�Ti�R���MN�$-��r�@�#R��۴t�0ҕeZjM���-�2"�E҈hc=5{Q��FV3�+O��]	����d}��`	�Q��L4V�N�����]Z\��~�����V�E	R�)Z�vC�ͺj4�n������3�9�6�&jT�nˬ���@#���(>�I���@4��d}Αդ�:�h$ԯ�z��ֽ��4(e漎j��G�@��V �瞣�=��������2�nh�1}�e��}�����~�kz���Zcn�,�!.������]sN�L�o��o����>i4�.]�|��~[[�`+MB"X& �I5EQ�8��/�@?������>�EYj,��o4����$0�!�6�ꞗ��g��	�( �����	E�ʖ�5T���
���Yhj���3}�����9�tmT�;F�#����*uB=?�t4����2���L�����%����Q��^�jeMW�#������ɢ}e�K������W�|�5t�c�_3��0=����33s��3��H�h;��#�S�S�)%���1.�AS�������Z1�ڠ>xI'IЃ0u	�)/f7��*�D�^z���Zω'���4 ��no��
@8V�y����v��I����4,?�c�p���o��l^s}�L�~.`N�x�ƒ!�������y��*�Vs��O��>"a��l�np[���\R��@~t�3�sw���a�Ք&&x�	�X��r�u�L@�#���q%�L�^#Fݲ���1P� �5cZI:ԭMg�n4}3�fD�;�@��I�J�
Z�����^�'�i1Ji�|ي��m������ ���l��B]�*s	��aRf&n�1�¦�"Y%�Zh��d4FK���q��2�ڔ�$O3�>�i���\��$�NM��d��Я]�J�.^���~Bg�9/ ;��s�}�����:y���)�x��}�nh�+#0�d <��V9>�W��-\]�s�s��o_��1���i�~kZ���b-�3�t�ez����g��k7r?4�F� E1Tn& 4�v>o,,i��!� ����Z�4��f�ϐ�h��7�i!�֪��&������i-�~����-��� Q��LЅ��S�)�V��3M����l��2ì����2@j���AS���XB�hʌ�5���,$�,���9 ��L$��
�Ԏ9����ዃ�0����7�w�q�n���f����`����Am��Aǻ��?��vm;����wO�lb	�Z��m0c���+3���ޯ24���t6�>W�����,����ܗ/mC����;8�f}�Ξ>ÌG��t%�z��cQ�1���G�����V�wo֛��$2n%�l�%�3��{ts}�V�QP�M���2��̻-_:;m���<��p�c���� �.
�t�0�`4��t��;F�[�~o�`䧒��i/͋�)��r/>A����՚����W�i�u3���]�����w�eE����u3�s$�h��p�l��-� J@���7�}D	]�z���p0�e\��၃��|ݩ���A*���Μ���A�*�h���q�̮��LB�R9'�$� ��!���a��W_���e�-�s�5��� ������
-,� ���B����ߥ��y�rլ�;��rP�2��9~�7/����p�"�Y D�w�<����j�pW�N Z��L׮^�[˷�	A�& 5�662�z��5#����6�Yt�T�֊@��{��M<O-����Z����K��3�$Y!B��r�N9HΧKL�(�z�d~W���̳��̙�L _x�qc�Ln��%�'k�0p�ی���g�7��g��4�l��L5?������x��30��ŵj�9׈c�YG��f�g"��=L�l]7L9�~�5࿥��(��������Y��~6��7󐌏g��=�߭I=3{$=r�
[�m�vC���&�Mn�XG����(��0�J���9Y`FȏW ��5S�t�4�PQ0��T�X��\��,�w�0Yk4����+�Ы/��n.�`-AP-�L��h-���,�??o%^����s��T��}��Uz�ۻG��$sZ �����!n������i�hϽ�����W��`�e�303 |N��E� �YfY5�p��^{��݀�!�/X�"`Č������Т��n#�`mĵG�.yԜFsq��V��xkq�fH��7W�hl�0H�k��zB��NDH"V��9~�֌�ُ�����d�L	"')r0yc]�:f�g��׿vK���bZ����w}.�����5�%_�°�3~�̜����;���i}�i Z7�91��oF��>rԗ�hqa�:Й�1�0�T������i�_�X� hX�kf_y�e��$:�,O)3}`��d�f� 
�="T����>�x�Hj9��O��&�[�2[�8��C!I�AϬ�e�~67����q`�/��y���n1Z6��8N�D긔ɗm�s�.=��invϟ5��Oa80�!�d̜c�#b~f��$Y6_�A�FQ�3̸�$50�Ԍ'��llq\	D���A&��u�<x�7}�u�R����#��*�� ������*�]��?��=G�+���BC������U�Q��Sgv�th믽��������stwY2W����rߺ�So������9ʉ����xL�"�E��i���jfJ�F;k#�E2(f��i����4�TC�'��T˛
e�!NAc� �J�63e tML�����B6�+t�����C�����7Ys�����*SSF�5 �.�$�ה*��ח�͍� �����;t�6W�(���0�p"攳��A�4.�-��1����/Fd��F��/��%�E;v���{��-�Z�w�>�!���oeaAsB�WB�����>6xj������&�c
����ݎM��PI�G��m�l�!hJ� \'i&f�$���0ھ9����f$`���%�g�[��&�6�>�V+�E�k E�BFӓ��В�����)��|_e��%��Eh���z��L���{�<lG^�/��5�kN��T+W�6��&�祫K�g�~�������\��s�4�����9|��8�fq�����a��������������s����k��9�P�����JZ��$���iի��z=/��%F^���,�M�����ν�6���~*�g䥊hk$� Ӡ��G9�P�"�y����,j������Y�%�9\.���!�k���P��g8jj�R�ݧ�=b�c��D`MM?ukr��c""��hX}��(� ǲ����0�F�M��2hǕ�l�E���ベ���o��e��5����U3��ןҥ�����5��z��O�Б�yZ3l:�4��n�DTekd5v� ������y�k�P��A6�-Rӌ��������瞣f=�hhhTo�9K/>���׹��k�����7|���������E�tm�	�6�F��7��[M6K����hɾ���Hj���wb�V����fr�r��	�' �j6��������!�iP�2҄�f��y�r/�  ����صA�`��c���/�L�%P)�B*󙰺��f�4�U�!W�:UF��?�|CGV�l��~���MMO�1�]�e�}�!=o���Xg�v[�Д�֫d��yf}]ef��ڋ�w\��2��c0����3��gӯ�+s0]���[��K/��®Q�h�Y���O�x�������fh�,2�5B���"��ރ�n�DM/\�N?��O��O��ѫ��N���O�]���z��4�7ۆyil��T̡<�ʐ2{Y�Ѯ�+����Q3n\g�痿�]��D3��l�8s�v_�E��6�)i��#҅���}�N�z�Z�\���ٷYk�\[z�9A�IH�NB�f)3�ӌ�l�n<
� 5k��X5���_�4�i�9(��1B��NJ��'�R-�y������LNqJ��N����:Ò����~vP������k�~�2�*]�hcͻYbi���!�y?&����2E3��y��y�F�6;��D5:3����;c��8���HR�l�RE�C��[����x&�'N&RfA�
�j��ْ�QMJ!�Ń�Ɛ���Б��@1֭7��X�����Ij6bl̙:��"���yg�Ih�м=姟��J�f�f�%`.U`��$��V5 �߫�,r�Wu:�y�1|i5�w�G�vC��1I���!�����3|}��}F짎��O���o;R`��0���=,��k��3@�9��A�K�����r�N{}G Y��l_�F����1�W��i�g0�0�0-�d�x�Ka�D�/�O�S���}@������A�P���#E��6��`�36��_�Hy���;(Z08�=���m��믞�3o�������aRMf�l"��nƙ��J�_��H,X�k��JC�C
bh� }�F��5O��8�>�(J��_�q38�W��iM��7�mI]
��� �� >r��%����gfiρ�,� �-6�h�|��Z@4Iv\�K��#4�6�P�����p�㐺�Mj y�4�'���$us�µ��̍.��l���Y��9�xLO�o�ײ<�Y�9�N��j���+cW_�j�h�l�X��H�x��1}|ad`�0�#"�fR�K�@Z \$q��]�C��g,�%v�����=f�H+��6���0����G�C�J+�p�����9؈��g
�a� s��B%hM�	R���<����[L~fz�sn\c�,Ա�0�1��
��B</��4ɜ`﬌�<pQ#[f:+�x�}�� \��YQl�ub�����&�[�YŃ��v�u@�O�u��߿��߁�#�����'@*��Z���G���9�5�� �#�3����B8��h@ c�V�Uб1<��}�Vdc�(k�6'X���ėXb����k%�Ԯ�T��������f���h�)P��0�AX��U͓���S�2����&����cC��߸ef��G����x�-��y�{Y���5"|��-��֨q�!�m���ܩ��ϋ����V��_�@ � xж�׻�+ B�X�I��4����Ђr��/�UZ�p�&����w3xX@���T��%k��4��` �!��rHL�<~ʍ��=F���$��_��_�U�WfY`,&��M��[o2�x��~��+;�t�iԻ.��|[�=H��G����}�����oj��󱖱�P�>|�~��Q�ʗ�K���O�WR�Mn��9g�Fߚ�<�Ua�qZ:�;A[]lJ{��쩃������Ӝ�~�[��X�N�H�K�o� �`�����mX�1}�.��n>1R�C *�+���c-��������H`�`Z�Q��=u���Z�c�K���<��K��-4!R��Ƞq�8rI���a`7z��-yלHˌ�mk^�U������'Dy�.��A�Wv5����"��^�:������P�Q-B�)���y,Ʒ��YF�K8�2�e�Z=�5aS{���|���􄙿4g��l܄�<���6Z�E</"f�h��x����V \ő��ͨvf�!�I�Y\�F�� �����թ��i L��rAc��%�, HW4L�
�zN^�������^��o��^6��߫���vw�mD��07�v����Z�����Q�1���x
�U��[�<g����}\�uy�cC��
bk#�t�g���5�Ot�Q����"`�i�Y`���b� ����O|���u���}�Y����h�ݬ+�%6C#�ض��I��vGڎa��i�{XG�7ٱL��(��_��|�������ƅ����B��y=hFC���O�Q�&�����HY����Dc�m5M��j ��3��|�Vmb3/@S��EAs��������-�(�W?@Q�.��D�O`���P7�	k�5���d�)yY+���F��0�5�-{d�|��F3'��?�R�z6�s�3�>���m�BJ44���I��u�����;��kq��	����3��;�/�"��|?�Z��L��Q�~��u�� �]��� )j΁2����ˀ1I*���������GD��ru�r��v�����c��@��"@�UM�zE�ca���ƅU��{NR�'�Sl�!	LU��G;�i����\9���=QaLnm`-�M������EkƧ&�����e�0�؟����T�ݶ���z��ާ0��T	�03z���wJ���|l����5~�x�:H�s�_��������6�η�Ea�]n����3>9a�+LM̲9Qe��]S"�5��aA<�Q�:]����8��0Ł�t��<g1i�wƪV�D���M���n�<� *d��\�'u��F���5��F����~�=/�KUR��w|+H�Igj!�������'NL��Z@WV�Fd�+� ��;y��H���֌!n�����6 � ��c�ˀ�uc�&m�y��-Ğ�2��l���H*S0�3�s2A��u� B����X�`7Q���98��
`z=?�N׉̽��ɋ�����}��oe��_|�0:���[<.+}W�d�� ��/�6-�sz��9xA��;\��mgib��Φ���χ�01��$v�z<���JbO�����}�1*�z���9CO%�����Y ^Z\f!���y^�@�g"�z������Э}�J~��?h��]�O�6uIj/o��D|}$-���4���g�#�-��w�u_���wT��9`,��E$pn���h�D�)�r�]f��HmdX��ɓ'���{������Ƴ����!8~���ۿ�͌S��𣏸k�޺�=�P�艅�u�:27�|&~�u�/�<��ۼo_�W_{��g��D1�2ڋ�IJB	��qpғZ&9�Iʦ��S(�	���_ä�W��a�Xp6y>0��`M�0�
θ�b��� F�m��G��������ܹ󬕣vv��pk��Z=̅;AX 5�й6���,���11n����f<c��ZY.�ʎ�fEᴌ5�f� �s��"��&���~��a´���ZŚ)[�F1u�}X��b�o9F�����5�LpdXk|F��m��
T
0c��C.�����8��ji����6�l���zA�zϬ�s��х��!x�����غ��/k�r��v|��o;���WX ��W�
9����'P�뗏�[y�?����&[k�~�cǎ��`�O:36-�5�0vD�������g������y��1?b�
���|�	���<3)���~ |�sO����q���rH���q�WA��.�8_�ڰg�����B��O?M��ַ���t�������A?��_�f�͘�'ǘPe5���֕B5�Bj��

lf 4��9�h����n��ps��Ɛ��$pm}S�U�C[}��#��й�?�q��w�C��S\pdem����.W[��@��Gh���r=Y�uɑU�F1��5�� D3�$+~u?S��KD�9�о�E����[�D0A�23�HP�PPF��O��OO���RK�2r����, ��y��\e�Eƪ/��i�<�R��Rs�<�>f��<���<�!`��& L�=�[�`v��B�W?a�QXd�:e�|oj1q��@򞅪�z��@F��L�A��1I��'s���u7 ����E���$��E_&RUǎ*|S~�V�L�0�;�F
�Q�,���]�9�Q�ѱL�4�+ް5�%T�޵|+6(��~����q� �A��/ T��h���[-wO�ׅ�:�h�~*~u5��jF	fJ�� �?�8�8q��6���Nҗ��yz��_�����is����$�)&�r���?"���Ιu`lH�
�/ЧF�f�c��]_|�66;|�C=D�=�8]]�A�y�ejwz��&��;3�j�z��>��/�uEQ����p���fx�b9h����e�vn�.�,EB5�šY�@���0���>^}�5z����7�.̟�i
%����	��`u.�1�z`]���P�}��h���$ר>fԾ-�j�����?��/Xf �([elj[\�2t�gf�0w��G�EC��\��M�P.�n�,�;ڄs:m�~� ��g�����S�1�ۏ0��7�M��T�=b\�B�_��G����&o�z�	#�m,���JH��O�T�0W�.�<c\Y܃����*�M6�,�fU�=޵h�2r%6����v�j�" &6��<��ɘUf�i#�y�-aJi���ϡ@k
S�`"%�GG����(�s
�ܞ9�e�����n�� :,I%X-4s�٧�� h�d��E���V7��q
\��������.w�0�?�w��~��; ��d�r95���3��#ꏄ����ξMi�����M�`ƜA����{m�z�Q�l�b�#�{�j}m���n�_�Ϳa�. ���o���ԩS�j4�f�%Ȭ��R�Y�R��U�kvB KLbL9�B�j�~�ɪ�^Y���W��Aט|՞.|��ΰ���[8����و�4�W}/b�LM�az�r��G.��t	���f�ԑ�����[�s�82k5�}�`�%�!��r��X"h�w��>ڶ#�H�`��(Z�?w����Ze��m�� �O~�	�fV���K5t��xEW�<z]|ǂB���j	�?:�4p�+q�-����>pM��F��}�,�{Ncx4@ΛΪ��"��������IQ%w���c�h�V���1�#HT9H�|V&���`�;нp��[k�-_��͔�W6�m���|����?�'�x�&�'QK�F�~�/��$�?�y�c�\i����y����5��1IRS�2+$ZO�^7V���d簹�a��}��df�),�>�(=�䓴���y軖̓�:�/w��)6��Yq��]f���4~�~������j��/�Q4w]ʪ�9���U��A�Q�`��6�J�(?���m���Z��8岘>�`J�'�6l�W5,f��kH�����-��,C����/�?-)�*5z�}�kkb޶~v|F�2�f����֤�©pa�0��bԜu�(SGt������ɢ�:_�^¨�:��o'�6�<��W��t��?R&�(&Է��t�)���4�q��%�7�kRm-���Q�H�~�,iS�h��3{��7��2��4�8�y�� � �5>'>T}�hΒ⭛о4��E.����!�qR�V'i�5�8��0]}Vx	�w�����g�=��#To���i����z�az�����Ɔ�͔\$7
� }M�GvQW����Ԯk�O���|�?����[Yy����
��=�ޫ|�dt{�_k��R&�k�zm��$� �?�sFy�7�J�e_��F�����3r��R�7�G- �֚P��P����@�U3�߹���2���0�P�����+�S�w�0u��k�����NΑ~�B��'�4���1ٴ�����n��14r��K �<
�׊�������Rt8�$(1S��(�(MpI#��%n��a����!�!Î�47{���9f��a�DK7op< ��A8± ���^�ak1N���6��L�1�����1KlrW�ŹF�����ϥY�Ĺ���G{�}���,��"P��_��g$8w�� g.4�bªL�W�!��CE5�߭��<V-�#` )� @�!h��B�Z����ł��6^G�8+R���6}F�Q���V%�o����d4��J��2��z���a�+
�Z������,|�3�m6���m��4������Y�Z�(qw���.����O�V6�%�`��>e�����WZr����2�LҒԏ�LO�8�*`�gן[4M�{큱3q���ns�-q�>��� ��Zm��"�J���L���"��,4���Y�������%��b~P:35Z�J�ڛ7�^C�7�FCL2�������G����1MFW�hxHU��5�a	��`H��B��C��pI-s.��׹y#!�zoN�B��R�7��,h���q.�����I���_)kk,X�{g�ָ��ͺp�ٟ�����r�����g��S�����F���b�������/�Zp�^��c.�rڕ/<W3��>,��-^�:�=�:�e@#�@o����1��IQ��r}j�tc�!�0�s/<�˅NS�,<KhT+X7��Cb�m�ێ`葈�wD���~[��h�Su�Y��-I��{=F��>aR�N��r��a�T��c��P6��M�:6I�k:���?�Lt}�����Z����"��R(b�H4(1cY]]g�F����%0���;���[�k��A{m�~g�����Q���|`����32��k���j�aq=���v������U�o{ߞ�g��y���Ufzr�ſ��{�<!�L}��Бc��7�`���^_P�8���Ȝ�����4�X�Xj�.[q�h����a���41ŏ��?8_�<��;��~h_~�Uǖ�I�cS�����R뷝���WYH�}��߁�#z
l��Ιq
������o+%qK�����+3S�t�����܇\+j�N�M���e��3N�1�/e��H�l�μ�y�a������`(z����'? 2dn5&�1�P�l�M�;��d��3o�F{�R��$��&��azS�!BA\���~�	O�L3@�x�!�L�,>���0"��RȆ5j��kR�A�!8����k�J���[6FA�G������WV�D��g�ͅ�2��U��#��MON���,?l��S~�0w�I�i��ƍszvu]��; B�u�آ%�}��]�t��e�!}�ð���B����JZ�0?��!��[�e�or�kĚ���Q�4��r(�i r���tn��;L�������JE��<c:�v��j;�� پC~�sw��hU�_������t\69�YV�7�6/�U��ɀ����e&3h&���f3�e,>a�Ҕt\>��C}��<��TM��.�_��0I�Yj`�?O��S˅�j�cͭ`�`j��^V ��&����#��tk��iOOJ�J�猂� �iZ��� ���@�<s��:��7�A�7��Ζo-x�L��]�c�C�e�1��	:�Qr����t}��4NLO��b������1�q�Z6��'�&���� 3`��k�R��P#ew[��k�z��}�NPfB�����O׸fa�f�[^��;��g��l'�����N+��o���k�nea@�l�?�~�s��4��h�ro�;��x9Pˈ��q��d���hG=��ֿ�>��3z��HC+�^�7g��E#��r_��aUG��\7o�xe�hy��Q�'������4�v[GJ�4Isߗ�C͡�G��ͭ�LW t�1_�R���~�jA��jZ����m��K~-�AN���
$L#�����,Dۅ��Ao��k�w���㐡]�{C���� ��Y���[���� <�s3�Ġ��i��\/^��i���`%HDK׀30N��{H$ 	jk��HD�St�=���~��݊/�d-H_���u�i����U�	t��}��@c��n���jL��?z�0>|�� ���mx<o�}�������H� ��3��/����e�|�\�߳���&�f8/4��M� :�(���5��Q���ݫ@�"f��L��� c��P����S`���3Ι�B��I��Ã����;��S݊L\��/9���>����>��!�)[3|�U�� @�q���#��R8p��Z��ֆ��`@��x|��n�hێ`�4D�,�܁6L.�W���M�;C��a��I�c��mݪ|�U}�k|��&�/<A!��5���Z�SJKT-W�
��J�s���%����\-q�0/��!��L����<�6��ُ<֨��HEH�B�>|�<��x�U���-�H?����"�l�ևZ ���p��:g��C�p)��ׯ�8��8&��������a�ҟ���J{�(>,�~0t�(���`;4"9�A�Y�WKȕ�<�n*�!�ʥ��I4{��zʨ��aK�"(��f�˃ Ko��%@K:��;e�t3V�e8xn����0�f˖��)0m�~w唊Z�^���1��n�#mG0t���l��D;m{f�a�n�:�d[0'��G��	��^ňo������.��G=��`?د��ʖ����Z 4������e0^��)��XC�҇�O�8�>��{��q��*��n.ܔ6lE��0���5��N��9��5f�/����sL�\(P�YN�R�k1���f$�8�q`A�����˗\���`���(iy��I��S��&��z��ss(.�?�\k�߳��K�s�&��Sj�|?��,b�ާ&v���{��=�m����_��0��{:���{��p��^�B߷���b�ߩ�#z�E�7�]f^4!��.q�b�[��U� ᾿��i�۱�K���L���}_{v���n�^����k���%���<u1�000���Xֹ�ff�F�̮s\OF��4�2a��.�#�u��c��/��n������\DV`p���X���MR������Tk\�[m�X�?Nǎg3:��fRcl��J��Cϲ�3�3�s�83w-�a�C-<>8GJ���dS�Ԍ���Ve��7l/m��>���7�+�t/Tӻa��~��U���Ҋc�U���;�vC3���ѱ#�`��6�ܝV *|_UҾ?���׺������������`3\��H�ٳ~��T#d�4;j����9tlr����1T�#1i�7;|�oQ���*f�;E��4)�h,}i
ƂT6�Ӄ�clHuc�F$��\�~���J��T̽�i9t�5`|�?����ُK�Z+C��9O]��`rg��^ʌ~���x�-�,�!!����<��	[�`�@\?ck��9�[�1h���b����[�%�N�Qkm+�S��G�m5_ۡm�Z9�����l�QQ|��v�j;����ͤe-��8�p|����n*7.W��Q��l_u���|��Q>��>��x�_�������gVS�;��&�I6�<_0�]���s^�>�bU&�8�Z��ݣ���j�B�������"�h�0�7�c�28�o51��9��c5�Vc��+Mpfq�u��O�ҷݮ<Fqg�����_y��WW����,G.̡\1�ذqXD^��Ő�����^��{^M���W�1�&�//�;*|WўQ�n�>& l��d+�QZ��b�h�|�l;����Z��� (v%��mx�c^���QZ{�$��V�I���K+����(aE�.��N�9T��ʌ�G�+�M}�Vc�kJyS.Y!x���=ڔ�M��"܂���I	S���f<t��qq�I�og͹���RWxF��=�մƼ2�<����a.gd����aA>����E�����Qv{NH����h��)�� f���#��>�p������j\@ܩ7ߤ�^z��m7����DL�u�cGx_��O"�$eM=�(�v�19�L�:*7_�)�Ķ�#)�;(��	,���a�ou��H�UAZo�ew�d���#z1�ض�ܪ�A�;���a&��m?�}T�Î�q��S��&_��Ui�U�(��C�Vݗ�+y�5Ynr�[�m�yÄ���<y�.Y�_�Է�l@MSƤ�&��~��z���5()K�T1.�E��p9��kS������u�m�Y"P.�4!���,�B֊@*5�'̘�0�^C�Y+�Enrz�͡�_ͺи\��ሃS������Q�F�6��G�բ���c+|����6j�|��Lc�hΰ}���cn��>>��>>���m�k;��gY-?zNH]��;f4%??�<�����1J벬�2A�3n�^�~����y���e��?�j�ĸ�����Ǖ!<��Ar��se����\��Ƶ4J1hye������M	"��9�:-�[k�!�e��0t��]�z_�9�_ڲ�!m�1�s`g��n�5��٢�����f�t��s3D�[�>h�d��7-\����|_��7U���kQ)΁k�Zk�e�q�i�hQ#�K�E��y��l��A�k�]�M]��~J1
ˢ(��aO3�=q��̵���g^�F���4�2ƒ�U�A����a�(�^�\���*+Y��/�V5�������L��:�<��� �7x�'�)� M��EQ�M�,}�e}#��Y�G�f��w�og���Z^{mɶ��ɕ��3#Q�@A�H��`��@č����U���EFfdvf]]��U|?�Bu�����=9^�B�ZEN�B9���A�\Ce�*@=���B��Q��^�`e���2�K�M=�$l�!z�[���9�bV�dH{�WP�r��޻K4�F&w N	�M���B�����)j�|��������Ʉ6�d̋�	�Ӣ��`[s��t��Ô:8(PW�=�f;w���֬B��n�X�R�rӶJ_�̝����$-S�JM�,0�[^
Y p�>�Ұ���B��~$U0+�b�r�VR۱X,�8���b�)uۨ�r�F�`WkA%�A薥�ɤ���q/�_�x�^b��&1�s]��YjP�(~P�<N3W��9�|�U]��,�=�I8j����u=�ڸ�,g�%ʶ�¶`Z޳g�kzD&�5�=���t���"- I��:���r����Ct ��:Ȟ�v�M7�$'\`i˭4&�ON���-�j�E�i��w�����A���Z����;|x�����5���=ț�I[�djNh��J�>y��o���~&s��{�%Q�nU��(�*���/;c^nM��?W��37C�R�#Q}Ly�jf5;c�;_�֠�Bp��\廢�7��S�MV�0̅�N���'�1���;����~hB�l�N4�T?���iz�H�qf�2�{髽/��83��.N�i!��%��9WC�j��LwQ���m?Ũ��YՀ� �M��>�v����A�| �b%��Rق�I\��ټ?5L&Ӳ&-��K��tM�-�9[p���7��kD�4�%S���e�Sd�d����7aӊ@� � >��&�|�n9����L�DS����n!��A������W:���&���O��#]����Ķ����6W�.��Uqd�κ �V���J����a����9��łP�{���~�P4�ۢ���f�&<�O�Af�����Ǭ�#���䈭h��u	u0o�c�������6����e�`�Hr"L$���a�?y�4;t����G��ujw�K/�?|v}މ� ���0���A���ӧPK����]RX��O�"򮃯�v���$v��7�U\��TJTY���`e�9�@ֳ���L����U
��u̺���tF�gO���o#����}Sӿ�{�ޑl�7�z,�3��߸7c��'";_�L��1�$�}K��V+T*�{��X��L�=J3W5tyu:h��we$�n������R�$uF���	���j������4�r~���k
y�6P�q%�|���a�B���K��uG�yB��+-�4g��7��)`�ز4�7�
��B�m�&o U��s"�4r p���x��ނs���R��P[����t>I�R0��ȍd����`���/�̎>�	ar���n���m�u��<@⨹gE``�-������Ν�b-���ė�eLpa�	/^@�p?��b%6\��޽���D�?}�Ǭ��rp]��㠒zx����?lzWǰR��%At���m!A�p��^v��|@��	��^�|�ɡ�\)M=���s�(� w�����Lw������a��X�,��~yVD�oݺ	r��G&��c`�s��b>v���:CC_uȐ�ͭ_���]�$}�ikmm����gqlK���LnP�	�ՠa>��Dh^�9@&u�s`I�]��`]`�&=��A�`�l��쳺w��hk�˽o/�r���������)p�T`~���~�ٹ�F1��>e�,-Ej�z�O�aӼL\�h�~��#Ԉ�$.�P���{/?�%%	��p� ���$��b,/��AC�m'l/�v���lƜ�Q����vK���	����ڿ�Q�(s_`0���e~z�7�WY�S^�z����A���fRc��*d@�G�A-�N��u��` ��y�ˍ~uw�9o��,��;�b.w�!����X�5�&���1g��U���3ˉ��"���i��S����:�~�5��+�`#C���h�ͳlrb��q�9h���,z �&&QKǴ��y62bzWp:[>�S�o��6oތ�&������p?�B��j��n��dn쀥�~+�K���P*{��K���Z-]L�Rʯ����ХP����1��i�q�L,��,�R\k�����f�ɷI�uI�1�qe1�8_�rm�T�b�z�!�*�P4Q	
?�2�E�>��z�ã?�� ��ҭ���A�1�N��nq�� M߷&ί�,w��^��Ķռ�F@����/��)r��C���[Qk�t�ɢ�8�����q�cb;�֭W/ϣ�R\ ��Z��� ~ڻ:�#�יJ'�}�����cx���6�.x:��MN��k���T��FP���s�E'9�'RL75~�9N�Y,[zۮ�����g����X+\V5C����,ˤ�Xd�p��^��=ɋ�a;o����d��w��c&p
������ƶ��m��6���M��sr��y�Ўɩq.��im�V���.7�rz���{����c�7��ȱ��/`�Ly��wn��C��Xp��Yf�@K��'ѥ�'���inz:�/E���#X-�-<F�����G.��s�QHհ>��X��~����
r���`��4_6�����Υ2��|��D�gu݄4}[�ss	3�e&�5V�����*�Ďd2��cW�����G��+�{釗����>��p�,<��o�o���.��-�G'B����M�1D�t��5i��R��,����
�\􊾽E�cI�R�29˳�6��m�6$>�cn����f�^&��"�sy7K.l'͡@�8�oY���@&������ߞ�4f9��cƝ��fVM�#�
W_y9eI��d�;�'�޲~|��Ⰽ,�
Z#ng1o_R�:0�À���t��Ё�!-�|.(���X ���e����ʣ��(�/)��f�˾��I��n� �����q��8_|������?�������z�����y���>���|�G��k����/^4���SCCC=��������M�L��u�z.�m��������
�7_����BR�e(�zb��^/4�'��|�vʸ���`�f�8_�Jx�\�k�M�گ8�qC�Uֳ��b�)b�\`p����0m�	S/��M78�v�k����� X�����V���J%@w�Q��7ִ���0�$��M�:�_��<S;< j���ɤ����wO�>2��2�$���fP�T�%�y�r`nkK��pm W� n�4�b��dʍ�V<7���\eW]���!�%A�w4�{pwww	��m`����0��;�py��q�K��k��>k׮]uZyJ�y%�|i�tI�8b>eܣ��^N���m���Q�N�\D�t��Kg��{Y�����t
dL�lM>Cjڎ*��F�������jU���g��0���U�˾�N�����ٜ	�֋.  �\Vn��\5,�O�!ՒO�;��N�X���p�?�q��V$e��W{J�Oۻ����W۹���^���4I�2��iN��O��L��#���B�����=�����e[,Hs�F����F}�|�JeHz5(�^�!h�XpS�RЩm�)#��|��@%��i��n�G�5�|oG�<��ST
������1�dj�!�Ag4\B� � ��+RT'�J�S��R��z��]s`8�N�{�p�G��} z}j/uD�C�E?Y�8�r>Dr<�(q�q嫔���<���ܯ�w�w���'-iv���_'����W����vN�����F�6��AHZ
y����> �~h��/@�?ȶ��4���T}u5{�L�I��J	[V��@a	�w�p��!q8������aAG�^�׻�YUL���]����2_	���j����8� /^q��S;�C��BAZ5��Ͻ�/��?:o&�/�Q{�
E�1P ���4��4P�d� ǎ��td�4%o!2���~=�pc<4����$d�cj

t��`��<�����5�Ft�8��z=�j�9�6���-=�'ޚs�6[�3���Ϛ��s���s�Uu�h�u�-,��D�R��M"M��9�\���h,��_��
��~OOs�����I}�'�9?�_��ҙ�ĺ�;�7BEfhF�)�[?|Jg`
�͈�r�J�B-SQ�����c@���:��Q���v31p��/'�J�ooߛ-�c����Rt�{-�|MG�X^�G@⨬���	U�"'&%5����po��Dj�]��u��fw�#�D��O��ג�\~���DZFP ~�Y�͋b�
&BѨ�i[+����B���JS��ĸY�"�9"	;F���7��s�|gI���r�|>��	��룫-���4�J�FQ���\���4�]�{���.�'�&Mzvv̢�Ky�S���&n�����H�zƻ���SZ�d���]�����A�.�����'�[���$�����m�x>���3�Z#�V+�%%��ך_��	_;g����='Q��t�����ߨ���X�h&'��ddל�Qzw�i���ζ�B<��u�4�/�ˬ��RHmF�]�~�ᱩp��ptcs�������~2��S��@^ff#R��/h�&\�R���fQ>Qϔ��\���!i�o�o�<��ǯ���>3It?�� z��H7D�k핰Y1D_RK����٪�7��߶�?	h)9�$��W���|e�[ul�z9=}��hGࡢ{t�:2w�L�`�7��?>+�4�F�r�]����0Ie��<�;������̛O��$��qm'~f9�^{�O��/�B�u���ٱ~;��i}�P��Hf���&��Vy��W��QP�8\�p%��&�u���n1<�����V�A�D�(�Y!j��(����gںn?�j��$wll�0T�8��Y�-�Lx�ȉp�&�b����Q�1�� ;|�G�v{t�N؝|�Yn��i?���e�=�t.o���5�����<�r�.y�n�L�nAv�ki�Oi�r�\��P?LA��2��+ʬ��g��O�
6V+>�K���"�8�36	��&N݃���<����u�����^�6�Z��։w���-�${_�(2�̆"�[�(v�v��fv^��"����q�We��	?��Ƅ�����礵3�Q���s		�j Te�Yz"��dp{|1�0�lB�����C-5I�&h-��\e,h_Cy.��~��]���9 J�ƻ������,8�t�b^�hM�*2,�����R���[�=������{�k-M��f[*0n�&�a��o��6L�Zvs?���m�C�"���S�-��6I�;�j�&�ۘ0Ȅ�h~L�6w�y�OT@�r7`&Wn��ٺh#��aL4{C|��>¢JAo���֕�D��2vㅯ��g�f��� �Myfc*��7R~�wͣ(,��jg���r���T�� ��|�٣���ɬ���tz��.֧�G�
�:zc_�g����������M���gH��y�H�	)��{��[������s���u\��m!Q���Ů%��=����-�*n�:ץ����#�ʯW�Y�iXp�K��4�-�	-��P�\��P��E1�P1p�>���;l2�-F��>|���s��������ZԊ9�˴�RԞ��N�S#<LT[��U����goX�g@D��{au�����֚\�~��~�`��8(v��07����N�ө<��v�B��$E��O�<�"08�iю�V(������f��}Z�w̑T̸hr��7��x��׳�����(��k%�	�0N��H�ghX��V6�����J����ҭ�sp����:�y"TL2ڒ����,P�S)�U����fi1�~�|#�� ��)i�ݮ����ǽ�ח�����a�Ꞽ.F�S�;���3���D�#}2֭p������5^�*�5�YU�V�n}�s|���gI��nP��� d,'R�K����� �Y��5Q:J�P��S���lb0��$d�K�PCV �ק�{��0�����C|�?��?׮>����2��3�ThMq��'���9�.c�ڽ��X(A�� �v�s�	����vv����X��pq��xYa���qD�oX�݇�b�JW�c����'�����8?����ǧH �4r�=�W�C�k�������3{����8��s*25XM��`���E�@�y�k���8�|��'�*=��\ۜ�r�ߞ���{첇�������w�����ٴ*���;�rꀋgaW(9�]�+�[)��t2�T-�[���̄PMz�0��W�R�DD�5ؑ���tdO��G��9�:�ҕ�`.�����hȶ�`�� �&�������J��0�Om�Ő�6��孈n��:���������@�<��`)��ZA���Ȭ*8d�I��"u�Je�öcIɆ�o��A�q�ԫmN����I��]>�[�W����s3�̃�ae#���*o���MɆ��(��z����,q��r���p��+�0���+�97C�_��Ћ�6p����O��vT6X\�.��y�y��d9]��i����44d��?��x�A�<Z�_�8��鯚�a�A��\��R��M��5�W��ٰ�L��֯wc�v��fb���[>L֦EF�E=`E��Nδ$�9�}��6�4�<�:q΀B�Br�C6\�+�.u1^����g���چP9�)<;��<���2����I�{�
���mv��J�$���Q>4�$
�����`;q�֥�;���7%hm�޼���r�ŀ��;*��)
�H��_�6I�iL8b�� ��i��� ���5������Р��)L6WO�1���C���}ư�Q)�{("�źOv���~��ƕ�M)<h{����ԇ����[���?r�B��h�jT4j����G�Dq�E]A����/���w��,�KK�փ��A_���hy���عMmC%顂�̖&��nٽ�hJ'���݅5G��D�u�)��Jx!$B�wFv���Yr���tf�����N��~G����nol��KW60^�[����t=��lWWTT�<x6�_��]���`�YY�o�%���Ƌ�'�Vʦ�1�ػ�P����j���E4�0z\�)�c�1a��,gߣ~�ń���wp�5�I��Lr�+�x{u��e7�TI�K�B�MHIIt���4�d~����,��b�ʁ=�vU"��Z9��z4����|�6�N�]Lu:�`���vb���ʤ�Ɵ�� $vljH"�a�	��UK@����=Zm~C0�Ό���������NO����g�^�]��{����=ǽ(ہ�]��h=����`M�a��r��p��N½�_YhãG��z�FCZ7�� ��.r��>�	����D���T��S�B<�=�A��1��f.�i�}���G�*�p�P��������ɷ�7rzm���ϯLt��)�苰;5��j���#yc��E|E�X����1[�%+���U�(�_����(/��%V8U�?	�R�+hGg��v�2y%��x�b9<?bZ�xb���%�;;�u�-Ƴy�R+*��4��xغ�Ե8B��$ޠ�ˉ�Yx<�C��$���6�2�q7���lQ#�n���E�@N���� ����ȑ�g�aN�t�R����O�������KLw�1{�FF]4���Q(�3���؋��'�9�ݷ{�=���%����k�?�_��KvȺOǽ5�����O���8\��I�ZbzԅO�㻟�R��j��9O+�>E�)��K-cS2$���"��S��Z�|jW�xl%ݠh���NU�z��vtB�2Ș(W���4]s�=��i��>L��ː���/��j��2�,4x�|G�ɪ���=�'����3�Ν��&z����<#B*��
"��+�l�~=Wr�r0�`ǡڰ/��y��Ii`���
������ ̌�����������iU՝�ǧ��B��z%���n�Kg�|2���z����N��zk�p�����y��hTEl�����
x�!�Ɵ"��wm������J���?�U(d͎�|2���Ns�d��r�Ҿ�X-����k��%��d�{R��ce��oi��R?+2G`9�l
s����9�q��ҝO�Z�=�NpTn��v`,Å
�j
��)�gA(�|��5���좐#�9�]S�3�z��2۾�+vpE��}v�n5�^��
ׂ����ml.+bD��/���3�s��2��?-x	�5YѯJ���k��O�I�b�J�+W�:I5K�3��k<�Ӗ�D�}���?�Q��T�1�Ԓl�y|Մ�\^c��5�X���]5��V��x�f�������w˛���"��}��遞~��'!�ۻMO��6$�U�*�l����Q3)?u�"B,�O���/����s�6LK���˙[�JW��H�bϭvw�(ɷ�Z�@$l"�S�%P�25�i��U�"[�3�������{	�OR`�� �*�9;n��ӳ��wQ4�c���1 yƂ'�XozYrϕܞH����)J �-�j�̰wƳ¿)�Y�X��;��eB�����H?ӊ�K7J�n��CR�W�5������%֜���������(CC���ym�6����>Qe��"Y+�iC�?#����n�˻�@�3��'��x*����/�����^��9�iB-%���Y�Ns)i����:';�Eϳ,�c^��[Dw�� UR4?U#ѼG>T��V�N���FV������%_� )|U>YOGS�6]�����ȕu��ƓC{��舼��YƐbn�F�p�Khϭ�)�yU�a��
'�z5�]M��VVVn����z�?�wLEA�
*�!�Swӣ�u���J2�=���Juu��}e�'�	*)~K~���iu��Ơ�����pI�o�l-�g���КŦ}J�%Y#Ny+3h�4�!�"��B��F윕�Mv�����o�ݷ�������O�Ѭ��ˈ/��@l��}wA>1����g���${YY��=
���m{��k�}gE��c�!B��;�2F�2����6jMd��{���uaCRN1����"�U1sRQl=} �[9;���Z�!���Ƥ�E�K=}�����^w�W��{��������� ���S��K�
��.<��T��؋;>>^3��'��� <H�f�3�M�2{Kab�`C�m���~�0�_��%'L�"\��7�*�X�u�e���G��f�͋��<��.?I���ƥuY���Y[[u���p*���$L"�t1��f2�>0,�,��Җ)�9���l.騱L�����2k�����<�(���T_J��s� �L��t�1�NJ0�]b4���F���
;����g4[H��r����曞��^�CM��NK������**�Q�gO��23%�2�P���K���^�.�	��F�<����a��wW��9 ҹ���:G͙�]��UP.5Xb���1qo�z].��|nm�>�wT$��z�y-��Z2ꠋ����&��EP�+`U5�դt��~`@vqh-'7W&����Nl�7U����L�ɜ�s\4��\Nu�����<ti�._ӻO��P�Ҵ��	���y2yC�{#�%��!�q��K�+#O'��b�AF�%to^��˝4g�c���\�ǯ1�ew�ns����{���"�.6{;�W�M�\U!ssD�6�!�1���" �ɖ6@8)���M�b�l������]E�H�D�i#`X�#}�
*�q�=�Q�D26_c������H��MG�2rdF�[�=_"F�Uh�C�w��~� !%����mo��,5VUV�[~Κ'$LyAzkA����$"n;Dnv�#Vs�]vœp�.��m��p+''�խ��5��5O�a�$Sߕ��gd�M�/�Vp~�r����w���DNYl��8'*�(㊥�t�����QI���]��‸ݻv�����A��0�C�t�'��^�j�~�����
�4�T����}F�|(��a���Z��x��Y�\�� *i���*4llb�UU-�����dX�E~މ�J��ȹ�w`?��(c�7�M�k!N���dY>k��伥#��2��Z���-_t�*��T/$'�a��ބ�tkn����V1(��R���^s�d]�O��QLb6O+�vx�__�">����^�	{/�,�"��ߟnN�2�?���
��3��=r���;�w5��u$v�P�+���}8��O��A^6��>���6��
}|G�i��6�ߖ�P|Z�w��e-¾ۼ�2������[H���'	��)�0�RCut5t�@फ�UT��;JY-�7V�,��kw��'q�hZ��]���i�j�P(��|߽Ar
����Ζ+{�nk����z�\�=�:����~�Cwͳ^�ѐ���L�:��<�H�=�y[݃�f�;����P8H�3�8�>4꣣��ܸ�ܨk\��G��9E��o���;	�d��|&��h��c8l˗@���,fbJ�n�#���ٿt4_����Wb�݉��5�?y<��)B�Lz��@U��ܮz����[��p��.�C~֒N16;��ѓv��amɤ Å��t�d�/�i�����rҢ��VtW��<q��@������� �:V�R���M�6wO"<�N�onD�(��p�����J�{z��:0�A����;�&c�k�ܪ��ho7���^Na^�1�ɛ/5��@O`�:/�]����d��2S�w�A��.n���\1S��a�`���� ���@�T���ѽ��z;kzz�	郓t/���,ɚ^s�>2��������$�����n��`�o*����Z8�ݽ�%R�$��oԵKE��|?@x�M�T���L��자Qe�mm�x�:�z�&Us1*�L:;yt_�|n_7l����_7to��3���5��@Of?�|<�W�I�TT,J�&�P)�z_��W��K]� Q��o�9B�3"�6|#�"�"�'�^���M����Y=eߦ%�+���r�Ԉ������`���܃l�})>[���>��u��J�9�{�~�*��c��|�\75��އ����u�=��f�OМ�-���$� F��^VNۊ����9DwZ@���CFP��O�g\*�9.���n�}�C_H������ ��x���J�R����"OZSX�U+ݓK�4�ا�����5O^�Ի_�+ېJ���{�7���;�^����7g�΅�p�
2����1���5�ܚPG��Kk�#��eݓ�>��mjQ�9R�x�E���x|vf��D�0�-��������x&�{ԷY3��z}y�ӷ�-鴴��}ʛ��<l��"K+`����[dm�i%��5��5}��qc��<H�����ӂ1Fq�җp8����e���}N�1�+`E�և�<��%$W	�>;���{Ǻ��Kz��˄�9��#��4�І���S��T��^Q�Zj6�!:m(��1���2̒�D���X^��߹Q�� �)��]��kXS?s�&Z��l������e����hy0	��H�È.��p\�*�t�a�K�c׮s��f�݊��؅�C���X�oRjl?FM(�1x(��Cvhrif�r���2�7@�7���:��u��yᰥ⥇y�/ к\dH�-���-//�� ��:���<3�<�LE:K���~br��H������X��B��A��X�|+���|��#�?�s�թ�='HT�Ƭ��[�Z,�8P{�0�z,F��IN�D�F���n�~��]Ⱦ��k!`�ֶ���Q���cZ���iWv��>�OY�ӿ��@i��L�Oq�y�u]pN��@M�g�1_�7ܟ�D+c��L��]�<V?x��ݮ��軳:�;��;k5�v���'��5�r_�t|���ʎ����\M��::�����|��<�N�쏡��qҮ�B1ߏ�b���S�Π�|""c((����jN-E�&�j賹�WQtA�u{���ƂA�/�rSח܂q/�5�Ė粜QN��)�

8!Ti�`rq���E�@�Db�S�ҙ*{����hE����HNy��[�Y-+���10//+r_ d	I��;��Ĩ�����c��<�����k�� ��Wiؿ��U���OM<Y��R'a��V��L>���3�5`�����[Yfǚ�o
����S��VGN��t�kz�!�Q^�D�� |��>쾆�8k�6g�qJ���K.���k�_J�+�*љ��ca!���*V.c�۽5?2�������}����Z+s�����-���Ȉ*�׸�AG���w�QR>'
Z�©�Šbֲ�B"@��5'���}�q������\��G�ߕ�=�P�{����oe--��~�Ð@]�	u�Su�[�]�/��k����J{�閵��	���곀tr5�����Gt?�s��j��s8:�f���;�Ko|�����Ѝ��.O�������z�c}@z�W�m�Q=|6�^��$I(����I,3����N2 R�>`(�d]ʶ����?1;�Z�Wu�y�T�/ |z��d���A���5��/�A�MaQ���$�lG�������.���l8F�&.�㏩��ÛV��WA�]��$*vS�����N��|*�b�(��Mb�C?��(lgG�ۮ�ˁ��3�T/����j�z��Z;l{�{�d������\���6����X� 7�����1=^]R��'\�Og�O8�4�R3�-'������)�)��B�P�w�͂�?e�����"[K;�$P�G�B��e���Qv�봺!�"��B�V==�N��b���{�ձQ����II(+��|Wu�Gh��� �;tv�� ����_v�=[�D<Ef�Q~G���7\g]boFNT�x���D�,�&�<t��-,�XhYX�y�ᑂ��v�KY� d?�:��u�8�.:�`P.)���WQ�*��q�ڨ�ѥ� )��	����������� Z-���X�#Sf��I���[�0���=�X{�iθ{+��D�ڃX"�w�y����Gc�W��p�C���[��כ1,����2�&mX��еj(�WB�!����3����x5��"��������	2<'v�dx;�V���MgN`�3g[������(��E�u��K��=�Xs��)�HD>Jff�j���?�.���&N�(�ޗsgaR�ռn6��{��T3"M�D�,v����?$�?����Olr����z�#HI'l!��g�}P�<��p���d�$�UVK���}7���A�����p�@tAc#�=�&E	������%^K*� ;/ۊ��9�f�8aX�$� [���\H���U�<n\"�S�WF�/-ςp[���ѓl�0Es��l7ϵg��)!�kL{ض�z3UTk_ग़Dd�%R�s;K��q������^C�v;��C�K\�v�l�ff��0�	Yi���$-B(��P��ѱ���0��;�M�ۚҌ��9�~n	~���m'���ⓨ)lUo�-[`���R�

!L���g�e�+Xq*�?��V�Y�o.d���uZ+{$J1�fl�N^tlYX^�5�f��'k�y������Q�4i샏�r����P���)�á�ޟ*a�	�̩(����ʾ��pKz���� `4%;��K��0����56��ݏ�YtS6�iu1Ĝ	��k�-|<�3�\ĊD�m�dg��X\�|�u�%v�[��8�F�$lև��]Ȱ�m<����2����X�-3i�g����/���Y&��,�+�!Όk���՗�qaohy�k�+l���x�"�Wt�G�n��y����x�x��WJdҔU-a'X�7�V�a�X��t��p����s�BKU)�U7ta�vn�D������C.�ٌ	ސ�������C���D����X�L�-���JPh���$V��f�W��H{l��{��zqpq�U�o ���4(!݄zJR+���{ySr�Vlf�!#<��K�ң.*�;}�C�71���*�Tđ]{�G;f{�]��5Ʈ�ƸM\��{�C�G��:|^h��r��mm���a�T��>��k����x�_Bj�n+?�%P��Xf�c%�>=z� ����M[-���Eh�����0F�I�y���{�.e�&ŧ��_;� 6πh��E��}�h£d%tC��n�Bt��*�jyvv�z�s�A��tH��
7xa�@x��_`&�A;�����%�ğ���'�;�ke��	5A� ����h� _�\�dc#�r3{Br�L�0��sXj���h,]|�̌�o����Ӂ/Rڔ����O&�Z�)~��q_�TM�S�ά�,N��cZ����D���pnb ��-�����'Ĵ��G���#-�Hƒ�E�1XT���}�ʽ��jpz�z���|���x�X��B��H�:��@����/����p�4�����e���1U�R����<j�ٚe��J-�1�BqE���I�W nI�L�Xd�#�S��0������W��kUr���d0����֢*���{e�S�X}-V��X��������_������hə�ܴ�ɡ([b�{"®W"9�ٖ蜂�X-d�V�]O����^r�R��;�=ǿ���٘Q��"�w�t�}ZXCЧ/7>�0����}�'0�hjٮw7t���z���3��oV�҂<��۹�o�Ke������$�[%WTR'1�ssN0�!;4���� ��3�½ѝ�ѱZ���j�_�}�Ia
Ð�xSr�O�è�>����t0���h�GQ`��.�x��ٹ���l��m���/�5�{37�&�i��d��SYJ�G�O��K�^��#oM�>:
����.�����?��h3Fhh3�����y�n0�7c�٦��2c�%������d�G�$S /m�o���{E3��/[��$)C��H��a�ǹ����+��S�h����٘�2��q�zh#�3�kBm�YW
��3L�o�OJpź��V�٭���mEJz�<pݭ�O���}�<M�(t�����x�M�&�P�gۓa�Yx�������ݏ^���kcR����̮ab��T��X�Kv�-6���$������9�,�e�"��3�hb�}�9��N���I
/��H�((F��+�ۉɵ��ߪ�:2��U�kvz����e4?���߶g4��t�8>}���4w�va�b�R�z/�bK��ι*d�8�c2.�U��i-��7�nDj���(�ɖ�+Q}�n�d��uj����I���Ħ�S�J;饁qK?ol��N��ߗL����9�,Ea�,N��*�L�H�C)ICq�=r�~�z����0�č�7����/��ZS�57���SȲ��:��9l�}���bbO 8�PGЏ�l�wx�:��\N���� ����fs�R�3`��kA��S�����֣{VU<po�������\|fy��Y�Zߓ*cßG4����M�^�s2��'�ϵe����vz8��1���~��Z�0�1�\�M�V�I)a���	'����)��0�V�]6~�qu�d��L���+�@�s_�Fv�Ncl*�3�����:�)��/v��\w
i����i	�{�q���@q]"��q�����[�P�8춤����@�M��~ �Q%�|#��p73G��)7�_�u����ͶE.?�Bj-ZֽP�]�HO+�����}�:I�0���f���~C��(6TaWL����,�p��R� ��Ǿ�n,E�]�.*�)|�3z�g\��w�_Լ�����K}>kw�Nc���7��q���]�$ܿ?�6q*�3��ܥGl�K[��������n���[a����e����>��wj�?bԥ/ѼSL��x`m6N�x���yV��P+��Q:zyɒ���~�v������b���U���E�����!��ލ���/ϯM9�?� ��|��J��έ-	I�J�|R���ǳ��S\
"=-�Hd�*e����]�"�f�$1��姧T��SgfԂ��t*��0Jc��)ZN�췔��b�[ze�Qh0�E����_Ws��v)LGtT�wY�{�#��!��U��n����t�#?(�4
f	Fl�����;���&��5�v����%�c��9*��B��f���R�x5�}2B�t[����6����l�orƵ�V�G�����ڮ�5�b���+�d��[��]l�F����>��PT���Qݶ�Hl�ĺs�GQ��az�e��O��̆��܃?*�P~I���/�+�KXѶ���"��/��Q�F1�����q�����-a`oo��b��u������$��t(���c�vo���d������ttw	a\���A�1������#��tڲ�u�h�4����n�����A����[&�E��36�����룼a8�qu[`��v���/�2ǌ\�+$�glQ�� 7�y��"��	�V��m���lW���(j�[AAW'����Y���6:ؘ\R�;��C>�VM���Æ����M����]{f�r̙�(�3����-O�����~q�����4��$�S�jBh�$/�Dn:p�!z-�D8�~t>�&����0��X�������?=]�n�3nD�Ӎ-����L�>��p��Ru&�￾R'�	��ȿ$�a:x���i�����pd����`��9_��n��®vUE����V��F�	�$b>�/��5��1a(NWU.]��XYlx
%)Th�K-g��%�0����?S"���,����
�#�_t��5�.�=�P	ײm���פ���W*��༵�'��L^&�50�.='r�&J��pE��ɃĽ�r|�\�'EU�M"���rKF���h�BÄy,�t�[<�c��eYY#*M@��H-�\��{+�Xܻ!a�U����#+U�G:�8<�3�$�r�0�崪�4��p��*B�[���ɽh׹5�yv�f���-هn�ڱ˦w1<o<CC?�����g�֙/�����s�Gq�ב�?�u9gF�?\j�j��͋��ڱi�i��v�~�vc��@�"1���ɠ�k,;_��Z�X5�?zɚ���'�>����?�=��^�D�QPPk��W8���&����f���)�h���n~�	��v^�B�\V���@��X�5lGA����5�JM�H�h,0�~��S��6;����:�!�]IL�ɕ�5�+��$����� �wE�gVѸ4VT�F�S�{Q�6�i�@�w�gmם'����/sΠ>H�3;�r�b��{���H��\!<ȗV#��;���`���5��C/���?�_{6KhRuG(�D
>��r�X!���d��C�N���%�@b�w}l,� o�D��s�'^yװ�F��,pk�?�_�/���#ȕ����q:0�^20�j�4N_��3��;%n�Ae��G�63ʥ6��Ya����������W��<�1SF�폯��&�Ծ;��=M��e�n�~�Ư�������6�ߴȖUc�ղ�C�±@�� ��́<��3Zƈ�V���&�
O-�?Q5iWL�8���(����ݴ� ζ�(o5'��&Z���G������`���Ã���]�t��� ��1=ӹ6���[
�������I���f�?�l#��W���	�S�<*f�o>z�,��9��L���U�����	r�����2���F�oL;WU��Bw=�]��G��[������DQ��J�7h|/Oo����z��Ty��-�����Od��ʖH1p��q2�9<)JV7�%�g����}\�j� 
�֖j��6kF������K�h�Ӄ�_
��3Y�����/�-XbЋ^�7�0{����LV���F`� ����4y��X�Zp�C��{x8uvs�m?~s3v�ˤ�P��Ɔ��{� �n�:cr�����@��1}�k���Ŧ�VBusk�S3����-w+2�톄�l�(�h�ɮ�A����YE俶i� b����?ol�'�J�.m)����V$+I=�*�f���Xԉ��q�����J �ھ2��'" id�%D�B�>�.�d��d�g�=O�@fPO����ʬP���[�r�;���C�*#���{0q�N������3e��o-��*<{�tw�3��$DB�p�9h�W=�^$W �r��L���o�Bx�3L����=.��w�ԋ��WW�{��֪�X�I�<pz���e�aC�MK�1�B������6N�(tk�/��v��!�O1����ձ�V�
���E&�S! +���i#�&�e��T���kM�߸�9��(�����:b�?���$:��-^�֠�������y��Z4#O���T������G����6ۡЖ��Q������ϡ@mT�,����z���ݷ��nWvJ���[}r��PF�< �X���T#�������(E�����x`��6����-�I2VN����r�/�p: {/V6�2��7{����I�JAۢ,�㗕=[)�|�'��t��FF�L�	����óԈ�)2Z�@|��ǚ����'��3/F�]�U�3��M�m��!�Y>�١� p��g�7��{�����2�%r��glaR{h[2���iH4���Ub8.JZ>"F�z��s�Oh��ӈ�IcyF.�;�YL>h7%�~jy�<!9��2�rRRV�~cp�	�d1;�⹊Xf>a��6���P��!o�J(3��3�5'��u�`}�� �4����w7�|�-o��QDɄ`�-6ZO���C/+�&T�l�95�I8���'�����t?Z@E�W��O���듨�Sl�]�y0�{?�S����	i��0y��A��=PՏ��S8�GTP��?����widWK����_]5P��GM.�\�Yʛ�m��<��A�؃'��Gq�����/�HȕYͦ�y�M���Z_����6]��Ii��u"�H�6������$��������������c� �l�����r�@3%[�;��)�.
��胧A���(�2����Y b�mb$uc(��:���QS*,�6�̳��M��#�U�:;�1ƈD����}����4��DU�
�'&dJᜒᨙ\@��LLM�>�+�t�6m�*���]�̊�/�lc�_������>�(Q��[o������v:�X:'��6%˞=�n�R*t����en�|����	���U��,|�<T#3alA{|��L�!�K`�6]t?��c��X �j=��\�p�.�F��I��[:��+��Q�T�͂7Q[�^�}y�tT~�m�/�?�lC�G���NY��.^x��5^�)��{׭W���-Y���+|���"��/�G�uF�,B</6$��!�,����넋3D�'�0�4MeZ<��8���=�aZ��G���B����>x �e�� ����L��� ���ESH�R�o�#�K��@�?�������q� ��}��"S#e�PK   �i;Y�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   �i;Y�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �i;Y�i{J�� � /   images/bbc1753c-83ed-490f-889e-b8df35028df1.png�W[]Ԯ]��kq���[�8w/�.�]���^(R��{q+�P
�x�s����/�@HvF�^k�{^�\+Q*J��HDH�޽C�J��{��� �A��/dw��At긾{���z�JeD� yR�B[�RN����w�"` �߽#z���T>��3�����X���<v���H��8�'���I�kxe�t�;/d����d@��ÿ'G��L�#��"Š+�d�Z��o�L���am������ء��w�W�sԳ�����69	(W�Ή��<�oƖ�8{���1��n���Ȍ�1)���sm6�x����1����~�QFq���1��.���%N�o����0h&�����w��y��v���>
�����ŝK��L� ;{�%�j�ʁ?.bD��Pɤ���(nFѝ�x�%('UT\L����}qq!|Ղ�vP]���yU!��&�h����MMM,HI�O/�:�98���
��y�~���'��7�ko�$v4h�iW�)Z�x�F��--�����ڼ�J�"�/���SMⶃL�o��k�bJ�W %M�T�^SS㾽��iB@Ġ~zz:�b�����+���SR�{
Hu�����|�3��̘Y���poxAtF����]s���5;;�$�/--݅��I��������I-|��෱�T��X,���߹vJ����5�������p����l�����S5󀄘
�QϠ�W���P>l���;����������}��L�2����Y�����ťv᣼�����%�!�����dC��;n�	A�	��vAx��P�(33))����D���ޞ����dɁp��u������EkgQ@��rM�23K2���?
EDn�6�"\��M��/Xo������%UC��{��r<3�?�����tg�'T�뉤G }e7����2=.�;�2�r������W�������L������d��_�.Q�h�5-P�T%�Zh@l��A���´!�+VO!X���C��l�uZ��BH���A�/�U.,�-s��x���w��kq?�������߮S%�|����I���I�:Z�to!����8�'�uaxn�븦TS]9j[���|8��չn8.���v��
E���J]�k<�ц�5=+�49����hT\g����$�,"��eXSiԁ4����f�ߴ�����,6��>cG�ܺ곧�sss�PQQW�j�]vG��;%�L����&���D�IP�!�$O-,������_�o���l�|��_�m�W���{F@��$Wk���z�{�P��\�ķ�j9D�"�M(�E)E;�0&�x'4�-q�m��i��Qۄc��������_^Y�jhly	�~q��������t�t��ٽ�8#�
N���+66G{ss�_��bQ*���c�.9��Tu�[[� K.!]�bm���I��$�9�:Ӽ�Z�?�@5=�/�/��m(�<+�JL��Oy��dG�E����[\��v�&[[[I��ʼ�����/���M_�,�UՌ����"Br`��W�������Rb嫎 j^�G*�r�sg�C���[/`
Bc���ȣ�G��~*�3LI`����d*��_i��.�����hA��V$U(Y���=[L�����nX��!�&"����l	�U��3������� '��<3�O�ݝ�?��h���'gtt�ʂD�
qpΤ�anV�M(�R5}=�R�A_hT�M�^p���-���U��M�\Tfɬ�����F�GAj�hr��F��f�Lu�2�YX��L�^^���;d#D8Ʉ��8n��o�d���~�"L�ga_�3PHy����������+�w~?���u,>�����Z�D��27��y
����l^6=y�
��R��&��C�vw1�?8�1t�K����T��q�Srw\��/T�zx�VX���&��uc�����I�s8���ʆt�Ӧ)�p�����o�~�$��/o`��	�ż�K��[т/���\Z^n�8a�$n����>՘�:� K�E��5RP�	V*l �VL%�s%�W����4�D��O5�D[�>l�V�	�Il�`ȿ���lN�8����j	�(�3'��˷�5�>�����֨�UHd�  �_D䬪�&wۥ?p��#0K�D��a}7fAħ+��D����V�.�C_�ᆠf��ϟ?��l�����{���r��L�aJ�qU�2j����W}�$|rHI���p��� �E�j�'�:T��r+�4��h�!u��~ڌL.C�����PIA�ĥE?M��@K��nX���������&dog�>v�~�&�}�?�←?�e5��A^��='��P�� .�X/Y�
����< ��%�aV��'E	�\�N��I�;h�<�HK���B�������l���]z��F����l]Z����5�$��5����#�ss�OO�֧؇�Jk�#cj��c�jjj #�<�
�2`@����-AջnaeM YS�k9�g�}�Y;��yž��XZN%������֖�O5'=}y�a��JC�y؁��d�0&��c��$;�?ٵo���o,-uoNmv�j�y��)hT�~��J>��	P{����n�ӮX��kɯ6�����*�diT�}X�=#'whhH���w��������.�3ƶ�FHSw٣H��+����{����0}�'CUU�C��V�~WJꮟ͇��5v(�>��3�ӫ"#!���75�����RYJ!��׉}+���/`��E�9󩕬�F���V������8���ki1D+�%����JR�������{#2�y�,���A+q�����.�?�9>��]���th�H�@sp�c�I�a�[�T'�{�z�c�7�<��T/�g�jjX��w�3SS7��4�0�I�3u��k��5��� EY��y�|�8��-���ҹ�j��pn..�Ϛ����¨U`��l81L���}⓾|)��0tm�e�؟�E��׆�hs�I$O�c�IR�O�T/�OK�p!D���t�����1X!2
|����M������Mx�b}���3�ស�E���6�R����a�.+����T��p�P�#���iӦ��z��22 d(o)S��2[���fLa���l�7lL?���Ӫ�����9��t=�6ѱ�I���\S0���+��=�����tT	7/o���&�-+4^ۥ*ʋ��P����&�ʮF�5<<,�G���mH����K����<�/�G���#D��o�
�1�d�k���7"�;*/��S�0V�0�i8���8�u}:���),4C"��`�t�Vbt����],�嘽*�`e�K%�v4ʔJU�x_CV	��8���bY��G[��5�U&�ѼK�tR(}�7����� �!����(��:~�=�����{O�oo�p�*������>�p����-N�����^�.i�E�e���Q#F�:��M������!���<c���x��Е��'�X @��|�a�d��e����y�,�˾�WA[�͠�!J�n*7� P����� ׋�Fm{���a��J��� �j
˟�]w>�°�����'N�ɩ��Y�rx|����{Abi��0�AOuȍ5��5�����l���Q�� ��ѯ̂;^>�V�;+"���7Cz�<��,^G>׽��t��F�dxx�/|P@����II��5�l�d��޹ۍQU�!�%룘���)p"8� r�4��}1�LN�tXn�T��g;5A����d<�}�5��	xqrtq����}*	�sX�i��9��Z�RI�����֬j���0�pB������j����k)�c#����~�AAP�����I�}ٚ��������fg�!�6�?�gT�=�����G#$�i����JQ8^E���/5P������w�
$�Ʉ}�t���U��F6�膇������(��� �=�����GS�	������"ی�:&����p�n;#��xUI��Ia��V��n���D%`�<�_"Ne�{`��$]���eIBQ���&�q%�h�O��-*�8F[����`�Mw�iX$� ��^[�2�6��X:�9)N�O
δ4��*�GGr�4�1���`FZ�)���	E3V���/Q��?.
2!�A��A���͊�A�7||�S33�'6{k�DAIx� ,v}���N��N%E�Ӓ���
�.eI�Q�)
���O���e.�;;��m����
���׾\G̺���O'��zZy�--/V�(S�G�MQҢBb^��	�4�Ʊ|���(�3��W��d��cR��O<z�L���`B
�}\
X�q5eQ�2�P��J�c�%sU>Aп"��Ŀb�GvY��b��/�qˑI�(K~������%�@Ŕ-�e�Cm�V�a3ee����-��C_H�܊���(M�{����k?C9R���Fo�z��mF���
�k�nO�eBB����XJIdN�xu�8��|�2]KOO�l�H@���v�`�aAK�R�t�/ �M�<?��G��п�4ִx��Ik]}�S� ��Z�l�0W�dy�	zfV*ƎH���F���JƲ���(1� r�C��z FN�1���I`sd}�|l��ϊ\ �$���}h��ӪɁ�0�v�¥��������XXXRpl�+���;��Uҵz�,��a�6���˰������5��������:�D۷�U�%����GD����v>^f)�D7f ���՟5ӡ� U��*6!�*_"�`�e���X<�n�����Ap�Ni�+�^{�}i� �|p�}a�����yW}=��[��Z��/���PyR!K4�SGS��E���� ����16�tP���mw���b�9:y��Xe0β�^f��|�@�K9��e�����:Lj�:��E��2��:ݣj��p�nB+x��i� L���O�'3���}V���xӇܫ*�؃!�������Qsrr��|O�������`�k��!��)�FUxx��a��]F��f��'KDn����)NJN����R~��&f���2� �&4f��f�z�����vy���d<�{�� 0J�(dp:�#��w~�|�����5��Q��2��@t�fA��j�kO��]��;=`���eM:�>��T�����,��0[�n�����嚃J��Eኄ��W �+ETض6��F�P�]o
��Y&"`��i1	�M!R�q��|5\�}��#\��_aш��l�Rf�OOי/@N��^��c��k�:�J_���	ѸQs77�]ۿ����%�с����0�P]خ!N!
���4ڷ����%��Z�^�q�'��>F� �,}�Jf5hm(((��B%kDJH�<(%Eq����'���Њ�T��,�B�Z**:�Y�@#���fJ��}A�ҡ�"�(J*Ud
u���o��Eu,2�(����r[q,!k�E�4~XM��T�b(�ʭ����d�J�����25l�by��e�ӊL��Ta'�9����3�糶�i�I�����I����x�o����K-�l������ku��QA*�2�t=�eU�t,_0���s�F٦�0��x#Rj����Q�,��U���nj�bO���^���C�x���z�\QQ1�Pk������3t�ć�[>0H�m�\y��p<�{�By##Va�ًp�.QrPC�z ��`�Q��4exdT�-L�\&t�q+aH��`��h�>CG'zv3���PUP@���4|%'H�✣��5'����;M�6����d�tC޸[���n��7���0�Gd��v�R�xc�6$$���({"o��&{�<�e�,t����*��J�rZ� i�� i���wG��Q�y�����t����l��P�ה� z��;��F��hA��ۭ���芿]^B4ȱ�5y/���d����s����U�T�kh@�3��.���1�S����B[LGxkh#��*��0����1$����B�3-ϕm�i�i �9e�K��k��;<{�{7����hl�/nkk3��eO��?�Քи6Me�ATW=��!�` V�spp�xd�OOO�ߓ| ~Ûi�p�לSH5!�||߅(N��l1"�ۀr��&O���09j����E���o����>���<��x�/y�����M��l""-M���7�q壛�$Ρ�j&���^'Y��kwG#bbbBЗ�e8@N�6�6�EH�DNKSi��)��`��Zע�)���,�瓃g��Ut6���f"���N�=���R���(���$����Sr9��,��GA�J�˻���l6:9�߅8�{���8:��̰b��������;���������9�e���$ƨ������m-.!����0�;������F�e�Wu)�ȣ|>�G8��`���0ؾ�8I�t���4<ژ�Ǐ+J]��A��ś���q�i+*(m@���h*p�'9s����̔S�SC+��B,���ں�x��*�5헴 i�EY�ݹ���O>=�/����=7]��������Q�[\_1��$�G��Q[�CSyJ�ۻx��N+P5͌U���,J�q��rX:����9��9���E��f9=6�ddֹ���/����t��:GӒ��<�ݯ~����1:�U¢̐��G�='"�#Eny��l�&5�0jVY}3�8� ����odd�"���У7i�O������<L�˵ɮ� 	��'tYc�<)k���;f�g��W�e6#�kN��z�������O/"N��̖*Wrԡ��)�?}�dij
�ԉ�" �S�$�1�R�R��9m\`0���ϢBg�Lc1����{��%�8��.�;`!��>�x&���'F�"Ep'`�h�(4 �H���?�e��H�Sj�w͏������i���� $�<닊~���z�w�;m��=�c�����V�*++ᑑc�r�N9c�)e��'�ޖ��s��0('j
��5G������	c�A	$(�
yo�^l_��=�ZѨ�tBL>T��*�����J�n��)�W������y=�ԫ,��#��Fo���!�����'"I�6>%+��B`C��� \�D���\�!��'Ze]09�5��D��&�8��mOgs��^&��z���I��[T��L�~w�!V2M�%-�[���j��§���U�" !�jT
��##� [U�:� ���E���󥥦����&fd�˹�Is���러�[�8wu�O�13�Nof���1�[�q��h�td���?����o���+�喨�R�7��j�g��'�f�L��֖�'��a��&�J��G@�`#ZuE���L�2E���1��wa�j���[�'#�������R+v!�!��m�A�� ���6�yʏ��P:W`l,*Y�>�c�� ��ݰr<���mP���EB`��7�\�Uz|��h>�����U������:�t�J��XI�)�0�6��q�wWy�z������^	�ʕZ��O���cnr2(�����x�\����^X
1�k�Jʢ�3�y�Sx%�<><}H����~e�QS�p�ꋢ�<[V Z9��;�\�����N�4�p�e��M�����櫵椷�eDG���7�����.��
�������G`��5��4#�Q~^��T3?]��	�e�R��!M���IzNx�M`��1:����S�H��$A���!�P"��{�h�JVM����X�D���'G���E�
��ZR86v��E��N}��l�b3P�'���쁘���������p���4J���ao;��Hy������6@��j��#��N���GG��T��1���Z[LgWp���b���ôC�
z�>
�fp���+�t��V�v��fOYAur�ے������ȅ/$���~z�a=88���(�����86-�+9���hNEPdv�Kǰ\W�=�ޥ�R����]u�[^^��G�t>�*��w!X���`ڋ�4evs�@a���B�2��p!��҉��u!��Bp�tTT�T;{H�'�����rl�ܻ���QM	-�1��4���p(�[=/f+��'߄r�����PG����<�*mbb������ׯ%_��Q���H�`��p�H�P�7���&�D��DE_��L�KKK����k��U�}[�܀��������7�ʰ+`�#/��DB��#ܝ�j� ׆(GSӭ'\������ݨљ7F�����I X���8?����z����;��L6kb.֞�p!鲡�[��2 8.h�5x�	���l<�]V�C����p�g��e!!� �sR�jw ��������333i��L�_*����c�D��)��&\W�h�=N��ڽn��8('�0{l@܉�+��w���t��ld�w�3�<<GOO?jq=R��
�훲|�����l1T
9ڂL0�F[m��&{R� �4-W��:����U��=��h���	^>�{�eE���y�ZZ77���H���~�ڛ���!��s���Ó��P�iB__��G�ػ�5�o�MO%�-�H!a�hs0�k�2�wW��V���V]��Ƞ��hӚ��|6�E�.T���҅Վ�e�I�.�������(�:Yiv�Y9U�����36![$U�Z���umWY����Ѫ�oɎ�>fI;�
��o�Em�kv�BeV��x��z�TH�2KI��챽�5cZ�j�cV����n��e|	�7,+��	�*���ss}lx?��x�s�������4�\���M�� -�O�nZ�
*P�Rɫ_@iSE�[1<�_����հd/��������}���\��v{.�������:Y�>�B�`@"3�t5w�T[!J=Fy���I�8�&�[�S�Y�~��icZ�c��ӯw��ף@y�,�e->�B�Sk�T~���e}}a�2���az&�*�:���������z�DAЦkqc�ukxw�A �D	�>�I����9��M�y��n��c�S7z ��Ϧ���B��y��>=a��`�i=�����𧘢�HLv��wRc�F�n��6t=~��_J��|���&�/��z�-�3���x»�P��� �����C��2Tj%2���o�< �Z���V��=µ(�?��>�Y���՜�����I��pS�S�F�s��4�#�!�a�ߝ�@�����o�Lq�����9PI��zz��H&��j ��O�\'�nں���ܿ�"B�q�O�De�nC����?�P���8(���OZ�p�p8)���y`�kIU?��K�&&��R$�2��9�C���R-$�A�T�?EN�p��듚��:"@��|��U@��"uvrb�dn�Wзg�v}N����n�}�����s���7�E�;��L&F��Y����ɰ�������c�i4�Z���2�� �#����%�����e���Nk0ț��� ȧ��^�ڼ�v��w��խw��>?:��[��71�� ����5��NB�]�L���Z2�S�貿
��ߴkD������6�+������$w�V@���$�������M!���6.�X������yĉ��v����դf�����g��}c����;w�T���e���Z�ッ�X�yYY+�N.�o��^;ǱƦ���;;�Es��M�A �.��i4:������w|\?d#ð�C�n� )@�8��y�
`y��G#�a���t!x���X�e�A;|��~�+-�&A_�J���x�����L�ݮ"Μ�*Br ��<}8�#�x<O��ѹ����'��6'�˲Ѹ´�rQ/��|��_*�����Ĉ�;#%��ww:���)/�Qش]����z�>K��G�|#���N�O��#�y�A0_�� ��+�7���ږ	�����e����?9	���LUS�� ��PxUQ~�)p�C���Z���i��'�j�o�9T|���b��m��� hx����1ee兺@����-p,	�� �2:�� M��J��j�����w��Ӥ��V��л�����}���^�X��9iL�-��?�Nj���;���`�l�r&����ËJ�\#-&�-�1h��N��A�/qQ���?G�6�߉��SS*��[	��?�++?�kDd6�����6�S�G��x�O���{X� }���t�T���j�L���dem���/3�j��36��`�!.%���!N3�g��֑�󻫯+�8�����p?��s�Cs�-GFc��i�#唄��μi��������/�����,^Q-�y��j'�*hv�5SS�ܛ��|�r��|�ێɉ��Ј�u��\]�'ÝB<�LK��\)$��L?E&R�Gx�.7�@Ԩ`?�R"�m4���H�K���\dmc�(ܽ��i�w���[8e��
��C�pz �/G/�q����+����zf�?�_Vޕ�����R���*�2~��(�a�9&>}MI�Ҭ��W�Ԝw�0o�qȣ0Ь1=���Q�tήg���I{�}�ؒ�/�Cl߳kjXm� �T�qHlH��	���j��=��.9)t9��f�3���f`aa�����,r�� a�/@:�i��as��O2c�lU�I��U�P�	l�9�뽁�hu֮o��k�͌����S����ȏ<�Z�/��Ja�m�	�w�R^��Ƈ���h��O��*AaYkѕ�n�K+#."ddZ~���P���U
!�1&X����md��n��E���s�0�hD숑�.�<(�η�[o�pXkE�}y��Hlº�҃������,GJ\'iY���i�H�$�H$" �w,B�F���F�c�d���ٙo�Y��\?��8o�K�TB��/jt+$����oNh氶�.�^(��4Z_vvbc\�b�꿻r�����:�V&�TX��O<��[I�����u�Pwvu�C4���H*�@�β����eӢ��{t�DE����"tq��V�H����#D+W�<ύn�����=u�2�"�a�g*��5���l��XZ���h��Fs3��V=��5�&i�u���%A/��ZQ��xg��_eQH���_~������RGO�(;����}l��}pv&3��ΨCD��}!1��˿��z�R�(ioU�$6JI�o�� ,�x�Ⴀ����B-�W뻿�7�m�++zn������)HI��Ͷ�o�z1ۄ	$�E"�W(]�\^l��v���z�x�7��Bec~����A�oz����>�L���,i��b����G�
f���������܎��G9 haX�`?W�vf�4]Vt��E������m�{��BF��j�+|�_�*	��QE7�:]�-�Jf^�����ǞLnہ3��2���y/�u��YYY���x�����w���I�ճ�djR���w�b���|��k�>��uEz�h	GZ�JW.(
ߋlNZG�UD	쮌����z�%�JoL��'�n����y}�vQ��Ot����� ���LHD��{�ڢUQQᢚ�s�:2u.ܲ1P�+8�J����և�ہI��}Ϭ� V�^��p�����y���{�d{+��,P]���Z~$���i�A��,�H�a`���I2���ߌ�{)5o�U	CD�Ax�������q$$$������|�iaY"���+j�����cΡ?�4�������-�n^;Wc�l�d$$��u����WH]��SU��Kx�/X��e��$�R��V��$Vx̺����5�+JJ,���;�!9�
~�;¸t�oS�V�ط ٵ_��7�^W�{ޱ��r9Y��;��"����m7��������0۩n����Lإ�E������a֕4)ug'��A���0��C#�m=���T�K�o�`���[��삂-9�\��:�J��#��Á�;팫`��e���qa��������	d���	��'�!Y�c֕(�6ʭ��O�a���ڙص�i��/�=��z���-."�IHw��߈���J��V�i��4lq�0���MZLˮ��Bt��<��Ҝsq���Cꁧh<<<�ű5]���ޯ͌��X��n���K��KFyR���.�:gJ.HiKa`Q*H��V8��RsS>�=,�1�5����2C����2����r@E-""�_�u�����Iu��f�
�,h���c-�Y�\� �ya��q�{it?�v�(��/""�k?��ؙJ��I��d&�f�`��3�`	*�&z���gP�5�k�\<SzA��)��P[�4�M(���ڹ��f�W�N�:=��=b����ɽ�uW@�&#W����x��h |�B�B�h�hEϖ��6�ӊ�Vw��l~מ��+�|k���ɾh�����
㷯���=8��>���:j6�\F�E�'�N��+�/�8M2���ޜ�4>�]�\��t��<??K-��{ +�:���xl&!;
���v�rv�2vu���=H��cÿ1�#���J��^H����&����hK�H����C��BZ��>�O�e(�ID($�6$�y�#tݫ*��X佮��y����������ǌ�N��/g���J��bRa��`*j�)x��S��L;7�J>�B0����H���^D�)��UrDx�fsC`��iR�'~�'f�X�!E��̔.��[����ph�Ϡ (
��
��E��}�~�oI#������&�xx��XeHx��B�C�tM: (���9�G� *"�� �D�_���q����Ê�5N�MM˓����T��E; �8�|�0G?�����r��)2��լ��J��hC_\�x]r�_/!ە�e,
�y"�z�� ��a����;s��R�["��#�3��q\�W}�A=�h r�5ϛ�}-�<b!��uu��>�jjj`"J�()J;�em	�X�jF
�g1���7��oݒ�,((8�N"а�I�������j;ˊ�H��M�[���y�7��{����A�ו#��q�%�y�BB��[1W������j68���b�$�*Wnx���P��zRۃxN��p���tEE�۰�3h�f���}�%R���i遲i�������w">x`I6�+�XH���U���RY�����o�V��4m׽�sD�!71��LBM��f�b;�Z�4N;��>)��x����c#�����f���G^��r[�ñeG�����E����D{Ê�A^�NN�{��F��
�}��~���XrU�|\hߍ_= E�C�����T���!&55�4ǂ"�W��Ke>�zɮ@�ghy�5���U�^���߿���+��E��s��G|^���>�~�P�@HG[�O(UՊb��Q
o��_|�|�%r��޵��y[�{B���@RR���d|�J�_�]X�������1���y�����ܓ��\��4�,a`�2�L}�?&/���B�-�K�m"bb�򚚳��f˅�E�oE=���"�cq`멃��?}r}n�K���l!�=�w�������J9�������<mj����g��OA�'�4�A��M��Fכ������,^�\�t��888�/S��S\�*���S�-v��2���gi��	"C=iih�����F&�i��5�{�a?l�0=��$�ӗ�{wZvC\���׷cZ��M����ۗ@��b8hy�)ǌ��v�_�:i����7�����	̷�9|���F������[�I�o���`��3���pT�kC���Ӕ��@�t(���0*c2�D����CSCx�9�-��I,o�tzY�l^����DF�@��s���px2��Y�ޏ��ˣ,��|�uu�AX�,�L����P\@@��4���m��a�������'(��{{{}�~��a���,�;nu�=�Tf�E��xVSظ_BCa��B����IWTRS�8��*���Z�/-�

�X���C�uSE��n˂��|�s&�,Z�K���>T�	�� �ְm7�ӻN�k����������=
����(D�:/�e�p��������t;��C\\/
�d���'�v��̯��d]��F����̅
;�51�b&��˷��d2��5��.a�~6J�;����~�<��;��+��_�9̧��K��ԃ2�����8�2� ��Q=�tɫ9����l��0�F�cfm�DZ��b1^����(��b��URP0��ס�~���:)�#���=z�����11��������@٢�U��dN�j��5|<V�U7���6����Qs�&���4t�~��Uz�ԩd 8p�~��4��կ�fM3��=��[��m���S����@�ǩsY��ϵ�7�1�9�}9�/N;+o���z��U�m�,�7Q�6�44A�Ҩ\uhn�[�h�h����������kij�B}�����Ȗ&�9߇�M�.ѭ�KC�ڠ�p�������l�����ՠ+@���b�� �V����7��0n��"��C"s7��/�X+|oݟ13�l�S��Mefn.5�拾������
KJ ��F�ꐏi,�#��(���δxE=��`���G0��l�tn��d����H�b�,2�{^7�O/���&��I�XH�f�rVeb�/����̈��^��S��E��{jJJ�s���do���@,���Ѽ,�����,6p	0[S��dT�H+���c���.�¤��l�
q�@��f��g]����Dƚ���_�~%��q"�LCE&H�]}~v��u+��{�~�B�=�qPm��5���J�[7����F�b.'ي,�gL&�G�(� ;R�Vv�/�(!ѳ�����a�~7�p�J��MN>kg�����{N��oj�=&�q�Ħgh{&��("�cɎ�~�5��l��Ɇ��U`M��K=�1�5%��U���'��~�B׽�%���r&����}|�԰�5L���%Ǻ{��Pg��$�<9+���`�q�izD,>�!X���ׯ��G��%���?56��(���C2G+�M�'���*�,D9����g�����~�ߘ}ы������tԘT��-`P��T��b�
��x����q���eB --�)�	��W$��bs0���h�L)�M�Z���宔^j���4@�5�LB�IB��E�р֌+*ᜦ���8�]
�dW��}sVf��F�y1�齭
wE:@��x,,:tk�U/w��߈�Ǡ�I�D���r����l�ѣ�{oush�zf�8��^���
���۾E\���cUK���dZe�̬�٩�Oa�e��\�!%ґI�~G��p]x<��.'''���g�F�mZ�vE�"�k�
�1d8l�FF��'�m���.C���2`P杍���=!G܊���qX��	
+�3���)%V�\��\:f��jy���e6�z�Լb?Ҙ�F �Җ���*���E���Y���ϢYBm���)�^�d��#ͥ3j�F�m����X5^���989�����f���fQ 6�45�Z[q�7�����MM��1����_���ߑ�j�j���D��m_ ��qyxx�J���Z��+	�:wvv�P?��7��	W�}q�������n�4V��_�k�]�6v|?��� '!�d`��S�`,����q�mMH�C�h`�R�B�M���LM�"SR4��������N&��I2�m<��0%��0!��n�T����f⃃���y�_\Vv`�����m����5�_M::aooo����5>���!ϓ�$0/a^ւU����D�#�j���\�]��_��7�
�K�C��v+�Ÿtbq�������J?�|�8]�mv�X/s�yx9��j�vJ<��˰�~~��av�8��S4t�|:fi� ��TTT�h(()��8�?4��Z:S��4�T3Ɔ�~�v��)x����y��� T��+G���Tׅ��7���y[C��Lq��pub��}��;�ۼ.�x}||�utt�R�[yM�J�Sl������|iOJK[(rO�d��� tC3�wt4.@�+%kT�d�&1�?
x�xx��������e/!��(~k[�v��6��H�9��DTT��C�oz�[����A.\2�=9��l]r�:�nX�b�c�g�*O�:o��� s�{N����@�g$��*���@� ��'3=�Ȣ������������v[DD���*�' @����>'�x9�&��a�񈙁A��P���xQ���K��bzVѧ#bֵh�A��)���JJJ����!����|]�F�B������iI����߁���%LP(���a�&�1%���}����䖍'։�n ����D�h�V��Ա�F�st5گ4y�1��T�a��eff�j�͑dry+I0&�cHss{zz����g�	�gkm�-��w�>��r.��Udᰗ_�����)��:т��Y"�ɷ~�k?����W�F���V������e^�Ʊ�a�"�������h[�
��
�B*����Kgq��n_��	���Jֶ� ��۱�>0�MWCC��r<��k���Ձ*�p*�>W�m�Y��\��4+���������E%�2�/~����m&�'���J�Z��gUe�O7ENNqW1���a���������k��%#$ԙ�����CFP�Q+E[e�m�����_������mk����j���·3	&�����hQ����OX�X���M��������� P��ԝ�������8��}Fl�0do4L8J�ivǉ�K
��6�Ù�����hepW��`<���$x^�@�3�����gC|,��@��؁��К��]Y���2*��i��tJ��4ҽt�twww�tKw7��-�)�ҝ�.����{��9{�=s�<3��W�f�AM#�"�U��^uD���;8L|�>5���6�17���v�%��_��&6��z��g���R�kF�����I�
�v��2A@���+H�i����җ~B.xZZ�E���t���Y`�e�~�$jee�"ocSu��ڿ���A�J��ϯ�S��eW��:/>�9<>�b��u>����L<=5������T[(���o��ڟD�#�azytt�Ԩ#�gN��V�H�����G6���G͇d���[��<�ϊ����m@"-v�X���C�Yk�Lk����Iz�a(�$f�R�v�++���{�JV��Q,��v�8s	������o;|��W�\�Vʵ���H$^k�Ȑ���d���#V8\�QK�R}j����'f4x\��|y��<#F[�'���Y�����L�Z`ya{�Q��⻁ n�j�Ck�κӣ{h���BQl�n,gP\��\�*d���w
����w����=��:4�a�,+�Kܖ��H/w6WV0ěcU�DS^h#�����LP�żF�D�!�S��m��RP��Jz��72�)K���&efz�C]onꭀ�G?�N�Y��[M�*��R�	R{RuzO���D%��i�?��	���ں|x|䈝�ȥ���֤V��]�9�X�6���KQ(�DCso�:�w	N p6����UP��Ra
��"=��i��2�ѕ�uf|!�W����:,�=����P�gHw[�¿(�`�A��+�^���yz�L�O�HLL�$�y�D�Ľ��O��A	���i�@L84>^���xp����R}��,��h<�G�f@�ӳ�XA!�v)��<�~��g�'H�Q���ql�qR��CH��*|����G:	ʂ�j�z�^`�)_�i^�.�3�O�� �%DGD����a���!ŉR
+WQ,�e�5·��S&G`��&����~�C��&'d�_�q�Y����D�q撓��ݛ�qql6:ڏ~w\�o���c<"$���O����kt�����V��~����&���܌�A�,�V�A��[�	;�/�G���
=n9��vS$H�pW���� ��Q+�3�s0��C��~ub$b�5���j�KJ6�\T�!�w0Ŋ�+b[ŕ���7!����^oa�"}p��d��������@�m�;RܥB��"	|�*����))K՚��@��v�s�Jy3���U�͖/� ��5��\����ۋq�������`���}��R����k�" �!}<)��ѭ`�c�����'.�Ɵ��V�6Ah��\
��s)`��*|��(���Z��8�߾?�k�'�K���7Xs�u9X`�\:�:��6����r�;�W�8�,��j!K�K�=�����|j����=� �_y�7�	���߯��n��+s�r?ҙ��[8�f���1=���������1M��ohi�V�%/�5�� V�v�[|g��h'�ꎘ�7�p���������,&�O��ԫ#%.v�#b�\I�E�ț�b�Q��Ң��������n,�{��f�M=-��0k)?x�\V�0j����Lf�f���]^Y�b�lR�{�:`��1�Շ	�?��S�Jڎ��c.*ڿG)m=e�D����_�^����/���*=��|�p�~u���� �'�����~P��Z�q��
	�p�=���e^�ͤ`Y2�ط����?bTRB�'О�;9%�����������!f<$�G���Lr�S��\�S�D��B�i�;ќ �WQZ߈��<2"4��"�,^o�:� �����###��r+���<̊G�����_��ύU��w�S����gD+�b����F�ϟq�6�n&{�4J�u��aa���3�8qΓ��r��g�Zz/�j�hi���!�X�0;��D���	�ۤcW}d��B���a07?�U�=��K�7,���wQ��W��w��ƌ&}��8�� ]��#+!a�����+{��zyf&	9�Xl�}�!%P9��6� of+�=mpkI���ߖ:�1���ve9�8j*{(!,'7�̄O?)Q9�����R2/�q�^.D5l2�
T�ʱ�F���}"���!�_�76����(�Ͱr����ޒ����"A9t]Ep��4Z���Ѩ ^�����	�	��+�y/�˙BT��#�=����*�.vF����*�&����/s���{A��<�&��&s�G��M�.3���[tZ��.��C��C�MMsp��4�&�P57�M�n��w�����T�L��P1<�w����W��M�f���J���>u�TH:�Bt-T��n�,����j����>��!��R^�6���SR�X@mX���;t(;��g�:<��U�:��춇Xq�VoЃ^�u��(��,I�-�E��>BjM:�B��g^��;�D�����p��EGF�@h�>O<�:�4:�sx�H�6�quw�@Uwy��@���\��Y����0$Fn!հ1AS�t>nn����$"$�/��Vn��#�㥚S��V�͞��U�-�F��$�,��dܚ�Th>��\������������S����Sޱ2'� ���(6x/��k<� T���7��V^i�F�痫"�P�/{�Y���zс:N�9U/��&}4T�_nf�Ł���p>�ąr����|�]���η�no�o�g��*��n�?3RL���h|"�u�U�p�솸�T�JԠ��voI��L��*f\\\T�I5�p�H��rf��Γ|�&k��W�:��?�<N�FN�o��t���|��v������<o(��$���,{%z^PB,��/'|�g
e��wZ�����$��[N�ß�E�)p���o�WE�caP��7��a���:�8�ٱ�w�����U��C$�]�%���|��*	�\��ёF :�(1�\���@�S�*K����
~͖8&)��ïp�R)yy��f����Po���7��p)=5��jzo�,���q�5� 	���lţ5�f��u>�#��pY��$����Ĳ)
�6caq�`4�?p�766�6%F�pWR�K*,���O�y��3I�)Z[�yN���7~�h���������n!��M��E� +�i"5H����p�혖�������������z��S&�]�QE�;��� ��qan.1tO�Ԭ��{1P��#��dy���[��޾U���=��������أD�O�a�W�F�Vs���t�y�������)�`��4d(�i��W��K2GZ�����%�k	F%l�e$�����z( -u4�b���1�2�t�RR֖k-춝s˝e`{ip�׀��i+ir��,U]ueVѹ���#���<'
�Gpz�b�o�:��\�(T�	���lߩ
�*����Ζ|s��es����t��T�J1ˎ�j��F�:��3n�u��=6���_\]zA\ZNg�4�>�O*>�tx[�T������O�i|�2�=r�����Z�5��U���[��f�b�zᕬĿ��j��3��M��;#?�����D��丅y�����jP��CI-fR([Xl_Cz/�H@����`�94��n�MS?;J�����%Z$,,�# li]j~nn����^��s����P84�_��n���(++K*�`���$�4o�bk1����wx=�j��+��O}����Ť�T���m�������ۺlnn���!�|�h?l Wq		epqѪr�'�.X0s��ܲ��*5K�������@�0AU�4�mA�#�$�$�O<2'e�Ųx��x�ݟ��a�u��Yyy#�K�tsF���u��cL�CV��Uj��d1G��O5;�5h��~J�9vn֔���rF�J���\!�|,�3S��č6ޙ��k�H�)����MMM�F�C��x�*s��EWw��vj�)����E#���u���:,�,۬�����"P�����΃����y)�8��dI���\2�:�ꍻB� �К�6jn�A�gj	s�i�[ʢ&���ck��=T"�,����5Cu�B2�����zfZb�i�]?�(�>&�n�΢��|�H���1�C"_��_8��$+��4e+��*��� ʻ��7~��\^^~����Gă=xe��	P�n*���������L���#�ᶍu�+^��ɣ#�\���g�Ҿc
K�"�+}%�4��T���*�2�ܡ��&�>uϚ����r����:n�X�]\����;�3ݣ'S�>f�+���OC�%/Xu�}�/�<X�xC&��(��1/3�����(T�"##��?w͢!J�n{���<�:�+y���l=�:|�Ju5�$�ì *���^�&�ƙa��6Y�d%�6��$Ě��ׅM�!��_Z����؅���/[�L�ӡJڬ@�8:��-6����Җ���F�s&�Rŭ?��Pc�y�
��E��k�����F%|X%��T�uM��+��y1L������&[�:�ȁ�8Zd���W��}�~I���jڏ�a��YxUkkkǼ^W/Y��I�#Ӣ*G�SE6����#��0��h5"Љ��h	S;J����ʒ�	̞��t��i���wZS�
�>K�O���l�Q�N����i��{~ç�t�d���ݬ״N��6�rt�E��}���i����X��e��e0u�w�wȸ���vEtʴ�`uH�F�E9,3ժA���>�L�&���u��s�A�7�2��H��M�#2�~>p�u��H4��0�w��d)Ao���+�.L!_��Np�_X��\Yq|����		6�|*�6/T���ݶ���(���{�Ok%�b_[�
m	��I�����R\Y�x�L`>s���T`�C<M����f�9��Y��C�I�'p�ԢO��W�?�ﱰJ��oU��,�ܵ,���%��2��U�2��jS��_�!�ϳb�@䡶*G�G	��m�k��	J����7_�Q/Y��+sv�9<֙��G�h0C��}��7���٦��998�iq��b_9U(�A�7u~��&^B��C,�Le����M��t� �U-5fT��!,���$r��R�ʾ^���Tv��6��guh8~�����%�b���?�˔2a�}��y��o츮��#����i�T�?GD������9#���8zA���oƅ��Ͳ��m�Y,K���A�����!��c��f��(������M��Ё��` �,	��R�Ԃ�<����9�x
+���c??dF4�ԇ�s��Kj���p�D��ݔ��̼J**���e���g<uf�W&�[��#�Z�ކ�T�]�4�6GFdX�mXI����01�o��võ2�<�g��]>`�8/rQ�nUsF��D^2S�|CW��1!�j,��p� S��'s�>�w�!��+�j���mS:-��k�c���Ó��O/��(�ߎ���~u|A��8����5��i{�t|�
�v�e�= n׳�;v�����p�dlr����,���B
��V�U~2 �����n�?}�[M��i�]�YOO��)���ĉV$R����IlE;ܐ(�� W~'ʌ['%�[�q��v�s��e�=�� n�j������X躱Q!��/q�oj��Po��q�Q�bB����MMف���1�?h��>Q�`l��h~D!�Wa�e������c�ҥ.����j���ؓ��3�����!�����Bgd�����U�Q�>�����S���^&��X��|���*�B���U/.s�LW,���.f����H{�lJ�7'����,�����D����Q����؛�@�1��Y�{<C�;�⁞�Ꮆ6^�o�.��/1�\���0/Mu�W��\J��c�F�
Q|uY��ۀ�l^5�J2�N���`��q��� �PU���AF�~OqlhT��h��Ov��S�?aԩ�>�n��S��2��uI������K-�����o�?��b�T���4���y��#h8;p4�����t��}�C/�)�����wd��UtΟ���g�Q1&F	�ҮZ8w㡘6˛z���D��AC�bP�H2�k�����(��xhh���܎�ۇ6m5���nHkP趰��h����Y��{��D�-�����n�� ��h{ee�����j��	���Q^,##�k:���n�q{9R� �.`if�.M�w4�ҹ�a����b[m���$c W��M1D`�}g��nX]'��G+�s��
|���mk� ��Z��J��b��hKH��Q�a�1�hɃQ	���7'k/^�(v�kB;H���]��Bɣ̎���*�OMykt��� �����r���5���O_���ۤ�8����c�Aݱ-qt
��l����|�сM�z�~l�x�az����1A������$R��7gQ!>���7K��dr��)���zt��_a.`1B�%?b�����D��*M�Q���zA���m�I@EA2��w�DT��Zq�ZS�j��AR�� Q$>~��|h�F��FS��4h���¶9��xJ���#9H��'x��Y��^WII��W�����[�V��z������[ �X	 ����i2�d̉����'����d���'���6�����~���;��6�?�@Y���v��]��s�*�J�b���)�$&Q�"{��U3zx=���4��k`j8�ڧ�D��|����Eădا]�EZO�@�9��������q^c�*����F�e�R��H��5������m��n.��kn��n%�ӫ���:C��J-��ߣ)�8�.�2�POiˌ����[�ba�A͞�Z����7'��B(�P�j;�Ӛ=��� u�v[���S��ҭ�A�f���x2�N4""��������H�96{cl�X���S��r����*���D�V��(�^g�O!jw�=��?����ǀW2���J!�*��4�b�,�h�6d��p���ÓbQ&f\z
����D����wյ��K{���p7���L�e�6�O�t*�R�9_i")�>��N��Oj�iX϶���Z��f؟��ȁ�n\��ǈx]ϒt^^�@���Q&�7Rͤ7LV�T?-�t���cP��|_���/�78�:����_Sy I�7�L��xb@���iޣ�&��w?S�8�)WϾP����Z`/+���y��m��W$��MT��V�	?���x\U\F@�����x	�+@W�0ϑrttb��C�N�������i���c�����-kmj����C�)p9Z�1��;Wv����#0mgYt�fKoX{����T��be������	�y��%�����d��z ����6��ek��?�I�#��J�EXn��9�rssg�6k��֪`F�x|�)D���F&e���ʑYr�p�H���ˉ೥���xFi畫�3wb�׃�0��<i,�R�Hd�=��o�l�8oV3��䟓�@�ό� eYYY����%�2�_y�2
T�q�Ғ9���F�,��IF<acx�rE�W+xѼg��yW9?�����p7$}�>��o9zw�`�`���z%	ƑGS;��awO����_���Q�TfS;1�+��5��\�(��H>p|�a�jQ��9S��7�hGC���IR���B˺�~�6�7�����prY���N�[��K+F�� ��ӎ��[b�rbY6+.I*���k�q@ �|�	���v��v�L��F�����\:�y��4��}M#Ae�x����q��#⑃n�*��G7v�E��A�H
���<[�@�����'�7E�A��y���z�v\�P���qS)�= <�1��2���W��:�o�$�j�1�C�a�~
Z"o�<��7���$�/�x!�#�@��F�D!��S���. T�P������ٳA4_�3ذٕ��;�T���sU�-T3�X�yǘ��{z� ��o�(�c��b߉KK#>������b$%&:=�
�=1�����+W�_�¡����V�K�K�A�b���v�+܇�Zj�֙N��z߶�u��q�]c�M'�F^�\����p��-'��唍�0��X��Ml��d[��~��Oꡪ��֓���g��������}���KJ���� �i��ZT���r*���B&umj1)On$�Jt6�h:�֖n�<��-u�Q��D07� b�����<w�3��>�r�!!'R�L��:�����Mw3��;ҟ.�49��\(Wc=Ka] 0���0K�P:�c`��K�E].��Ψb���um'���C�"�
�5��ݫ��|]'UP驪Q���F��y�N]���ި��������JI����TL�W��a�V��k�#I��nZ87�����U��;�[������7�a��-�.� Z�&�wtm
,�^�;Ȃl��y�:`N�C����U#@£{p� R�>⢗�x��8���5���B���}��l1_~n��zjٕ�=��CJ��P�d�������\gZ�pc�a��1�5����եW}���bnK�R��e(��QQI)�8z0tp�~����Ol��2'A.��{7��?�R�A��>>�i�2
��{8~��AI���ذ�=���A��"��^��#��1���C��G?���N�Z���/!�8�B�#�V��	�+�QE�^W. ��׫��`�������8��W�o �Ov73 A�����5��B#Y�!��"}�v�o�CNr�HjTe�>���P��I\�^���r��y�9*Z�#>I�c_i�y���]�Md�ΜP�K��(�|5F2�>�v�t�N1��P&�6|h��=�?�A�*���O�啕�J��\��і�x���i�@}��^�G/���vvv��p���Z��ZM^��6i�P���͓[~w�lt��w�@z�D���Մ־@�ՖA���Pܿ��̏��m��~�<��eE�U�t������H
����PH�
ju�Ta޽�U���w�Ӫ ��e�UQ �չL�K��m���ٰK4���ӫ	D%���u��$�����N[+Y����r�<��~�d��� �a�W���w�ǁC)N��P��~���B���3�������&�H��X�����+.HfFωn~O�8 +C�[��.����w�!m���	���s����^5�ϡ�Kݺ
�1��E���r�f�䕔�o����ͯ��~���GZ�L@bJ�?�x}�Z�.�x��J*J��R�ۧ��P������RưYh^�'z�&u�/��3!(�H/��p��j�����{����@��}�Xp������n������*s�v��!l���y~
x>�X����2�=Ysy�i�̐,C��;x./G�@���dtۘ��5Ư֣&$�~��#��EX��X ���{�8B��W�ݙs^U�VLB@�@M������P�$�̏���+��do(��Kgse�f�M6|���Lc��6�B�t��baHE��h촵�����䦥�fH�=�=d��u55v3�ۍ��Tj4NÁ�5������(Tc�-l�f��a���F&��N]@g���@�)�k��={
��^v�����/6������&	�����umT>O��,�#�ŲV���aК�*qM���@�!q%����=�,�F����q��SPF>�w�n^�Tt}�0�#������)��P6�.��1��>LhD���u���n���ޟ���];F�&�m�铵V0
�D-R�b�y�I$}QV����|
mr�$݀�v0n��ԁ�@ŷB���*yx�(���P�2�}[��#�۬4��y=����x ���g��ʸr�<�����`�y��lh��J�a_���1:�!`Rc���m��zQMl�Z��$�v�+RO�N�⠤rK�O�[oMW����<,�љt��>>.'@d0��t�inn�*<��J�V�Qqy9�@?M������ǫ'ũFe�@���_��{`��d����kA]��"��×�S(��,;�c����������
�µ߮{���L�z� XV�*�O��&�nK�s�����+:;:��yܞt�mEr�sp����=�g���-	�e�K�)=p�	�{�hv���Ô�{�hٵ�9Z�Vo4�t
�����L��*A����������]D
W��W<]KS��1��njW<������L���+�|D�w"2m����.,���w\�̃�i�|qPO�>�#^�>�P,*��a��1w�B]4�����[E��JT�Vs���G��,q����̨���tMn���'fNI���+�P��O�d*��L.`�F>�|yv����!9?���w^RRR۠������%�/e,�U�Q$��7��oe2��VDP����������_��	_������� *&�Q.�i�Qg*�jC��M[�Қ�O�`��6��ʰ�p�J����L �G߰յQ�ujt��I��ҟ���� ����r��t8�B¯)8�<-��%�5�������0�&::��O畋ϭu�bA�x�x:׷v0HP��S�-
�.�pc)��p�,�7�����v �
�07ׯ[�1�)�6����k��1�ע7��$T'+�,����IB>�G�Z�G)D����Q��#�ю�?�YKKA�fT*��z�45|��C� 0f��v�@�::����GGH���8�{ݮI6���TL;�� �=�l���٤�Z��z�)��l�J'��F�� �!	P�!��/�'E\TU�jL>d�rG�⫚���^�\�0s¤�k� ����&_�Ev��	/��������gB�Kc���N�i(�wP�װ�X)J����S����R���-He���*�@e�{=h��m�,8��%~��4$�,�pP�m��]���g����z��J����m#t�t*���=�|�@�@�cB��u5�B!F��)��Ěp!�_?nQIE� XnIV���^���v�G`��|_��񒠷�󼭉��,_�-���ݿ���:����xрò}����\!�������@f��2�s<G>!2eL��y�^&	4޴UŐ���/H{7�ΪZ^&�3O��?y��Ӹ��������&*��O_�2S�U�d��B{.P9����lk[}Ӝ�cö������o������7���9���Р��,��[��p�"��-�Xs���\-��vCu�_���E-1?yg�5�nS�2��e�,2&�(��E�	�WQQ���q���	��t>�w�1����� K.�`���e�^��F�C�g�^��{��r�]?ӪM��|h���ݒ�Ǻ��<����
�PN���**ɭ?~Ï�?"�ONJj�Ly0�K9�<�HJ�q�y�oQ���8:��(�|8��=�9�%��E�d�}��6Qx =�9 ��'���Z�VP`d�������������lS�p�*�}2'Ϳ;���y�g��K�����r����]�p�vV������s��+��2�5;0щ�OP<�ԛ�	�K��))�X��ϭ�Y�"!�zx̪�J8�x�Ng
e=��ڸMAGg���U�`q����+�oɝ&;�J8tz�����z%�4俒�|�Q�ӾU˙;C�J5��P�ln��U� �	Bc��S�ҏ,S����022�c>�LtV�>J��:_퇵���*|Jm2�	:�]up�X�Y��e�/�Ϫ�|k�%�d�ey=����~�9�W�'b�����>�'*�q�y� 88� 22R#�K�G����D���ztF��jђ�G9�lïd[K�w���D��to���gd�UHN����Si,����u䞓�و�QW��ϲ���z��[�?AV\�t	�E(lK�)u*]�xh����Rb��ו���qv:|-�ݨ�ߋ"�Y���m��w|��.̮a�Z���=�w��ǜh��iY��7��l���L����g]Ki6)����&��z,�����$3�ι;�GG >�+��l�ı$]��ա=���DWH4���1�R&��2Q��������ԉ�9'6��0�=A���g�@��}0P�I�%�~�[$ئ˙S~dt��½,�_�%x��u6��0�bɋ��J ��k��j0��������(G0�C�T�I��t��K�;֦��_44�#���AL�I��U�Y^1���ƣ��|(,��@��
���41%8��|���t�����.��s��JS�5<:�{����O����cs����h�$�ruu���! �{'�&b��߿C,���mQc�޹��ר
X�\�e���,�l�lxq�'7����Y�i�J��Be��|Q������M�nʯ0��XH��1_,������Vt_J���3n�\6�������U���>�C;����P�Я��6���0��u�R�x�9�=�a%�x�&�B6�!v�$� �V�I�8o[۱���`�R(��ɕ���oEd��C2`W��u*8�R Jc0���Y�#ĥ0�B�kU��9-h��l�7�2���xߏ�̓��ڋ����@���fw_�R��Ӻ��T�ZX��uN{�6����.�&6��~�H^���hQ�J�-V]_9	!T0�GelY��S�v��;z�v졠��ґ����0�y[��K�b= c �*�,��8V,��ɪ���ך�M���aU'���|���n K�����aٶ	��
=N|>F�;�H�I�âAtA�.�)IY���g��诊��j�z>���Մ0�n������¥�9��1*�N�U2e��G�Cj}�3���u&j��W���_�'�v i�3�E��8O�I����m=L� ���|8�^vNNW����H��Yk<� �!Q
��X�[!O�Q����"(�?��o�X�ayjj���2����/�P�9����p���e0���B�0j�49�B���x!�R3�2�K�g��`�RD>�@�f�|��Y�5yg�!�4ӱ�'(�f������:?�lع
�����\۴�Èmp�,����V�^VR���a��1 ~8��T@�O��:�c9���l?�,/�A��dә��3��<�A:U�#+����ICu�w��---��hl����#ׇ�kk [f܄���r����#��~����<!-td�8��O���~�S��/�[d2ekw�.��T�#�%ژ���c	4��O1l�����S������fn��z�ݶcY�W��	!��?ob�uӉ�1���|�/�-*�>a����g���6I���ʈ~5����y���������U�� ��i4X6[�ǖ���gۭ�I��,4��KKRL:S�W�;XX�6�w9����,T	vp���J���F��w+u�4����_�a�߇;�=<<�Fm@J�w[ؘ��6_�k�d�]<C6h������0����Z��r���>we@�U��4�P��!yP!%H���d>i��vq� ��w�����:r� �-�;����&����+5����Z��G�9�b�����Fؐ�'a�1@X�1�w�����%جn�S3l�L� �з���G�xF�lz����:˴E��k��m˅�YMbv��(<V�6��cE--�W�g�*޿�ԅ�����,��7ɻ{��nQ��H�[�4����
�MR$�M������D=㷜ۓqus��N�Gnˈ��lf2�X������RMB�fi��f�_牀���7�I��hr��߮��x-��ٌ���&�;O_C��l�aK�)��x�3����.�N���mZM�~0��Հ�3��/8"�ţV�U��HW�YԂ'Д�E����l��b���u���7gn�_�ٟ��v<���:����a�(5����_����Hc�q]�0.
�"���>j��rc�M�(M-�~�bz!(=oBe�h)B�3��i���|���w�C�C�MO;���2TH���J�'O�xVr�Z���G�g��cP���Gk|<aF��?�omx4��^��a�MIeJ����]�t�'�0��K��9N����\ߝ�AL .Y���-~䲷O��U�`�?��G��F˓·���Ưl�&��"���,����c��#�� "�(ă��T��{td�Q&�*z22�s�Wڋd��������p`�<�  ܠ���VbAv��n���+-?���[�7OuMԮ�w�����I��L݋vl��a�=f�D��Cq�5f�-�����I��`�o�[q��5�M�uj��,D7Jr��"�1��a���*�`{ "�x]y���W�ie�+Mz�G����k��$Z޺���PC3��Ţ��U��x��x�py-;��C��`�8B>\��C!�i=s�e	O&}����?;�K��!E)*->53�wk����q��M=M�	N����f�~�1����.ߞ�f66|,44V�����>�+
��*����2Ꮝ6��%��u��:�ˇ��A�'�;�wc���G�j���gNj�[����Z�����Fv�Q��v�hq<�A+#S!��!��:�}ۖڀ�e���p���a�<A�ua�Q'8QZX�PI�8��n>'O*
��"���������i�=��Y�(��=��k}��L<�4&�O�֛׫ֻp������1Lj)�73+����?��W_�-�Ev|TD��)��x*Y�z�n"�r�ftr�j,��`tņ�5���O�p���̮��k�h�.mz������l����S�q���y��i�|�~r��P�Z:ZؑQ:�Ƕ�Ⱥ��:-�v�}B��d����7�OL �t�M94���̶�3��)�sl*q��T+-�w���S<�v'M���������Z���G8↶=�yy�1��/����k���vu$������*�<3>Q���x�oz��co	�!_�v��˞�͵��5'�"Վ'��cv����,�\�ěv;A�N��:}�_����צ֍9e���+xb�q����H<�bŉ� o]tN�tE��W�.����!ZYYm�)������cޔf�;o3Q�q��~`��o�F1Q�s���'&$L��F���X`�u}._8LS��^���hf�����G�A�����5&[(�;?�ifZi���B5�&0�=��᩟b��X� �|���~c�����)G��J��7{niI��nk����y����/Li��������H��y�ܺ~�U��WiN՘zbB������(�KZ�����fяN%vԋ;;;���l�,i�
Lg��Y->.�-����5覱���d�9��BW�B�tL�����6VV��`�t����BnT��0m�[UJ��L�!9y�\�ԹLR�^��4�ih�)�w[OG�*E���L���l#L���m��m��#'�=��O�$��Wk����k�-!cTw�BkA)n�����KkK"��k#a�w�F\\�=�7���J�#l\*���_M����6e�`��w�=�ǚ"�GS���L�m
4���]�d�̨퐚@J�`UK���(B~
�g�Ω�5�U�FP�!@$�V��y�ٱ�܂����#�A�%���^�����f�fM}S4���D�Q'�i�����X�177�$���CϨ����Y9PʸZ�W�����XR�}����9�xy�=P�.���r8����c/Vc��j&�)i���|+�0m�����~\���m�S3�z��R��̪�>x�p�k�6��dm�Բ��z��t4>m����l��f{�����k��?xF� �ozVv}p�K����"��@�.�|~����٩)��0[7�uϘ����_����~���v�v�g�3��9*F�;h�$k�����������>yf���vgI��3��ƿ��}�#�Ǥbʧ�18ħc@U��� ��2)	�<��kZ����.��J�z�C�<�I	{���o��B(z�)��П,x���*U�H��@�$����s{f#�(���=�L���O֬f22��*��0���p�oM�Č��r����(�|��CE�&T�R��ْK��E ��[Rh�4�;�w>�X	��� m҃�H�OЬ�)��μ�̡��fb���Φ=N�g������V߄iJN�H�����]�u>�u�_�9��3E�B
�~"􋘫X[[�٘��F� ���7֗c�K<�v5���4s�%�V�]�,�����U�t��	�s熈T���b�}���l��&���?���2)�>�p���i�!̫��6��I��G2/��:d�#��h�C�1U�]m��:^i=u�ƫy;L B�K'|�7j���+�"���TŎ�.���6y�_܃}kY^e.c2���1daEuus�Ub�Ȁ�+&�h~����U`���}2ˎ�΍IG·K$Fz��}C���.x��ֶ�o�?a�=u�z��NH߮ۏ2������_n��nϛ�g``�Ī��i���_)õ�W�.�������>[�Ie��q�'M�*w���Z�=���׺J�|B�����s<L���?3��8�צ��u�n���׾��z]���̔qXG�ǿ��=n���7���P_B��5��i��D�:�g@E���a�q>�뇴�Md	��E�xf>7�2�c�(L�������~��Hu$=�|�c�k@�:62�!#d��L�����i�JID�E@����j?������� h�`[�!F)�M^K'����%A�TƦx]1�o��Tn�3�ȷ�n�'�^ը-�k���rbz0��ӝ����$��JH�,&&��ܺ:�O��/i��T�����QX\�����ܻ�������Q��[XX\�>�&ը�ѧs��KW�H�ۅ�M��}���1\\����Lwwww7����\��15������	�}�s��ԋ'*݉���@�vu.�<���.>rrwwW�_m��:j�3���6��%�Rc��[k^��Q&c���I	�	�l4O$ y߈1�G$�B�� �E�� �U�aXx�4���A��Z3�r|u��b�e�8�"?�}���5?CXoU�w�5�BFFF�)�"TO{��}�϶�<5vZ��:�|yWt��P���8��hq`��ǝ2��:��-L�[�z����'��	�����9 L��*�z�	�2]v���+Lf��m�!~�֔�z�
�AZ�r�:�W�&�C??>�/kuM&6��{���������_<O~D���HƓV�w�M�"��)i�f�M������|Ge@��G�{zv�B��*�,�E]V�S�u^"��?��)q�f��f�8�`p�;�*2����Ɗ���	I4� x�,��qϊ� ��p.��5��ǪX\Z��Z."⻞�sa����i���K�����~AIC���.~�(T��|�fm}� H>0sg��_k
2� ^Y.�z ����wl|��5.�F�{K#*-k��~k�-3{%Ӳ{��,v@�ȵ����I��K�����4�0
j�F�w&��x!)(&W���44�N('��C)a�����Z���E���Df��(9Bc(�I`M�A}�%�D1�Mdwޝ/H����.�/�.��p���K�qȉ4��ʔ��98�jnkó����?��b2��-lq���s���.��u]/^����� 5*Zx�E���Z����/��<����ǝm
������^�k�j.����4(�^�(G����z_,��>b�PA>��6؆u���O�*�n��F�n�㆐'�^����2:�F�7�?()%�|����<L^��g��G2C��8gwڊ���?�{�Ͻ�x!�#%.�vp�>���ڝ��6�[�����&G�'��8B�$���{H>[�a9TH���n�6��d��i@�2���{�p�N�"��=�D�Ֆ���3�c)3��doJ�t�<B��ll�bE3�6'q���0�F��c��$�X�x�����[�L<�ڥ
z�������g(�����>M�Z���x��^|��������՚�p���_n�XI)��{����(QAA������C(P�#,zj�!Nk)���(|�ųN����� �HC_�=�̶�1���Y��XB����o/��oz{P�����$�..��Ӆ秂Gd ��h�.B!i��)�E��تǺ~u+U�Fo�6�{�-�(�2ӆӬ5@��[98����%�	e�t����(:�T~�Lyz=I����3�b�.��`d~l�U䥡�����a�ա��=���^���`���!7��`�VI�t�?)�!U�%��y��s#���[v������\��M��m)�_|Ae� f�l	%�]����	3��`��9u�@d����:0�����{D;g�ycB��]���T��n�^6���(�Hu��{�	;a���L�ٵJ)������VC]�.�wIc�?��S��?đ��lʳxVz��!�6؉|�Ǉ��B��N]5�˅�Uz��A����d���t����AQmw{��d�7,;����r{��^i�KL9��Z.�q�/-��!�!�����֬r�Y��S��s63�^?�N��.Hmy�XI1���1�+d���-���VkD�!$Ud���E~J-�Y�����q7P�����ё]�׿��W_�܍m1��9� :2�eo�V@���O���Y+����N�d}j�G}4A�2���X���>'���&B��b�6)yѧXM6�>�:�!���]g��l�K�_�Y��u>�ߓ�Ib �oǉ�1�j�$1d�+���4b8l�|[QfD���I,_��q��h���ߺQ{d�Jrf���1�i!�XW
��f���-�糬����ʛ�(�������]�(������#ES�}��� �n<�ܜ����
���s"B���HYTs�:-�,2����A���5�w�%گ�J����B}Mm>�'!s��.���O�8M-�b�k[�����l��2�,iB��h�B��`�bB��=�d����u77�ܻ�#����V(�+2��E����`��8�����P����U�h�ߙ3	�y�yWzf���:�A��m���*�2mRKY��j+Τ�y���7�SSϻ�/Ӻ������ *_��r@�.����m9%=���J��Ck���1{�1�W4y�QڙK��S�^y��?ƍ(A>�ncؐ�}�nT]l�E\Gt���!I�%J���I%]�~�� ��Z�@C�v|b�/y���O�U=W���\�J7NF��ks�@(�?��B�P:� b���V���z�!�o�[8��h������U���B����}4l��a�i�m<�����ei��wJ`�G�+�dd��::>�k���� &��������'1��e~�E2�M�ùM:���������攽O7��7.�2�te�ò�0��ҩ^lv-�Hn�/ݢ�����W�^��a7��F����^ ��QX#5�z8A���z�u6�g��BQVH� h�Սmhp;e���f��$�֤�l�ek*G8���S]}�B��c��=&)���v�z���Ζ���^J�8��=ڠ��QS3�_֢L�1�Y��#{����56����LuS���n��ѭ���b-�(/��$H>_hJUy9����|���l��*��+���'_+��Ta�wI1���\&���T�b�J�"�W�O6!4q�-o��n?�[�ɠ��bu�א�m�=��^�ZF��$Gc]�Jkȓ�Բ����/�r�/�;U台��N��1��5�������al����m�ʍu���e�Sv<^����1��L�('
���:��:^m�ī��.�lvs�iw��P�F�uۻ�9��5B��o߭0��_�u�����*����ҵ:��4�C�s�HV�.�!ZE���"Ȝ"f-��Ȉ�������0!$@؈Q*�_��/O|�*��PhA����`�<@��kͽ�B���.��EiT(��~:Ru2���Z(Sh�o5$�iqhԉ�#��>Y����rJ �R�Qr0Xg\.��m+s�;t�~z��Ǒ!�1�I��K&�,rz�w���M0s`ӌ/��o@�=F&���Bωwx�Y�ud�_{����"
$�]������[f 9{��
��g�����Ģ�0֑����I4����J���`��j/�-UI)����aɋC���1�0E�Y+�d�D��QL"
��Z�
�҉w�o��!6+��<n�#Ŕ�.$f��]���
��^W+�|���g�������/��WD�M��ذYT�ue���}�*h��y3��E��F��P
��7��[\rr��DL���o倫����ql����Ö�(!����Vj]��fՃTl��͡�'�鴚�)n�pRe��v5J@++1�:;ehĘ4	n*��&�<)���W7t#�=+?�����"��P���¸7�hdfƌ�phd���Y��cq�h�ٳ�(�F�%���9���P��={M����sm�ؙ'�=������0��E���C�l���;�7㻥�Z'Aj�eG�J%4�D��I�f��|w�v
_����O���TVZ�8���8���j��ZZ��);�8��ƙ�yc5nqs3�(b�껴Bi�av�l�JqJj[�FF�T�Z��n`ם>��ᬸ����KU�֖���r �� ��a�
�BV�-��
��WS�
���?�a�ՠq-�?B|i�j���~�}z24w�ւ��TD (���.����`��{����+6r�^�hY�����wY�3
д��6�^��z��L�N7��._��$	�b��q�Bmlm�/�o�Q�Q_.�kmj��k�TT�"d��X+<RI+��N��+̫+J�a�=��%�K�B�J^^^�J��@�w]���L�b�ގ��T�HY�|�IB���䪚�^�cU�zSRcf��)�E�Z[��|f�� ʼ�c`e�4W��)�sfc�m	����f����%'�A[�s!�	�b �{�
�����ʠɕ�� s�k!�AҶ>����br�r�U��3�Cd�<�= ���;�B��OְeFG���Z𑰝��R�(���i!�^Ŀ�6�~�hڜ(^B�z��}����Θ4aB��6�� ��n����/x�!V�C���[gH�lf�p?yB�])#��%�0A�1�9������ʔ���{%C�s3q��v��r�<.�9`���.b����d)jh��T\o1�Op��Z*�[Ԟ�hhn��v"�C�t� C	K[W�vg����]��v����i�֜T�&sCG����]�#�Ԭ���)a-� $HHǟ�A~$U�Z�~�:�G�mܮ��������E�Ӊ����b�PSu@Euee#�ӟ�];'��[��6�T41D8����V=�GF� ��Yu��k�Os�Oe���v���{�(�D=�׏��{^|��B� �re��>a�~ �X-DEQ1!U��)��W��M����Gu��ΜJ9a+;��<ޑ�L�o��P"�'�9�]��ҍƒ?n�<-	
�}�Y104�&v~u�_J)0�d����}�M{�`��T2�7�NR���f�x(�9o�`TC�q�
I�'꧸9%�PY���n~��y�ߪ�$�::X�C���"��7俚��9l�oY�p
����<D�b"|�!���J唪a��b]hİ? �ެNs�`��Ϫ:Q�͔���Q0O.liÝu�Ԡ�!OP"�����q��	_xm���C�M�W�M�}��x�FH�Ve���f��z3hm�� aVa;��������*���x����A��OV,&�H-;h�C�����BX{����H�&B�h��ƌS\Z:	¬INV�j��I� !����~���V���Ȇ��v�F����F�wiO�������m�v8�p\� ?�����ä39;����������	�Q�ڔ����&�6���2`w�2P��z�������"��[T*��y�	v��V��N��xӿiLW���h�,��G���8?GpY;P����X��v�6���ȁ
_�
��2R�W�]|/
��Z6h̻����� ç�ha�p��p��M�N���=�֏��-�[㢢Eߠ �ݗd����ꙭ �qċ���Q\�'�яd\��=�W_S���yyyiVzhp�,�CL�93y!JAZE2��yxKT����Z|��_�L�א0$������!�:+K驡�N�"�Z��=*��wAۥZ�W�������h�bpw"ñ�F�:6��|zXl�B�7��k��(��f�&��gW����=��H����}����$���8gZ:k(��� �U
��>���脗��+tm�7��=�rJ�3�� ���-�h��p� ���jto��W,Ks����<N`M����:��w����K���~������w�C�gwۘ������h�]��f�J�R������6��X���)��]"v��@�a�.c��',|������R���Z������O���ț�lw	q�07������B���(�92���d�@�յҷ�0Y����<ILE�띬�+�f�i�p9}ܷ�9�߼�(�kȴR�EVyQ�0�����j���au�f[f��v��-ć��t����sX5uuiͽVf3�=>˟�S���`bj�Ze�EP����O�2�50����V�7?����q`EEίu��gX������_�$�,3h�����J�	�ʚ�j�y��}��,p>�}G�e$QO�2�������)C�T��[�}uAt����MB�x(Z�K�ȵ�Pu7��y������!0���XR;�d詳��g��"��y��-߲�;:������Q��c��&w�lm�+Ɇ��a��*�]���*9�sUm��xM�I��3`eu	M�]j+�{��%�d0{��]̧0��>�p	j��;G��Ë8g�6�^{Z���:��/&-huj��fǨ��ˈ�	)�\�����U%�w��ȐX����K�7S5�Ƽ'aV��b��0�x�����Q�נ�k��6���.�����|�!a?�Տ�s`'��@M�>��eh�l���t�k�;�W�0�������Q�N���{�w�'�L�
G�(����	KW#��寫Ƶ{�e���S�hZ��H	i�rЀ`4Gî*����~����Q�/���jˏ�S�q�t�"5+e��8�egw�_o�
!�Ć�>QG�Y<�>��9H�9��Wp�z{��4�"|��gx1/{5ρ��]�͗B��X{Gǀ��ۿ%�������u����z����6��_t�T�a��T�=��.�O��JR����Ē~PQ��P�s#|�W��pB��s��8�}��	�Ϝ��#(�Z,��j����!/y9�������K*��@ԾF��w�l��֨D3H뜃*�6��x��¹O����:,�22N��#sE͵F�ue���!��V4�(U�C��2����70z~(��4����a��vd�a�%�.,p���{<~�x~b49RW�>wB�'3ÿO��������)�	������f=p�]���[;I^��Ǫ0@r�
y�[��B���σ��ާ^�QZe���u������3X�ԵԴ�b@����E!��~
Ok�o�6/˩	r��U(�6������"OD�Y���\F��<�%%�ﵞ$,��=U��ձ~G'��Q��am[4|~$�@NO�t�/k��0[KҖ���\�N�'�wW���Du�d0�c������ut�45oиK|Df�+�z�X�K�	b���=�~;PU��g|g���U\??bƬ_#~ݞ9|�`~��c�5j��
D:/7��P���Y5�u��]��L��	@�9%�_h�d<i��aM�O����Ab��a��&F���au\N�f*>R�}���x
a�dS����?(0D_�|d"����j�GL��h:���^�}ӿ�7oRh�k�.�����ŉ�lb+,�7�)|�P��+�;���i�[�K��x�9Ɨ7��T����\�.w{6|_�Z.�r.ie�n��1�Ժ)�{3mA��B�LM�4/0%���e�"���I��cT*Q�I^`Z���%��NmF��hQ�d!;/����Yjw!�Ҥe5�β?��D�,4v^.Y�bUf�k�/(P���N>�K(z���/�p�0��V��Q80��n�R5��5�
 _��,"�?۸�=}����j���}�Q@=�:(d��#����"�l����n�o������t�~C)����;(�,��L��(P�S������Y�P�牾�	���� ��{�c�2�ww�v��^�uu�=�a�
�#��������M�&X�U���0MsCK)����?�M���Ωi�v��	��K��������E�2"c\f��\��e�0$���q�J#�M��F:�wjkҍ-��%��Aj)J�0��h#ZTW���R���ʥv8R�2(	P��c�|�!c@wS�I3n�|1�3���]"���u!�k])�$�:�T��83��c�F�2���n}�|��Y #Cp*m�����F����e�M�5��39�R�$Gs�.|�m qiB �))�'R��K�����<z$�s���v}�9[��J���r�k����p�Ģ�,�0����ĝK7ߋL��Tu��^Zr)plX�V�l\83#Sc��f�?wt�V��I�����
�����1:����L�:�.�����Ѡ)C��N#�S"����hN�DJ�%GD>O���A�
`�G�ƈ��1S�z���9��$8��d�YǤ�g����P;�c��|K�
7wk\B:�ڪ���p|Bf��u���c�|D1��̿�
<ъ����,����MX��mn�n}����;%0�|Z�<���̂EE�qm����ɛ�>S^�9�3%��fH�4����km�R!��8�#�����[�ڕ���Ly��د4�[.ߥ�Z�����Q����#GFHXyv���x�����P��TZ�:P��Z�66���Du�gd�������
/��OQ������1����MA�ӣ��XScu�*_�Y�g��`�9s��r��0���QnL^���z�4���:��қښK�\��A;�I$QD{����ţS\;+O�Zfɱƞƺ���N��B��b�_���&�_m�Y���W�B��td����-� E$�˞x�_=MM�S�=��tL��,MC�K��bYY���Q�uv��m�S �D�E�^xv�ȓD�ߑ#�	�=�V�|��l6�5 C�]"�������8�/x_r�wO��,�u��Y�$�d�-�*&R�[y�*2<��
u��̜G�@��շ�:����e�75o�LZ�g��LN�R[�d��-[�*R3�y`���ѭ�7���2��ݗ'���SF/.m���J_\^K&��ϳ02��Yݟ�s�|�o1�Ǝ�=|�e�d�d���E�_orf2M	̩(�8�cY.�B9��v��LsXM@��v�����|j��'~h�(<�p7d�^!ZEv�oSm?�xx�?[]XX�081"T�BFP(�]H�?�΢N�H��8:ߦ�$;��g?1��P�_���	6h���;!�l'� �̀�c���%�,Ns�V$^��~���d�.Z��K�R-��i�^�|�T #>�E��/�E�KoF-^7���K����b�Ԍ4����r���%�BK��+�q7D���ٗ�G��p�ϰɌO�N���dd����E��!W�Te:��$L���t��2��B�6+W�����ʽ��;[AS�U�V:(�gPlZll�b�@�~����z�����ŵ��!�W��'w���Ce�+�P�P�����(����%�a��QXǄ\̞�rEj�^��@���D�+F6�Q!�1Ck�r�B �}}���qԵ���ӘTtWx�������rsH{V�t
x��Ls�c�Yl\�\�^U�:[�C���_�_�K�M���~
��(gn�̽S��M`�V��6Bn���|��3�f�� q���DG/΃`f㊭�����W�p�~x��;bC��!�en�'+[�O���X]��π��ᰵ~��211����$��|p	MKK9��5D�dJ`�ЫQ15F̀�OJ��Y�NO՚��$�
�|�����vU!�{[$��-5&9����8��i�#��3�8� ���tt�������<(�^�h��WKN|h&�����"@�E����5=�H� �o=tu,��/������FA9�s�18;�\�2Y�d����"s"�2tV@�/ڏi?GYW���l{������|T�(�u�tB������TN��4ln*�j�,����/F���Z�w��v!�d9t�	�C�q��rL��n��+��@5J�Vk ��p����[K�����ݫ��O�CŢC?y���㙕Օ�C jD~=~�
�Va�L֕[�7���2�'�40�������P;�'"cz�G�W�eҩ�mlQ�L{��O�Q�������^(�ː�����������Ru�`���p� dѺi*���*':�9M�ؓ''��^��`�� ���v+�b�N��7��Q�(�?���(G_־�b�^H�.�Uۼ����;����R�M�%�A'Z6��Ӛ'�6���j�ri+H�
�f�74}1��%����<�www#���13RO5�43e���S%��	O��1 �� �/�!�'�$2cƤ�΢�h��l�J�?T��	��QTZv���D�r[��� Ȧ!�yrD[ _m���1��@�o��	��fV�4� -�uVaN����yF@�.07����t�&�h� ���T�Z+N�W��(�9i	��H����Ă�ţ����z���.�5d���5w�Pn��e��7~gA�EE�۝?PÀǤ�kĭS�b�?��P!M�:(�|�R�R%Q̈;���]C�Z��Jq/���Ő�V1�����,
�C����3�����eG{���Nu�6�IIY�Zo<䦕W]�j��L��ǖ�uD@N\ӠP�������σ��)Z1�	��е�K�PB6��Gސ`Re�'W�M�"^*cVk�[�1ؾfM<�%7~��V��%��Nʱ�^�Z{ Z�c��S�͎��|�j՝�����Hi�4CxA��]l�Kt"�5�r&�`D��N�Iu���]+$�hK�e�K���b؏��.���I�������z�J��5�� ��;1�mB
'8�b9Rk�H	R��^Z��O�L��}��A̔+�L�̈́�"�Ũo%WZ{��(�i��p��T���N3l������޳ؐ��!eP~�9*�l��ɗד6����a���X�V�m=gJt����x�����ӹM׿o�,*���C�R'��eZ;:�<�w�����Ռk$�?K�8��KT]�	1#D��"�"	��:N�l��DYk/^j�x���o�����M��{DЮ����(q������)�S K�_��'����D�I=���N3x �6ڲ��>��(UQ�r[�aPwR��V�> ;R�n��K$}��2�nԀI�_*�Y*c�S����qE
�[�s��.H�,n��(0��o�s���2�!�Tʞ9J%Mf��ES�-���wSR��R�ϣ�>@�'�q����Z���4�2A�A ��a�I�kj�=5���_����H����c��QЛ�_�6O��6�$2�YY�J6�~���+�Ĭ�]]yd5�Q�����_�ؾ����������hm��&N���T�I#`k�i�������Vx���P2mRy�����~�����悒�c�j-��+7ϚS=���� ���HMMˊE�K�ְo x�P�6��v~�aW��Do'.�>B�@)��Ϥ)O�Rw2�ш��i����i����"M�����Tf�g(Ӏ[QX�5�����y�f�n����/n�B�U�Ton�L���p��!]m����Lp!���{u���/���p�j��!,�!�XҮ���iТ�ߵ�Ň��?Q<ߌV5�=��)���\�|��\/XcF���˔�8^�";�&����؛yy	�P���������]]]�\C�.b�`Q�
�ǻK����O��5F������q�������O������� zۀ$n�X�\����/�c��$�8�.��p�8�U�}n�}��xXXږ�|��<ݣC�B��[P�值t�#
��r���b�֩ϙ�����)�Ɏ�+sr�Wc��B�F��lË��˦	Q�5��L8IQ�~���.�ze�f���ݤQ'�Oh��E'T��\rQBs#����
��
� ��s�����+��{������@a��1�Up}���6�;@"y݉C��� ���zBoO�F�zA[$<p��P��L��~PMC���	�Y�#=>1��vE��3�p�=5}�2��a{模/>5=	�����)1�lC����2D�P��kIs��Hp���Y���v��UM�S���_ �zs�9�P�R7���gC�'��l d�|m� �!J�21m?./4�(<|h|І�8�2�3��KW�c7*K��j���4>J$d�E	7�8�9А�Pͥ�lӴ�`~z�ׯǴ�������g^A��d�SR��c^�5�7
��EXN�]Ik�T��u]��UD��-�4�<����T�!a�V�3��aއ-��{644d3*è�C��AQ	3RVQ	�ndˁ-r�)5�*�f��S������������������jՖ������$�BB��D�,�=��f~����{�p�p'L.�d�{Ǐ��#��ǤCwv�7�I����z�s����o��6�}�
|��"�EW��<o�c��f�nv�Į��ͬ�����.�!&ߪM���w���46�,؅�"��NMy^�D��B�ׂ=������E!T����h��F�D�*5	����JN�'
��OG#�0�'vww�~�y�:>_9j�����mVg'�(ijhuCRr��3M�G	x��bo)�a�*Ab���#�prq�
��`���l+�v<�&0\��s�נ�Ѭ^��`��DK�uuwCU?���G�x��Ȱ8$���2+��v��m��8�#f�4�N�n|�y�ˆy�����-�`�"DF����������qNۭm�m�ֻ훳���ݲ�@*&�,��E�5p�#1�)��ǻK�kvCš��H��ץd��:E��)I-R�g.��
��JF@�~���L)>����P�}���I��z ��d榬c�@���[�H�~���`�dZP��oD�)g�f��eAo�?������"�m�&M�@)���5Ǿ�۳Q
a�����F����ahZ���i�eF�D�J��
����^;%�P-�A�*-M�f���CY��g�oٴ�#��1�=�U)���e�,�y�ב軍��v>v�|@�/�t~�����%��E2b �Bq)�`ib.�F�3)"�!��}c��"��)���Y��h����t@�k|�ץ~P������s��V#�����yw\����cF82J
5���#��~�@>����sF�c~*��9�]q}������.!�4�r�$�	$�f�é�s-��S��|�k�������"J���306�Y�2�&�l�U�Pz��ZVP �g�~�:���[m��{����w�����F����hw�T(�ֺ%��9C2//���Ti�(:/nb||��2��,v�".��|�zCߴ�t4�Z�^ϫ�����z~����"�y��� EE��Y���2��m���e�.!����y8>!a��,���It��JIp��J����\LL,fp˩3N-�a1��dr�8XĢ�T(��Et�n�p�Lg���XU��vneӎ<��T�MN�v�����0�$h��N�Wl�v�ɷl�h<���?�X��.P�ah�@H�UTd\)H������֦��^����>�	�,<Qt������r����~x��1�fg��K[���ܚ�@��"UY=���GD8�A��!�����+�6�b��0rhbOM�d��Dz���N�����9��x�5ѐK�"z�]�yc��N�`0�wmM�D� �*����N,~$^0��@��f,>���l��n�ÿӶ���؆و#�@����dS��p&s4��&��M���dgol���Pt��X[;� !I��0r
�dD�'%&&����5Q��c���+�S�⇚M�(1��q���+���i_��e���*2$/����$%��b?q�_^�B�9�	-!�5^�|�h��$��M�>��Hiy|z�c����Z�k�W�RݭB�7�6���?{_O��x1���<�x]�9eK+E��K�H$��o�$w¡��%��0�%Y(�o��đ�N��g)��Q"�%�;w�Z�yjÉD�s+�=m�����\��5�K����f�/)9Pj^}*��m���P"g\  a�c/�&!4�_����ĭI�PD�妾�� t%GІg��ܠ��>9�5cZD/�a��,6!�����Pժ�������e�r�U1����iR�����V�1SFK��؈����j_ḣ~MM��Yxg�o��22��p�J%�;HA(_]�?5��M�>�k���� ��,]���nCu1����d?��.U�ۭ016ɭ�H��P�R�47�������a����{,7L{�e7�b�r�=d;� "���w0Z���]��n5NHVũ)E8��*2؉^�ӡ�����7��l^��s�qn�|���nU��)?�-..��y<�Q<s�<������*77�&Qc�/��.6�Z�>7�A�5�X�ס��	;�0e0]��{H+]$h�����v���lvgys���+w��T'J�0ߛ���]n2����V�@�����'ƙ���N��܋4#է�7�5���S[qH��ϩ���8?���#Z� ����\*'���n��'�1¾%��l��nN��o� _*�eH�w4��y��QЏ�R��@�Im�W#����{x}z���(.a�j�I"f=|��Z�r���ѝ?��$M��;�>��)�io3��'�s�%�WX���<y%�?��JW~�A҂HC���ܿ�f�.-^N�C��*E�a����<%���up��ۅN�f��~1����n�q�C�(�U�B�C�d�R���x�\��ly��1�.-Y�v�ۚ��� �M��9� e�����VS�HAN�K�Xc����~��Z'���� �z�+���½��C� ߵ\m�����AC8oN��6�)4qC�3���I�Ur�+��o��rC?��O�Cl��8?����S͛��cW��+d*�����5^�1N����$���Uge7���&��H�d~�߅�a��'kW���[�>ĭ�6U��=���2^-?����,������qW��f���~ ��\__��.KZtr���<C�N�����|�n�8�!���θuq�E�'��7^���M�k<��5��_�p�Ve�Ca���J,�K�~���� +P.�,��C�z_RV6��6��8l�a�����idd�/�Ǟ���bu�[e���R������4�K�~&�p;�.no��C�.ɴ�,�>�r�/�+L��f-��L�@�� beq��܄M�N<�2�"��X[t2/ઊ����ѧ�:LS\�~�p�J2� ��(1�/�X�t=
�@B�ݚ;P�'Qc��M�z��g�I�u��)��h����7�-�%�v΄�UИ��/E�H��~�(}�Q�;y�n/)���|�4�Q��j�^�~�b_���(�?�.R��nhH�Z�7"�<#nFA�y N>T�+�H��Fv�_��~�&X>��쫩��+�Ķf�������K�&í


B���X>�7���gq�J�`Z��c�;�.�*���u8:]�f^4�Q��&`���~�D2�����%��g�Q�J�M�i�E�A}�Ý>Ϟ󀂋�����aBM� 3[��D���+�V��	/T_
'\n��u�y9�����8ҙ��|=K�vb�Om���XB���_�����It\���@���Gm���kҋ�!D�A:2�cU�lj�Z�W:��a�g��%��r��G����%��bn��d����:��k��4�ş��9@�3|�5���ߺ���#X��	ɋ�Yܤ|�H�KU��F������u���R�"xAԱ��b,
�.�����.��A
���e�7�{wW�7^ԤYQt�:S^^ޯ2��:���Z��Ы����wi�+}���gX�p�� qbSvff���ӕX���k���K���2�R���Ç�ɥb�<�7��/9{sV��s+������a��̗+���E�h66�1k7��u���Z��e�|��������|ƽ��Ͻ�-N�=�s��U�c)%Y?�{k��F|8`�[|خr�٣|P���2`�%^���i1��s�"M��4lO�S����м	g�R�<r��ܾ����;�EL�ݣM���1";SU�S����oj� 뎽/677ǭѨӑ�8���;����*`��]]��M]D��fvV��0��&;���9�����<�H�)�񞯩�Ϧ6[(y�����0�_I�{{ii)��x�:E�����o��2������!�o3kی��-$�7{JI�K�\�RL�b�?wݕ��}}��Q�VA1�|�<��o�]���P��4#k4u!VE1ۙ�||�t�gHk)�I�:6��g��)}~��R�P^�9�V���l���ǝ{�ũ�d�	W�U(�G���Rn@G�Mۇ����F�l��l����p&���T�Ę���#���=Zjb���2S��E�R��?������ ��UŴ�77�{B��d�'�L�F}�$>5.��L�7�nnZ3���Î���Z(U^T���rgþ�g�-���{w'26jkk}������B:a���t5'?z�W���>�u��ijF�*+u>8󀨇�k�T,����L�6fZD��\i� ۫�}+r!Q$|��ED9����E[���P�(4
�IC�Bd�ϬVBR�xy�㜣؟���df�˒){��D(�O?�
�֍�n�C2�K��p�y�]��w�g�Lu]���Z��*{�z���pa�j�۱���y����zh�^�-�������S�:#��mz}ʯ,�@�UJ�Mmq���T�@�~W���X
{q��(e����%i�o�,@M�>����t���:ݎ�I����a�1g������JJ��Y��41#��B�����=ǾGSW���KoU��7|�u�~�§/C��w��UpDz�6��M.�-6�$Tr���
�%acmDZ��Mtl:|:Z���_�xG?�FI��'��2��R;�s����'꽥�Gb���ԋ��7#Ea U!���n0���)`�b/ 7<� �\�4��C���Ƴm{�mm��6�ٶm�6v37{�i�͓7�o���?��g�k>��=�!ō�t���@c���r�y$$w)���VUo`I<]m�+`"CWr�$f΁������ ���Xߑ?&Ƥ쯪���9xޤYSp�uL#q/�1[B�7juJ����oP��ْ�W�^M:,�t�IZIw�N�z���W###�Bqbۍ������S���D�Ó��fh$�E�����|N�	T�xX4��`i^5�_YVi�b�Y�����:�#Y�F`(5vz��t;-��F��V�Dn��ds̅�g��&U?~��k�7*ƅ�*�&������1��ѥt�=�9q�niҌ<�_��"�N��dt���x6vG3���=!P��,�A�;#���y�l�����f۞�CC���ޝV �*E�\@����n��Ӈce��"V�tT�!`��֜����Q
d����B*����� ���Rm�:M4��^�m��1�(>2�����rT�[Zz>'��=����}�C���!oA����p�T�q�u�-��Q�.�ZB���%ǜ��G��b���C�I\�ADt��%=�p}a�j��.m{X�J�A"S�d�`�Xi�77y�/f� CZ�;��:f�������+�����n��ߏ�D�y4�Dٜw�������z��0:��C�ݐ�.u�7��_�N�J����g�ST�/��,(�״���{�<�`6��HY�' ��ڊ�OHh��M�)Cxa*�w��@�0�+q��0-_�~����o�����>i5۾�}��\1�������"������v����}KB�1�
<!ЀJL�rTY�h���g{Ĕf褤-��H�dZ��m�(��L�Q��&mRR�!1rJ,R�b�*���jF�Z���*�Z�6.�R�{�#��*c���B�]ې1Yîѱ3��t%��$���	�әg���U�W���$����a�bC$����&Ίͳ�q>�r�;����M}W�[�kXpد��`~`� 'ǿ6?�
�6�3C29�� ��CXd3TUЋ�eI���WrC_�n-�Y�����]Ts`$�
�+DǄ�����|W�g2A_��'S� 	���9��m;��4=[,	��r8�״�����B��Մ���;����#	�_��m˸�aj0��C���*-���NS�]�Uص�?�����o��biD�����ئfR�dи�	iIV�����1���BB�:PYY�QT�5�����R�i���0��Va�j�Q߶8�mO�*~n��:l�RdQ��Y���`G��fc�
ǳɹ�Eɏ �ew�M$ğ2W.��@A.T�*�ю���8=��|7���Y{!�F>��k�<����\�$�zCFUm�V2��/#M
�nLM]|Ż_��?V���UI�g���z�fj�
���҄��]MD�wr�wuEB<P647O�Y�u���Ý��h�R���z���]3p������/��3<daT㄃��c+Nnl��)ds�����Щ�~=�)ãS����H$ Qu��z���V�\�RA������^P	����P�5�,���z�B)k��
^�P����Z
��ol�p���v��W�zHqh����bύ����֫��L�dS�2�|�th6ճf#uZ:�ҍ�]�O�U�i',�J�c~�.����[#][)���E^�MDpi���Z�Z��d;A}=����𨹕����D)-I���Cn���=��X.Z�3Iq�D���ā���X�ia��d������ؘ�շ�^�E5�1d��˜��\�ǮMĿڰ�@����H��43�p�N�>wk�
����@���S��%d��p�6�wA�.�&�4�GbB�`�x��߲t�z7�국���Q��u��+	A�=����>��"I�y�kzX<�_s�t�C�/O:e�a����w�i>���.�xb��v�ׯ�I��UI�o���[xY����Ă~cq��X�`�?�A<�������ƨ(��?1�/#�.��4��Ё��23���+Y���E`��%&F��INI��߇�]��gZ�H6�SSU�{��{6܈b�r/ok���<�C����G�e��;1\����߃q�� �4�J�~�h�W:����p]��=M���
c�h#��Y��*@�����P�_�i8��z�[�0�$F@O���5�ј,o�E�]�S�I��	 �d����4:)�K�g�pfBQ/�1G��g�K}_<2�b�yw�}�ȧ�x��zd
s��f��#����l�H�|T����C0 �s}xݥm���[���*�~?V�LU��T,��O����,�}�d$��I�Åb��gsm����^K���߆��5�������o��B�����4�uz��MI�	a��wc��ϻ��i�[��X�EMRq"��ۥ��4�<��쒤D���;jH��\��R��;17��,5�s�!2�X�����tt&���w5�	��Uvy����(�~ �_�ER�Hb�{+��]k�8�����M� �!�pݛ��3>A<֧J���3`�$�������tL����gr/ �,�ZJ%tÎI������fʣ��ή&Y̿��a��q*22R�� R��uN!�U���b-��y?�c(����,����_��B��њbB�����n�h�w7M���9Q��PX�YcT�p����j{��1�� M)'�{m�����+�k��m'Đ:پ��#���JT�R}�)]q��|�W��x�g�Qs�6]���-0S/3�*�~�i'�^f�!��ߴ*�����"����?7�H���W=7;�-՝6Jy:��q�LY�Mtۜ-�����Q�a �����r�<qHK�",[Y5ɏM��z��j(J
!���ec3��!�,�B����[?@��\l�%����t�a
�B�e��򟤯|��yB�[k�}��^����-��/%�E*�9���d]w�k�������20X�x�2͹����.�"Оk��8�Xb�x�i�Ah9]w��߿cc)�j'�h�(���v��"h��L���H�wf`~H�7�x1b�t�( �gz���k�s�C7�444Z�����p]�>[t�"Aڦ��3Y\v���>66U�1^s�X؝ �N&�y�3��@1\�^�=��R�x�2�s� �Ԕ����>�NOϧ�4����ǵ���;�j�����^BL����((L�u���_
x�B��DFE��(�&R�`'7���f�LY����4�����]���EρKC��Ǟ�rdh�[m�nL��3j�B/'���d��Rҍ��u�.=�]>�G�!vx���F���K�QֽL>Z��9\�������.�Z��z���m�{����Lի���f��o��yУ�D�8;�}�E��݂'���
]oh3�@D5�G��.g)JtZ�@��273�2����JII�$Q����,׽�VːW�+ss��ж1�?���F��mxnGP�ڬ�ԍ���tU���r��KK�!b?�ק���@���$�(ۀZ�59#B-/���$�*��O��?�W�&X'ÿ)]-�J�G��W�HQ�т�d�J'6~�]P��J>�����
��G� pz�V��L�i�Y�<:>fP-2�������8l���%M˞N�Idђ3kצP"��%�j�����Qlgf�[\��mV�p���~�$����?�/4 �[��t9�n�y:�j[��z��v*��L�F��'wI�D*��%IS� ez���Q��)$2�.PMW�knyyYd����R��z�	�hU�9o��8	h���H����u�����&b���i��+P�>��EfJeK���GN��л"2���M�4�m�C�DKmR���M/7'~eh�~�7��8o{mmvEX�[	 ��DB�	�F�m>E�]I��9���bd{DAPbm@ݜ1Գ)��e�e���LI��CqCN��b�Ѓ ��O�u3LL���HS��ۻ�7�����[R+kkk���ww�!j��� ΑP�(�I�L�^�B<OU��Y�ꈫ��kbp�?rpr�W��3�s�O-M5��o<.�`�.�IB���w	��	t���v��g��zg���X�G���M��N����:�N�@_�i����C�͇+��k��-V�sP�bH��b۳�ߠt]���96�#�f���2[��t}gw�^��Ϗ�NQ�J�\�J���겲�}� j��l3�䉸����ʿrX����^���0�O�
��u��v�����ο|xL�?���s�c�1A��Y|�:|rH� ���vg�4�R�]ct ���B�ç|�`,�B~���������/#��t=O�c	_�WӰ���ݟ��ۻ�L�?�w֡�3�e�jr�!�*(x*��%��:�Ǖ]���ow����C��P;�}�2���{�؟O�d|�T���v�:c�H�4�3�)6C:*L
p�DD��P�7�&W?Ր�kaw����2������:I"6[Z����h�w��� KeAS���H}������TUE����=�����g\�����?������8���<!��u��9d� �Z���G�t����� (YH�\� �%�Qa�XA�k\k� ����idد~~o�ےX�o3y����V'�<	e�B���y�;�.t�4��SH���m�EIETnQ��W�^ME��Q�"�Y��%�$!�K�3��b/[��͜J虿q~�R�vA����ix�DSC�HE�kAr��N�8���W]P�C"LL}O֫-߅}#����5�;3�~����ў�2a��^�Vl;7�>�����:�C������ӟ�,���/?�d��?��q*�)DtzyٖR']�/8Ҭͽ	����fg�Ɍ�e���L�һ���]sm�^=�����t\N;����/z|���Ҷ�n8�>?|�hafN`cb.9ѳ��y�������\RJ'���
G�0��o�/�03�4�*
M>a%A���� �&!++Ѕ�$5Q������'�FE��ǆ2�n"�i��8
p��� �%=2� }f����M򯪪��AAA�O�?�u��ۘdz~zi Go���P�b�ߖ%��W&'���UU	K��`��`>	m�_{fv�������Tx�3
�_4O��̎���Q�	�#p����u�������y��9��Gݧ�9u�N+��Ϧ8T��/�^���S��׼��Y�ʻZEff⵷�-��Р�A��˦��Wדnf�KMWb������W�������9$�I�_d����3�))pJ���c7�'��e����k��|�l�����:�(�1A.�Vo("��,�|WGNm��!�Dp�D�[�cr�5��-�G���)�+n���AױP+�c�陘��/ژ��� ��w�N�x��{�%m(J�/��ۚ��l�ف�[�?��=~���K�V�x�i�������STS$i6O�-^t���*?.���lq~z����=��S��y�^2���V�p��DֲV��y(�+�:�Jú��|\d��
$�r�'�E�h�|�.p<_��%�V��J���g���Y�R)��Z�t���8�*���$�D}7���]��ҰW��(K���K;�.��e1�[�
����ָ9��ސ�.[m�F/��:��Eze��m�~M� m�_A`` �A�%�t#|��Gy�
��"������%���P����k�e�U%��
��O��tBJ^�܃�&.������M?P>��2�E  	ԟ$|�i�*$�#�k���0������KO�ZZY�uF���@�9�)8c�>�U������Ix�~���!�6¬1T���Ê��N
q RJ$�$���j����U�XQ�Vj��u�������:픙YY���8�!�6)�H������g��(�ԔS�Eʀ� Z������XC`��yˁ��H+�6����M�#[U�<U^��>}D�����2��CD4�T�&�٩�B���#:������W��60``,၃a��S�����XO
l�!���G��M�������{���enRu�L����{D����Ū�T����SUI��q���F���GE��`1�E65[������v�a\���E��WiA��y�LE){p3������]k���82'�I*H�M#�8{p��M�5c-�' (`UJT�!E���͘�����2�l +[��ݮ����7JX��$"5�bx��0oGGݧ�tb�������wE\�r��Q���ޅW�Lxk�ş֭g&�Mv��F�$�$x�s���6vz��/
�ۏN�g��2\_��8Ȉ���2;g����'y�0����t�VxvJ����y|X���Y�t�����s�x�Er���i�EN�E���8��2���Ŵ*C�p=i6z�?8_�����m�~!����y����������[8�TKWYI	p�]�E�����E��,
A`S\�Y�q�a뜛y�f{M��Y��U���ؖ����Z���4�������+*>6�ӓy�W��$�V/�hV1Tk����5�M�iX9-���>T���9$,	�0�l���R��=}�"H���L�i@H�d�F~X�����%Ѵ7	VQ�0���m�s��[\20��)�;��p��1�VMEE��D"�W��\w�@deeY��[��RWW'�,�fB�Ie�� @��ԯ����'|�a�]SM��yQ¢�;�q�F�!1�.c�o5�.����\��;$��2�W�Óƶx�Ȩ6��JmǁA��/)����	LS?#����wl`�f��q�P����tml:�ٱҖ�ޭS���kvH*��n��������"�����[�h��Ջ�}╦���r��׼���$�O��,���C�n�m��wںoLHp����)��*}S�����yJW����B��!�YD�<l�x��L�ʠ���7aH[���_�����us4� �L��:� ����c���C
e�PTlu䓦�W�4ǘ�{�Y놹�c�o6����T��w�Z��6�$w.O+;�?
���l8ogk�Ts��Cp\S$�rm�[�?.��u
p�+kqMn�wv�i5�O�;99U���'`�M*ԕ����l\n��7v�>�R�ou���"���mE��Pc�n:��`�H��U��p��I�4,EP,,R�R�8�\���1���Q=�ԫL�_E��Z7CAC�D�%�.˕j�f������:N��I
p�:gEh�h���EW_	�(�c�~ �(EXX�ջ�=m!��\��!�,cFXԫ�ƠP$1�,�0}�#Ǆ���@u�Y�ቤ�UEW�w��g^������w�@xHl�Y^�1���s��������V�ɏ�V���њ7�9ӥXDP��t�&=�e���� �kew�J�;J281�b$l���񑏏��Qs�+�:IX{b����\���hL�$�i��,��x�Ӡi^�%Slc*ح��'/�/�D}�=<*g��8�7�� �	��������{�
��S>��fĳ�C�C���#�+�+�k��!�]oE�g���ã%1�}{0U�������(vI�D��,#]c�xb��e,Ǿd0R�"$�a[(��i�߆	�������<j�?�hMF�r�(�o�t�D9���Y��μ�c'5C�.Q�����|�v@���������E-l'�����P��G<m���pB{ L�{���ׯA��u�/���'A��T�ތ��t�QNp�M
ûQ��R�������go�Hu$�LBI<2�Xw�*C?���Ƴyv��ŗ�I��dx��t:dA�K`�uF
�����ު�����␅�Ir ��Xl�~��l\r!�k��x��{~�W2�3��OjF��n4�N���ʪ��p���|��Z�jC'1
��em�?�#��D�=y���}B/H8!{�>�#�@�ٌF7�����)t��4���y��ѳ:GG}^ʄ̸��v����`�Q�桓�
F�:����L�����b��	��}s~�QGᖅB��4�z"���a�:����'�7(q5�Ҕ,tg�~�ּt:��Y:���=V-�s^�T1Z��
i�ѧ�qT�Z���Z������y�j!#��,������J7/�gSg�;���VS]]=c������Im�C*���n������FwKCCC*�l4X�swx�������=�^WX�4\~^>��/�;ahWU�2z
>>>��r�B��wH��GW�������@�/HJH���W������a����)scEB���J<�Հ�r)فa��䨼O����k9��� p?�S_
="܍D{X1%-M�l�����I�^�餅�~$!a�ՙ�x��T/9f��.rȕ{��P�&#%�=oA���vŠ|L��� �j�����ABI����w��K�~U�}���Y�e������S4��B��{:�������'���X�'3nE��Em>8<��s���P�aY���0����'\O.<��D ��`\ �d��(����w���`��z�Î����u=%I�M亾��������E�]�~���"GT� ���J]���bڦ�<��)�מ뭠�j>�M����g$�VER����m��-�Ia]��J���Ǔ�²2����<(lom��m��8O�����d�k�^i���+��葿�v\lrv	�"r���C,�G��$���i����.kڠ�DG��A��e��t~��p���bo�'��eP"�o�/5~�#T��5d@�z)$!e�n�n\#���7����%�;�1P(���	�ɷ��e��p_hs9���d1$)��Ç���<�h��,)�l��Dj����ޮ��˚�j���7#zY���~�CT�������t�ҺK�������o�LB|�C;�`���QDOR��1sq#�6'?|��
;���M�d��EPk�o��7Y/
�\�e����i��+~�d-p���)�X�jmm���DF�;�	������=$��ׇ%�B������\�8Pq�%Q��;{f_f�D_�SH���-5� ����}��̽����<[�[�n��Ҁ�S�@3�׽Z�M��[V���4%�;��������v���4��t^�喲����W�	d�&��Ţ`R�![�>?��M{�&H����A��nJ{9Q��	�U#}��Pd�L?�鮿RO=�����cK4/�+���{^	&�J<[A]=���T���@a~�u����:11�A�R��3k=j濨 	��n�1��Nצfg��|���͙o�`IL)=4i@wuU!�p�[���G�'�) DW�&I|�r�Q��:}�\ٜ>9`���V�@�`#::ښ��p�"��q�2N{�Wǎ����N�6�}�gy@��cXd���&1l�@�%|.�d1���3�4�������B�Aڄ�7(A�Y)��7�#�f�g�R�b
�$�v�4
�Hv��@O|/--m�bX����<CZj]C�z�8l�$)�J7#�F�~o��/�],M�s�����S��;��n>n�


�P��)��6����ۆ��r(uY*M���m�{@i����:��r�[����:{xbL}R�!�C~�E��=@
9�`	)�'4p=�DC5���~Y���J���HΨj�Q��d�D:�'^L���j��_�A�N�����_Ð"�$�
]a�)z�B���v�~�miǽ��2��-w
�"r��WC�L7pt 0�l�;�F����oV�5)f��o�ҤCar܄P+f��"M�n���.��>-�u�7%�K��?Ϻ�'PD�t�8��#���f%�@$y$�@;&�K�/��k��P������^�^����x-�_W�orr�-55gOng�U�fZ�+F1������KC�P��WOUwC�yF��qi+=����3y4�k��/���B��`{�Æs��2�$0X�Һ�D�dG�^��Ç�y����9�G�<��ӹy���%�	�`R3�G�K�ijj�X����7���*]J<SB�����;��j�F�>���;������?������`ƴBC�����H��V�� �ӀFN�t3]�`K�v��Y�S����J�ЪP�b�?��K��x��$��Ɔ�+���[�,��Br�.�Q*�b�)u��_\j�o��W���(��<����?I�W���drv�Ǐ�o�<�u�577��!��k�ѹ5%�g�}��I�/u4��\�c�$��5�����w8���7��蒐r�c&���C�������ba4�I�6�>!��8666�O���fo�Pq�Z����-s��o��_���4�����T�b��}:З�v����{�@��@�ZO�������p����>���>L_n�iz��������&��>�7�4��e�y��Ql�_E&1%�Ѽ��!�C�Q|�۹�*�Ò�F����!´�p:�z0 o�+i	�40�{�^BR�������=��jO���R��v��\ٟ���f���B�ԙZ���z���/T­��f���&��E:YH�.|���߰c�Y�=c����,:aB#�}� ��T���7�>��i�]PUs��|���:�ct�z��^�����+'�.�k<��Ke�6#�� n����м��&��r#�Ï�js���q���uU%%&.~~~ �)�3ٖ8I$,���Y�MiS4�Gh��Z=�ap��U>G����<A,�Zd�p�\{�F��z�r(�S�M0X���	RmK�6͠�_8H���Z��?�K���$ԧ˒qD)�8�[ELX�71��Cu�i�_����;z�:�s��:Ͱ��l3NU����vpz!.o��ߘf���,-O����J���. 	��MLL�&=��*)�]?��A��1�{��vƨ�R	��m��)���s"n��co���zP�H�,34{!m�\,�GD݈pnn�|��9��y!cVd���
��(�����#��[�R>�����
i�2����zJg.^�b+Ͳ�Fj��pQ�΍k[!
��$������`naa%$$DMZ:"Dn���ILK+K�	�l`M;�ھ�Qu���S���DDM�i�/>~K���#� 3*"{��z����%��\^n����XdDD��,!���!b�Uv��/�f�J�fllL�=�t��7{C�*�إAē�ߵH����o
矒,U��� F�F��|�_C�r��&�_SS�]]�H�Y2%܎��6�C�����`�	CHr�}E�p���Es���.�����{v�ZvA��ѼC���\<!^�l��&4$V��W[���zWd�K�gp��W��%� O�9l�ù�$�����T"����u��iǜ_�T��_��N-�+m��ꊩ
��Z|��|:�{E]���8+wC�\��3�S>�'���1t�o��~�gX��SM��k�����fO߿	�6�jV��VE��3Ư�L��n��z��d��yL����o���MMM�\}�ٖ3[
8��3���G"���ܻ�t/3�/�J7U2d�/^ǭ��Z�i���/�y}�M��]��n�2�'~��e��?]k�b���g�?��*$ҨD��}����ƾ"�Zy��e�KE"��񕝃c$b�����=�>\5e�]X=��?��"�«��m��ݚ������ !�ᤷ����/c9�+��ƾy����@�Jf���}�ER�~�(摾�k�UA�B��^��
�v.$�oi���D��=�����R5kwL㋉�t]����Kwi7�i^s���|Z�aƯ���䤁-#��}��=}[��
�..��ύj{W�n���2���`gc���HR�8 ��T-��;�O��E�5M�*.a�?�հxf���\6u�ב�v��u��� sz��+���O��#�ܼ���h\I�DI~� :.�=h7�}� 4�̿�̿,_M��L�hZV#���������:���Ļ���]��)�qq\S���ӱ-��U�i�1�K���U8d=�T�o�y�GGⵢ�3 k�2��S��*Wx��L��E��(� 2��z�aľ�7��2Ӂ�Rư"�39ݺ�)���J:੧��Ph�y�4���'��m��K��؆|��/j�;����Jd11%��T���I}���QYY��3����ˢ8�epc�Ur�^Ф��� �3�x��30c� !�2�y K������6N��)ͣ�'�yG�+�����z����%-���&6(�{�A_^nK�� �!˵��A`��a���~�_�w�f�1�#�O�ֵS�� �d�N �HKu@����M�P��1RSעd�ݵo�����q�6�4r��8{�A���H%q��W��]����+���������:��"<����nW�ԼYc�평Y�	�O4��������M�}�����=�'����5,P�!�h��jħa\A�qdwh
��ͪ��F�z���<�k\KiF�8N�d�),�`���m�E�c�YM�. ̲%}�.�ТQ 1;������\#+C�� S�:��*�?�t6
	>���)��u��8k��,��ڗZUuEM!"#��5H���	�N�/t#���ӽ�Á�j�7��$I���z���h=�(s<�u�����w�O����4�Ո�e��<Yr��54���?��Wc��ߩg�Vk���~����3��&��&�N�<%F����?$�9���`ki�|y������S�N�b�A��U뮵:2(��Q�  8f�{;�_��	Z�CCA�R�_�@�p
������7r�AMό|�?���FFb��|���}b��󻛺l��w�:\�V`a��Aɯk�����������vu�b�;�z��I*�#����ã�i���Ye�]u������d3��1��n����M�}�n�i�^9�z�/��iV��������pf�� k���1��B���F�:\�������2!�EO�C���=���n.!�]��d���Tm��Bj\��	�'��k!A���O��]߿�x�f�{B=ˎ�9�6�LH�G� ��Ƴ-���_Z��ls�ܔL���~��p	
�s3���Mn��m%l����5��>��99e�L"���;��%�`K�UKE�4e��XŲ<���*��	�j���V��~�]�iAe+ge��.yР$oA@�ޤ�DT��t���S��I	M��|��ҭo��"�0�i%����1�x���#����{�q����
o"�5�"6�MF�_0���)�����a�;�B�Z�u71�"
u�c1!4��6���t�3�۾����ϔkm��*J�n��������b���R�*�rvrR���g>&���uH��
��"$�Iǲ�ɮ6|�H�SSK��Cw�[D9��p��.�lZ����|}}�Ƴ��6���.�W5�cdTӴ���PR�ZWQ�N��K]6d�Z)���+����*���������!����0C�j�R��_���Z�F2M>'�;��� f�h�;!���ax�A�����D��h�4���{p�h�����놞�?ُ ����w7�/(�Z8'�yP'�ʌ
"��*$���C1o����c@���A�c��l"7%���?�n'�	uv7�͇����e��ӗ����d��R��0R<G�ُ�X�����?���_�>)�9���x��=X�><{ ��&;�a'���&(Q���NHC%��)tp5H]`�$�t��Iz����1�c�=w���,UA:��y�%�yP%1�gyk�Ü�B�!N�Y8��S�w��,�B����t=gtL\\Lݵ������K;HA^=�6��/�xJ��p �U.2���v��;�����z�MT��Q?����b�o�c�cw�&]��K���!�,��;2t�W9�$J�f5�4�㜘n��^/Q}�&M����f�>���*��[��I� Va�'��I´��YT��ÐwJ�������ǸXGG�4t
M*�]�3N�����͵����Մ�n��ȗ��G��v1�_Q�:Z�w�_V�[,�fKa֫����FFyd�_�g+Q����:�4.%������ʹ{��ges�@�%H)�3}Qf��	nñ5n�]{ ҩ�I=����#}���~�72\��tyJ#�M(��zМ$��H��^+��W5���'Ϭ��~����&�;�/{���^����gPP���Q��ǰ���&���@j���r�����tD b6�]��-��Fc.mه�J6�+Z��?�"M"��x���L\dd�E?��I ���\��z�~L�8���̡�~�ѭ-���{>'��mg�,��R�dZ���~����Wh��G�h���d	�M�2�)n��E�B��W6J&��s��[Z���d��]��|�O����vu��)�B87e�t:���5t���9�A=n.*Bi������D��`�Js�%�ax�|r^���0��;�:�5�n��q��j����4�b|ȿ�3g��9�����vru�X( �T�P�;ӗ�����˄_�|�M����BG_�MJ���l�ʔz{w'$�f����F������3�4����=��X��f��s;��&������2�=��_�S��;�Ŵ8KzC$K��7��G�	�P�|ʫ3��^X���2����y\�>���<J!""���;1e��K��V���H� ��������O;@��'e����=��;������_���h�O����|����it�@_~d�ҁt	��4|mF�#a�ou2T�l��a�����i��N�`z|{�TI�:7)��G{a�����!BB���2[40�Pz?��͒���_-���F��$���Z��{&����]�u���y��F�UUU�ލ5��Fw鐪'<xP�f�[T��[����aQ��h���[zL8�]h�}�^1�Y`#Pi�xÏ?�S�!ױ=Ҙ�j跟�LS�v��B,�0E
yFG=�ou�Q��X�(`B/�T��y�Yn��pt�N��7)����p��y*�΋����������'��0a0x8������;?��t��ÆA#��Ϧ:4D������;�5��w* # ܳ��+p��f���3�g4����/��<<У@�_8��w��L�;�d�Z���{{ ��Xȷ8��1��+�`��<�=�q��
l���\�6|^�s�֭���n\/�T�*�L
�5��1���%�f�|O�@EqM���� �-��!���4z;<V�û7�m�O�V���$*�oϻs�/��"#ݦ�%�
�|W�g���@��#��P���5���o���}en�.�4W]]���+����b�6�*qv��A*��Gj��AOp�/����߭�_2�j�٘�"5�v��V�bH�'���/�YGE{�%����N��^�]Q��Ւ�����E�!���s\�����(Y�6�I)�k�X\g��(0�k�M���뫝{�s�ƫJ7�=�x�M-�iJ)��r}g�D��������r��[rT�� ����C��A�'�7���6��.�h4�
Fۏ�{���fd��A���c�TeK]�РV<6��(�j6�(�����.��D�<;E.dK �}<��Y��V����Z�˔im�)�%v60<+@ǞA��@{��St�f!/mSBMÈ���!68�/n�s��!�%��'7�3���"��Z��3rj�&s��jx63�h��ǭ}9m���I������̣�d��F�Fj�k����J�����t��n����^5ބ�& ��W3�)��-�t/b���M��p��
i��g�Cqݓ�+b�n6����c`��k"���Qk�L,ƴ�P��?��]1�|;33*O�8���$��@rbJ���}Xs�.�ؼn޼k��废	�9�v�9IC�/�Ējjj@�wNґ����Z�3�����4^L���tȂ=�sSSߝ&�6<�����.�(9�0}Ii��،ǜVɤ�� V�d���,�f��f)/�n��J������s�Y�7 |72P��o�/��d^Rbq�����B�����ͽ��u{i�,��,<���x\��eA���,2;!U�EMU:β��@KW��¡z{`>������W��*ܹ!�>���_�}hz����C�?��vlVd���7w�g�ٕ!CM*�N���b�3�	NQ�S�u]W��cf�>�
Y���w|�8�fT.Nk�f�_����g����>�	�q��>`?���ܬ��~�pB�k����w*9����3�}��l���24�ѥnݟ��_��5���f�SW���|Bs�.�����]}�x{wl�n3�_i�9v���P6��W�f �9�	\���r�&}��`�h�Lt�%>��������XZZz^�p��+�1�1�`��=o�k�w&�G�#z�� k_�lB�Mۯ�c֤����DU0
�) �{kW$?�1]M�2�a]YKxl<�%{ةmp�aL
���� �`��8$�o���
�	��N�1e�*��M�F<d.=Ǭ��!:��N�YR����[o�lsUl��N����aǊ�F�d����)܆�����C6���!~��"���M���:y!�G\�o����c��;_�F�?E���Yׄ�'�۶m�NǶ����;zc۶m�͝�_{��y>�9j�s?U�j�����K"bG�[}�i=���XL���r����lpuu�Xp��[k���%4Dt��Xd�}Z�;����u݊��j+̂��w�MB�I�ϸht��C'v%�*���h���}l�"	�>�	����L��� �����*�KDI_�g�S�����e�*^	��	/@�.q/������4�!;�s��눘�����7���� ��&�~GK▎�z�r�w&��+F\Z��ߌ���d������c�7}����A��2̦#}��&�Br�w|_��;4�8$�xH:NJm�2r�n��Zx5,��l��	�i6��]ٞz�N�IA���P���?#�{=VOVv�x���>���qWX07WJ.�>����>i�;8�Y�(��G��f@�z�!��� ��a�zp���̍n簋j#�S��婮�߶d�ё����^�IzN��aw8{#$��N�N���a�5���5e�o�`o�iv854�L�z�>�Q(�M���x�������j(,��n�.�
p\g���¶�ɸ�V=R6�2gϗ�JͩuZ��x:�R�� �lkl�tq�G��МG�BĖq�[�&�t�u���':d֔�_�ѭ�>H�����M=z�[����
��+_�6Ε�ǖ���vrɹ�:BO?�
K����CR~#�kn�
2{�ܚ���tnKv/~�c�I0:�����ji%,��B�������u����\�7kI�[�����A��ߏ��v�ƃ�a��:���--Xs`$1�8���<����'vKQs���WŇ�36��Rc��a�P�v��Vh�;�j�q��n����A/�'#���mi��#�'յ�GAV�b�`Gp��g,�6�%kt���}�����$�rk1�BM=UJ����]�s�e=�����'�P�N�|K�M���
x��`�%̀�M$��8�A�Ɏi{�,"�{8�$�;0~Q7&ޙ\v�6'cގ:7޺֚�6~�Ԕ����\yb�#w+F�|���K϶�ϻ��O�^@I�`'�E@Ѥ�1��֖�y�� AZh&q	Y;l��a��hU"E��&E���oш�)6�fI�ۘ3�����|$ɲ�~:�,����X��YY	i�����p�i��A�YiEL�p.!4h;/��n�l�B78�q����z$b�������6�l�8��4�A�񿞰-f2=���w�T �Õ:��Wk������T��8�����S�F=}=��5|���7 i}��ܖRU�}�#�"�M6�5�,��^;H���8Ĉ�N��OXI4Ur�Ҁ�b춿`o�...�n��P!��������MS[��x��괺���Z�"�����SM!D;�!!+�%���ݵC}��6.��׮4�ʩ�l�Z$������WҼy*��7J*G�jz ���j+�/�U�F�$'���c��<,<�Q�$Ƥ��C�P,tȴ􉨰����7<�pQ������  ���Ԍ=V-k&S��T�С����C5.�������μ3��E]�"֫��p�1jǯ��4�" �mǕi��X�(��ۖ���;�()����@�|���4IY=/�Դ5�L�<`��S"�)��sDPZS.�@O϶Z�}��uU��/iQ�5�����q�ū�/��wڃ)���~bU���Y�o��x��� �4a����	���0C��������������"�Q����&0$b�;�c�����b2��l��ȁφy���D��C��r����tp!'�|n�Ǆ:M���׉=���Nf��#��ޥ���v���o�d
|�c&�����|���knn�sAԔ:5��8N�⣐/�_T8��P�Q���(�C��b˧��lw�4[l��q��z�l������E|���3��e�0'!:ܓ���<��}���z�h�[ۧ�t����L�\D��8]���L���`��-��m���FCvP���r"Jn(v�������[�'�A����-'�E�_�|��s�q�������lZ~�f�KKHH(=�`�|�:9�-~Y���o��X�(y������W�Ƚ�"v�ܞ87�Eg!�f���
#�2��*I��q"���W��{g���7��������E�/���*�z��$'�	��������Cs���g����i�4Ҕt�X���i�g�8�n�n�%V.;W��\�����Xt���O�P��}��ӿ	�8�ح��g:����[��{������0f�h��Y[�=E X`�p��/H	�5��v��཈��|R��޳�u.�K$F�L�E��S ����ћ���&�����ʈM0��Z�џ:���ҭ��g��~
"��=_�>�s���b�v)�P#b�"�#{dgP��G�h��hD�c��3���
nH�����"φ�#t����<�ӑ:���T	5d�id�f��L�5
/�����W��L���+�գ�<� ��M&|�@Z؝Z��'	7Ӿ�[��	�bb��i���&�]͘~�
ܓ03}O�@[[�3ڵ��1�����5c��������������]�g��U��W6ӻ��V�.�Ӟz�BM��>�VFJ���|��]�-F��i�!�+��R��y=��4φ0���Qa��K�T`�a4����Z���,�efK��:������*U��H�s��'|�:Q	���\�
�:�\��?y������܏�L�e�Î#��f��bl�����t�Os|}��}:�i���M�����B���(��l��w��D3t����q1�q�A�MXBq��;+: ��W��gZ64���i��R�锣D�A8�kee%#%5����%�����z~��f�Y���!���
�^Pg��^o^Q�߃�3��[B@[Mj�/]��g��M�]x�1�xPK����.tw��>GFƌ�3a�o�+Ȋ��v�����FQ�2�7;EG����?����Y/���,��Lm"�-m�g]Z��KQ3��J9��і���{��n$g���^S��������5p���LG�l�64WT���n�zl�n�Ob"~W}�R��(j��[^ecc뇀�(��:����9����i*4OA�����|�H�ɒc����Ǝ�S�䆏��'S��W�TK�d^S���4s���9���'ʹ\ش�ۯ��0���4\*E�����ٶ'�@��խ's���e�.����8xcn�v�J���H��{�����􅱱��X�"�x�J���~r��>@h�y���tu�5I��ÈB���\�Z�U[n<n�����������6;-���0O\���������l0珲�;fTQp���?11ySc�s�Gp�h�z�'������R� 2�.[��~��x�r\}Y\��ձ�&q<U *��(U�a!�ބ������)e�D�:��k�C\Y�m�p_�1���Ɵ�������lC	�b��H#B��@T������u�b�u�p����"�.t�/J\��v�{��<�Fh�Zw���pn�uV�)�b�!N��u7��q�h^�Z��v&��<����е��$>U�w���M�W����)cg4q�����n�mo(%^Y�������H�O�F���B%�UR��F��*֗���RC@T����i���{a$��e����۰��;H�V�_n�����F�z�Ӯ�����n�,~N:��X|U=���Ee��y�֐�L͞�<b8���$%�DɁ�h�(�;A�Wz�_��K"_<+��j��������}	��{q�mJ�\{���58�-�z��
|@�dJ.�H�a,k��R8	���t�5y��t�:���騔��D�x*Pxh�l+�91��y�T7�ѱ�y-��?z�f�r%<C����lR�p0����ۿT_��<�zo�"�@C��O��9@��U��u���ܭ.߷���\e�n&��+>�!������>���I`>դ���傏'~xx Q�l����?�Qe1�����e˝��9�p��J�#��B�ZL���^�
�zy�3US�n�BM4��fs2���@$Sb5�k���}b������5II�����:�������s�*);-7�)=/M�l��.��J���Huý�N��Q7��t���W�!�)w7�+�i�"��n�7����{^���Ε�ci���B���]�U�I���}��n�d
�ϳ-Aa���vI[��;o��*O�������[��$�1Lp�����mY��ίߌ����Z7F�\�V���{�qW�OPF郌�@���PBW9dee�����p�!�t �e�� ѹ?�	������& r:l��7-��'Ml�����q���w�E��(�`��N�O���/*7Ư�~����
(g��- ���*u�`�k�_��s��:�vv��C���6��0��?�k�_*=���I���c��� ���K��H��U���s��Y�vב��{�aܰ��K|ܨ��A&������9m��I�y�>#�N_���^ȅ������:�=����~|$ى�JbH��AGZ�3���vH��JbG�>6�b�>�q�K�L�̢����Į�td�g��s��t�1w���$��P�@RT5?�{��Ώ�S���2b�h{\)�s�n�����h������XU��ţ��`xT]�p3D줢��aXf�O�*+��y�_֐ϬK��ɵ��e���Sz��{�6qy�l���tˤQոs���.F�qy~�z}�fqq2�ԫug��n���ѱ�����h;Fw�F��h����l2�}��F�N����䶗��LL��Ʈ�=.�}�@{`O�ȡ�y����[���s�ωLq�e���u��H}��SւR�
��Z�b�CA�,Ǟ�+TJG���K"��ET��mrM�C�]�վ݇�0oW�����qa#����R��qR";�r��0������h0l&�s�iӱ��j�ϴ�<v̩ό|�Eb��h������244tr3Lh��?�^���y�?y�|�Š �{�-�pu�ݬ��}�#�{l�������)kR��
������ ��*��Ԭ �"�H��gea���t�6VcƠXh����Y�@��er��{�54Lybi��~���pu�=��,��#��BҭE�����"�Ɛ�H����u�Xۺj�u?n�{k��&�$�D�6#�T/������6�H9�� �����:�G�t@'�C�8Zp���x�@���]�Ã�t�e�Д��=���>��=��
������e�K����D�x���3#��;�/7�,�G���ϳ]!-@�/Ck�`P���2cL;<��^��0
m���Uk}g�/W��5S�����GlP�{�)����a{\,�+K�R!4�<ju��"�)�v�Oj9 �\��*8��z]c��n�r�[5C�X�d����<�����(�Ŷ�G��+5�#�B���u�����KV�����#`�ӹ��^^^'���ig�O[$�Ft6�*��@+ ���#��6�bC�I�w�����֦����9%�~8Z�����~��/�"B�b�u`u��>����E��Zz~O�|ԝ5���J)��/�:�_�����;����D}��|��8$�
��MCq�ލ��d�;���oA#���'���Zb�Jep|�G�\���5�|�?!J��i9]`y�N�������х����/�}��1^%�K+&����S& w�D/�����-�8G�����qˡ1{N*b���P�T+��)梞��N)F�[ꈋ��
|,�T�#��[�&��at�k�Ɣ�9�=\�wd��Y�����qN��E���r��^ҫu��Z\j#q����æ���P�:�9&k���筅���<2�v8.�g�vܴ��K���c��E�h���x��=>��n�p�˔�f������~���2`��˵��ֽK��0����)|Z^a�H��Z5`:�{�s�2�ԡ��x��M`�^�y~U�����?�����v��c�GN��z�H6:(d���8{#L��mu�5����K22�St��i���B�>++i�|�>��n�}{�����q?E(�J���ʺ0���6]
�/�n��_ͣUh�+����`�d�ۢqԔU`�~U�>C�@G���A�����xnB��r�k��Uܷ<����.+3C�����t��h�Q.Q��,���|k�.]S�?T�=h�X���2�3�K;�1�%^/�Z���!���m��:!LRp�9���g�M�q�Ġ�l81������ �Ub�%��?�Id�{�p��(���Pb3':��� �[��0�&_�F�u!T��T��R�n��a���,�|�J"PmYT���~��c3�kn@}�z�vmp���+��X��� �=�g_!O�ʆ 0��wz�vd.�[�
M�tk������j���ne���J����?1�oߞ�iE�989WluAi`�ԑ����UĄ��1�aI�B��K/uU��NN��/&.�ptur���
�@����'��&�5b�9�<#�S�o?�!s���t=(5 *y�w����l�Z:�D� =���;�o$O�]i���]�2y|]��ˊ���U����<3L\�~���C���E3(Rr%ȗ 654L������)�T��n!kbi�y�hT}2��0��q��r�����1���2�iV*��j��@�DC�]�^��ʂy���L�m���_�������Ŧ��-��C���8=�u�1�q��� #h�3��*�腍Jx_�b@��{�����9�Wg�-�ewƎ�@�ӫS$v�>�G���p'���>�� +Q����C�”Q.I)�^���Dگ�M��Q&��=�8�v_�ea�j�-T۴���.��
,.�on�0���{��[����^/�ش�nqMZS�-����?�h�w�+?�y[�O�������ش��\P�m�-�`�_jЦ��v�a/.+���3�ǖ��=�v��g���)�
��� �=%����&�-/!���}�htC�o���k��-�S�u���ο��ԩU��~@�p����O��8����Q^ec0���O}F�gJ��]7��^���
M49q �[�Ԋ��#ؿ�/	��~�ߏVq���С� �fՒx%��T!x_{+47�&_���_ðh��X13|O�z?��R�?�M|�u~A�Ik�*3��#~z��[�gT�,��Vy9ڋ����荰ba�ڿ���)�ވ�4�����h�pDU�}c��SԄ1��������n������믤�� �I�^��0Y�5�F!c8#e�X��o�D�)��1�]��8}禷��4X�*��f�e�뽪��5|ݾ�7���U�4"�M'QP���EW�������������^q ��63��v.���^��j~WfV���FƟ^ا�Wm�=�9��|!��M�RX��xj��.@4ɱ���A�:ý0�g��s��^5U7� h(�D�~�13���.�Ø+���7W��V�s%�F��@ˋz�Q��w z��Y�������qB���QG(
r��59ko��C�ˑ��L*� ��ɣ�(V�%E.
���9�Ba&Q9��������$1:?�ʍYK��\>�	w^u��v�����#��-Fd�)B��ZK��3���޵=�������Tu�������x�B�{�?U��=��D&	]o6jj��H��,b.V[�?�`��"JrO]2'��N��6.�粑d�,����%�:�y�ӣ�*~~i��I�̠6����|��=��L��?�JR�.~%~,V�w}����h.�G�Q���'��O�3�ޯ���9"U��u�Z�''�>Ϙh3��E����@��Y��� �z9��6,+��������������cc,=x���ͅ4�oc�H�V�X/�5�Z�/
�9��sD�q���Z�k�ì�|\s�����򲶦���`��)�O����b���`�����ؠ��wx���/w�O��4a�=�sk��|�J��7�ң���1|l���HRW�3fv�xkd�Ɂ�Q)���Ef7C(��̊Q[�M�
��0��o祒6�w��}P��8�����j}u��Q��~/~E�p
.���e��ܶT��x�eA���-o��?71�ƛ�O�O�K�X<oG�2��j�Mzt%'������R*Cj�jR�Y�WYPҺ�PHID���
_0�8?88�ğ��eTK荣6�~����t���jT���dZ���d���9=ζ�LxyU��<9/����{{5Eu6���T�O�鮻J�"�z�>��x�~�=�	m/�o_[�x� �	���	N���$h�p����.����oB䝌�(�C��_�G���E3>��*n���!��_�w�B��)�F�KZ[='��i>���EA[�H�W�Aմ���G|�����B��i�� �쎍��<20Bi4'%[[[���$����l,u�>Y���6{ֵ:]ʈE��y��}��ەmܽ\n��%�d�)	p��`q�� ]��N�d�[ZA�\PL�)�����hu~�cL;�ӗc�5��C�W�[`�J�X��A[^�4�G{7Gmzj�Z��U8��@�7�>�U@-��9�J��,���f���Z�/v�׾h8�~j�PZO�/�~��6����I�n|�����F��,6���k��G�]�ݤǵ.�I� O��E��R�N�Qz���q�=�+����q�WGG�=���ʬ��O�:�� 
�ʗ_��x��m&��8���������`B���Sv���p���`������y��h��b�
�������/����n�yc����]Wu
u��2GVx}��]��a�{UX0����kč�h\����I���{��.qD�7�xi{{�e瓾������@$j�8������,N��6 �f=H��9�$P�f�֛�N�2pc{��{���?LTCC#���BI�ϗc�oO �o9@���V�B]b�������\��M`�B��h�G��3 ��Y]z(���bM���-$�.�K���=&��7���7]�i�7������Z5��m����荫��6^7�BZ6��{	0z��f���e������0�=�\otg1h��,�E3]5�@�Asj�=���F��Q�+�������!L�k��M���Ƈ�eT#�7������
���+�!�r)�������iϊS����{]��g�����"ݚʇ.��ޫ��X��s�l���ʭ<�æs"��rd;�b*���j���Z4JJ�)LcG$�~�L�e�M5mU]UU]]~��K#�����ʊ>�y�5���W�B~��j�6"�.�l���gw��X=��C���@��?t�}�L��!�n�&� -�`��[J����b���g!�b��z6B��`,�Uan���͠�2���O��pyi�"k�9��ɏ�{b�E���h9?����#.!pl�U̈ �a�(�Àh�c�H�u�O�%�[��L�F
��}�Po�B4 :x�	�*��]d�;>�Ԛ4|{���qJP_�l�q��{L�
���:PuF>FAF$FTH����
PT��>�K԰Q""5��=H�=Ƈ�t4R�v�bT��Bt4[�Or،ǌ58���~	��P?񞕵ޑ!e��[�E�0d���m3@Z�M��ݓ��6(�YY�%����*�N0�ݹ��`���U�%m.���xs����D��)��-���I�
p�nC�ăoz�5�P�O�bޡ�sah�x �p�>Uj��ctOi9晬(T|��;��|��5��{����=�F�r�J�Z䒸�v��?���Ǯ�T�~�dKE!�y첵�e�}\J)����ҢD���CTC&tm����&\�/66���N]6�xs��{0_��.Re�[�-���=�������Ŗ�pZ���b7t� @�K�l�E��Z 5ZyĒ5z��ë���l�O|�.��V��yC�%����1{3�7[��QĞ����8�������K��p���<T[���gM�v��?ZحՈs����G��{F���~��G������'�g� S��d��P��KH���fWԤ����3�#C�m��2,��!�\�m0�-�|U�D/m�/��P<��2b�^CF�Q0�h0,JZu$i#6$E����± zU��b�P���M���㗏��\���b�ka�b%�A\��0�Я�|�	�n=�i3��p�i��[s��p,���8]��	�BKɒ�A�A�0+92ӑXm�F|�C�3�ݻ��1;.]b�s�i�몤���R��Q��ĵhr򇖩���g\�s]�v�6]�$N�%��Z�ֶ6���Օ ���L��(���24�kWUk�EQl �?v�����-ݬ�&1���L���HQ�H]e�U\HZ�b�t�}��B||�����OF�����8�Ԋ2E�\�<�%X����Kr}�GA��_�M6�����0eN?��ibc;9�d@�j�iA�Z�W1��_�P�|⍃�r����i��h
����r�+�&�_B�xm;����%b������EH���L�Z��D߯�4�x��ǜFW2͐퇅UҬ�I�+1	)`@6�g�>Gq��
����JgB��,<x'�k�x�M];��o b�e>����C� ���?<�_X_��z��޾y��z�D� �R��*a�"
�!JקN���A,G�����֠i���~��D`8e�Z��ZAC��	���'+�$)''����*#3.�߈�V������VO����y���M� �ΐ�M��49�}�$�Fvnn�ų��_��z��j?����"ꍥsz���O�-�kU�V�<����h�4�&"��h,Ir�Q��yaJ�����@�lo�Mpr�X��ɰ;Uh�MY#�C8���Lr�s��3��Tɥ�)����.]��X���ĝ}?.�8�ԗ�f�tJ��	��D�l�<̦~h(-��G����4��%�$Z���oT�P�C��>zHf��0��L����.��ɳ����4�ٷsgH�3�{%K��� ��� ��!�����*��Uh~�c���F13�B�����t<B�XY�/�m?J	@kG��������ߞb?n��[�,��E� WVs�?Xc?i�j��M��L�Vw,�ߓ���B����/�\���S��?H��R�PGGg������mr�u�]9d���7�<��4H��� 1�h��_f��Q���Ӌ�[�qE�� ��٤�������q��~,�����9&���T��?�pM������Mԓ���aL !g�/��l�$$jG�ʰ�3�h��G�O�(����V�7l}}u�M����.�������#Ah�!�7�Ō���'�V��a�#�>�d���Y�C���[bX&���rv����%̃�:Y�}���K�B��0��.���J9"�"Xs%�
����V���82Ѐ\�Y5�T9�vLm�#9��G���ϸ��]�>����e�������v�,�=�OD6�=��|�K;��K��7�h��#�iER�q��Pu�ڭ?M������l|g�6j<�L�?<dcT�����_	3g8�υjFn/$G���N�<��-n�B�➻|��'��Q��a�D2������ێ��&�&�U���h]�0i���=m�?�tB�]��b��{Zt��}���)6�{�M�VT��2�f�ױl����͚��!Mj�Kd��R��&�u�[��,e�#��S��6�o���9	h+��:M���6��n����{������-��,�O�u�頟���z1�}������t�zT#��_mt`+_)�J�V{��=�s�2��^L�W��Umgȩ<S*�7IhS���˖�?���G�#��
 U��%nlnVT�wpPD@@8}F��rf����%m�9]�'�%�d��дR�7a�3F9?;�~�'��>̲k;��T�.�_Æ' Őj0Ku+�?,��$$Q((n���m��|���yL����q�A�k��P�V��Ïu�⟘5�X0iR,���g&���Mk����PL�����G��]	ׅ��V�MSs��{F�;F�99�"��4�Ҋ*6�����ȞRQ�����݄XO��d�-p��r�5��U��~��Yboj�{�u�s�j�U6[S����_�$ʾ6 .eb�8�&�9a�~�x�X['&��ډ�ʥZ�����|P�98B��Ij�q0��x����M&!@h��%���/���_�ޭzx(3�=Kh�5Uɐ�|� �^�C�=#�ޗK�*� ����3�4�&!�Eѩ6������v�Zg<�5j	<#��}���O����7R��P�U[``_֛k n1101�{��=�`l�{5M�CGo:4��CC�qa���6U���;��-����k\'JnE9������=�6��>���۹�T�l���������j�5��h�\k������r�{��?�t �9�Fw\������@�=�HO�e��L�@�t�`j3]P�!i{C�	]�7�Zr`+��z��[ѹn/q�qaW�� \�f��pp��8����g3�u��a����4	
����IH8���6���5X[��	�x*�&��ߐHJP��;�a��wBZ��s������iv�Y��+_3%Lt�!��6-/�#f'�h.��:M��R;��Q�~��K�S�jI��0U�yIU�B*HM�A��D'�m&���Z�"��T�f�q�@q�����n�����k>w;��W�*.�YY�v�q��м	K�����w�Rb�De���[ԡj�qxx(o��iU��ܜ��Z�I�����^�����-��} 1�_����=�8[�{�}<�Wye���m��/���*Hu���6�<�q�� �ʿJ���A� \��\�����ܹ����Msd2N
q�K�����PR0?ٵ���_��8[��6N��Y�pHl�if}�4�:���~��������5Ղ:̈*�����*8,�����3o�+_�����q�gM��7k��R'�@_˰������˷�.�tR ��&��\4�,�u��s�����|�f�������-��J���A;߻I�j#�yk�6ae�g������ j�;�@�d���K�+�@�<Q� ����[��;�!J�Fr�BB�y ��7��ݟb�U%/(ݎ�����������ϣM�l�?��&6b�;N��ܯN�K��S����4T��5I��>�I>���{�T���w��N�%A�8à7�:҅��S��u�
�ӻ?#����k8_P�+V)���������%1rtL��<�����UX'��C~ ���ű�B'�V������/�i�v?�c?7�n?Ƕoc5���P[����lu�N�VBq�Ѕ�/�iî�"f.N��&m�Ԃ��>�����:HGCWhϊ ?��w	��qnks3��ޖ�x���3/��A�S�v��/s�����O�T��&�Z�� ��[�r��FG:��q����L���,��n��+ϥ_��T$��i�Ujڤ��hI+wu)����:���jB�m6���4�pZ�"@��Q���?����l�NP����W[��g�m��u� ��`k^g��NK��N��_K��PN�^;��ƓX��q�* tW���7�c��������+�G3tY��N�3�t5��5����U�!Y�Db#���7��!��K�B��A@�}�짯R�{�[cɴ�e��l$� ���o��|��nX�X��[�G	�-������y�������.��R�s8�e��7���"j��\������HO�L����g]I�(�dmte=A�(Z��[�,H���6����O��O�_0jo-F�	wb���S�姐���D@8p2�(6�de�-�ߡ+ڄ@���I�=$zd,,�K�6SS�UzK�)��x�k�����zZD�-=-�Z[[-\r�*p���x��^<W��6q�kn?w*F��n�\�:��m,���/u�W"R^�PfC�<Zp!����L���m�n��Z�z$]A���->��N?���}��@���>cy�����Ȋ&#�s�/W�7�����Y��d1 W������oN1��4�o���/�3ԯ�W�|�s�-���Q��q�۟EC�3#�d@��4�O�e�U�=�\�m�="Ͳ����V��e�J���4I�*�T�j�0SҦ��ͮ�GP�u�b�	���ҝ��'�������Ϗa����e[[�pp��9���Wв�w��f�.׫���Kn�`��ƽ�E��NE�����PX}�`�5M�u{��*�\+����ADϙ-%�{ ��ܸ�cMC���V��~}�	�L4��E�.=�Й�k1�A��
����X�1��+%%%�:��b���Ӽ���q:ML�bj� �G'�����Q�`%V԰JA
�d[��dc�TݠB�� ��/�Q�p����눧>�1�NYmz]=H�����fw�.��d�t-EQ���������� ���`p�VW����U��2W3D��f�s؇�B�������Q�6�Mn뫋<�,v��Ѥ��wW���!H|l�����aAA֏�s�����/K�t�v;�����Y�K>A��i�KxUh�E�nD�}�l�4�t�Ǜ��
�Wlȱ����D���S}��Y�u���s��yK��fT��á2z3K���G��)���j��*K��A�"�����K�2�~�j�T'���Y״o�������K�����+Oې���/Cg����#L��/�`7���bߴYD�P0L�7f ����=��"x����0l�f���Z�i��YS=�1��<͗���ǾB���d�U�.㿒WsNϊ�����	��u�Wl�xk x�7!�z,�cD�;�Y)B:&�z�K�M4:\_�)����EzR��!()�	���;��;sr���Ese#�ٮѠ�ō4[,LH8�t`�lA*4��Z]�O<
�o����P��-���}.���%}�t)D�E<O�4,E������&�3T71'�oI�Qב�#S/?��V0$:s��܁U�=߃Uh�9m4~�)��	�G֖V�Q��K�֔
��� �!��G5��;v�f���~տ�,�2�e��t˼�Q/��H�2��5.&!�5��:u5��|���B}B��i��PN�Jm��DKsz�]I���-��Dy�4������D�^*q4]�~I����*��ۖ/�O�RU�E�������9�ZğȺ�{rܼ��-Z�\I�m�\_�Վ
-*�JA��-�ef�3hEԨ����eJ��.�u��a��\Ũ��oVkK����솵��� �OWA�%&�����ʬ�vؓUvuM�7ن�{6yGxw����T:@���|��ܷ��ܲL��gs[bFV��&�iOrkA�GyS6�Ǆ.y�;���4��r�Gw��xW0	\<��L��N��'f��܎�����ؚ�L��|4?f��νԑ,�s�����{$]|��qcC]�@�{�y3���'H�,��ə�i#�)O�qppz8�=v�o�r�f��r��D�o�RhJ2�s-ml�%�g���0Z ���ꐩ�_�����CƋl\\�2��_�����>��4�.��* ��� 7 � g��nR��4˭�V(�u ����b��>�J�Z��x��SQq|�hD@��}Z�Tѱm�&�L��Eݽ���*��Sˮ�Ě�a7�p�������MTSr������R���,O�������G��+�B4��2��Q�-���MJ�g������ylml
S3��^�-�ˇ	�fw�ڀK���w?�ً	��R�	gZƚ(eh6��H�Xɷ2g�&c����&�K?���_��v,�B^����/Q$Kh<���xVG�4Ɣ1k��yw1�a��00c�2.|���Q����/Z<|?����їH�]��vG�4wS�=#��췸͂���On���~�v�&B�48�/�����"íwh��jrl�����nQ�A+j	�:�i�ܜƝ13�G'Ət#�2@��b�&:�3.�=�2��۷��5|lhQ}i3@}a`{�����9�v[�Ҷ�_����v��o'Ǒ9�{��aJ��֮�6�*mR	�]�lC2�C�������m�,�%�}�a��Ү'ZW+��w;�s����v��}�Z�M3���_.��7+t=�٬Յ5]��*���o���64&�> 5]�{\���XWy��i.)�5C.c�9ʍl܋��)�����$H���a�8�<�1��[*3E1M�2�U�JA��#^�f\�kR)Gq"!� 4$�$F� �@>�q��\0g��&>f&S�|�c��kf�`�v����8/(��ZE��r��(St����z
�j6�~:432�b�:jh����fJ��L��F�����_<�8�2����u�5��S��8���#����byڼ�Z*�S4��)7G+��[!���Df��h��k)U*T���M��OMN�����,�
��G~do��b��eZ��������m#�#ۦggt�8��d?� y�!X0�/��)dɩ�,C��;Tղb�E!dY��˧�BpC�,��_�g��43Pf'����r�x�����w�<&;MwER��*�PUAWͭ��9�y$V.����@о�����A�F���ֽ�[b�q��r�d��[��r]����d�R�W��]���ommu7nܨ~�ӟjo�x@ǚ�X`�.�y+�Gv�d�8��KPd /+��)��[:���ɛo���5kּ�ל���4�*�o%�1���W/=u����}'?;����a�NA+ZTW�
����Z��󽺈�)�������r��d ��\��$��6�cb�"8�$pM��w����_�w�}_w�u(,��h�w������{�1̴jp�qE��� kf��5?�(��&�k����w��xvg3s�M4ͤd��A*/�y+K�@�ID�g��.�a�/�l���
�H�	������y�/�0�!�؀R���);�866���T������{�~�x|����ڇ�������q�X�MD�*�K�;9K3 D�մ�Һk�Rm)���_���O�'i��q�F�m�j��x�z>	�T��w�:rJ$���
|5hyc��eqb����C�n#.���Z���BnM�	����|7����{����T*'�h������������3��eW(&E�%_hNS���b�!9��^�Kd��Hg���,�@X Ȋ������+�+�h�������H_U���V70� K�>&���Q�J����mw�jג�о��h�
�*�
A�7��ƴ�������N����c�i�x�	U�A����ƺ�ձ���^�Z��r����hp�r���d`����oH�
�[I,�֜=۷���?;~��-& ��b`6sss�ʕ]�VjF}��Y�����M�P鶴�h�����N  0:X����5~��|�>�3Sp����ށ~y�W|��d��{ �E�;� ٭,���Bkgffڹ�8	�p��PϿ;������ƺ�㫦gg�I\�0(�aQ�3�\2��sG��X�D?}��h�K�����OZ�#��(�Lp�v:[!��얘���R����hI<����1��U���^<"�W�]���_�\A��0Y#|H��*r�x�GX��2֪��V��wP���t��E:{�5wjG2�\ۥ��]GMn�}�շ�K�9w��A����Ծre"�f'�����Q<E�i'73��"�����6RѤ��f���?JE�ۢa��yR���,�`}W�qvv� ���|q��5�����2 q���nq�����T��������
��.o~7>�OU�뷬UԱ��V��qf���eگ6�E�F�?�AύR]L)?��q�{�h��]68����b����g��y��<_	q�;w�t������O��1�3 �`�.2�� U���d�f��X�5ibϞ=�W_}�3����Q@�1�*�o�Q\�p!y��'{��~߉�mՂ� f* V�N�Ț5kXP���??I W�RyQ��f���$��ߦΏ2��Hzv�"���:|��Zh{�A��{������زe˾�� x,��EP6�+#�W[����42c������%(���`��g�bhh����?���]��@=�s-�Y���)��3(�U�v�b����<�d2)칎`.c. ��.�[%�8�5���G6²��2����:8��xp<�?l��,|@y�X�bf.O5�F��1��,��LM���R���2�3|l���&R���N=�멩��>N����|�&�|����@W��LWv�Q�Y�g_{W�32F~w���fjY�E�x=e�|�aD�Y��t�XXR!]�+���ܷ\!�����r�75Ԧ�ƓT�Z�����R��u><��5����k�(�2 ��²�]�S����#����1�ʘ"K@�-H��oUx"��d�\U$2�[��2'�b�(m���z�+��lW@?�J@���Z�����R����m�ۖ2n��I��ǂw���`ww�ڱc���/������f>@>�alϗ�-x�8������ի_۵k��===}�oE�
�[E��G?^�����w��C��!"�wc�R����f�М��>;������/(� ���Z���q]������zY H�*ƚ���E����<|���׮��_{sf��r����6�2]�b�H�*�ł�걱�,d�������f�?<s��x��"�{H���H�܂�
nyqSl����7�͕�����l�k+��v�_{Xb��LH��� LI 5��m&)�v���L2�X�d�i��,ŋ�>f$�a��
((pX���JXwgf種�Aէ��` �9��R6�FSQJF<QOe�9���e�b�~ʤ���ϻ�?~M��0m�^�^�ԦT�C�>s�}���]{�A�\����r���͍O�X)���zs�$���0�Ja���N�-�`��%J�N>��r�I�ӯ���u��֐y�ݸ����0z���4bJ�%_�Yy�l�]��T�F@vV�KYo�~��W���m_��v,�k_G�x,
$���r�=���_�Z6(24����@�ߕ���/6�Z�R�α�YǊb�`[p�f���[
.�_�k�?a�B�u�ֹ��w�N6��O�����|(���1wˉh�/z��7(�����c^�ݶm���^�r�@@��*�o1� �|����^xᏟ{������H,� ���)�K6l��ٳg��*�ɪ�S�z�xD�����멭�MF=+X�L�A]��d����0����jZ%�����y����������w���;�*sw/Ͷ�_Y���9Nx\M������(���ѐ����۽<�6H�{|��oln�@YHMzt�5G[�`M"�x�d	#8�Ԓ�¤h�v�~�(�}I�.�[�讶bY��t1c�~I<c���R:��o���K+:��s�A?=5�A��6�"���(��hff�Ǘ$STpy%]*�M7�+�5��+���_#c�*�޳�"mu����r�8e��ڵ��u����f�Z�Iz�W�����p�h�+�1UCa��NO*>v��A�\\�gs�s
T(˱o������ӳ+b���*S��(L��8� `}���y����^#"H��"Q��4�J
��,8U���`��]��bY��
�X�U�~����$�ߍM�o[�.���/u��] ��w_�e"�-[��B]��*`n���"��K>��I��z�/$�lAQ��Gmܸ�S���0�(xM�a��Ǿ�+q9�r�G���Mb���;w:�����x�oO�
�'�|�A�#�����o �2[�2cI��<�j���:�_?qB\�HٓɘfL�d`�M��΃oI�����鈆n%�&��/�'~���=p�]w��{�����a���`�h=M��&f�k���~k9��ϟ?woo���jҟk�b"�]0l��BJ4�>��{�]Z �'�,��*��>�(����biX,��p��(P�>*I��>��1oE�,��]}<
��3jxx�B�V9��K>�x�\9ˠ
�s#��r�Y*�
�G�Y7T*(�X3S�(��f�� F�Uhv����n�&�b5���~���Q�=���ʻ*_ti������L���qۇգ��Wf24=8Bwn��e�Y�D�c��옊��T_S�Sȗ��򘑵��
�A�P�	:��|.�-^HԄ��b22��9�h t\�$�#��QǪ���:Vi�X��#��k���8�-D���%uI�M����� �mѩ�e����yV%Z�y�e�f���Zp���_�-���^�k�k߀,{][�7o�~Z,��\CU��;�N��:V߼��.�DZ����O�R�}ihh� �  ���ϑx\�J.c�ڗy��uq[(Y���6m�ta�޽o�]��>�"�p@��*�˚�b��'�l}����_=�����5��c�FԖ-[t��s��ѹ�g�ٙY-0J g,�	Pgg'utt��'O��%Č��Y�3wMP>��WȮ�@l���k��[ny�?�������ys�`�+f��B��1Y�R��V>>L���s������naAn;ϩ�3\Y�c=��H�N&��Q�(IÜ��%3'B��|��*[�ȫce,PJ����hO/���R[�dH���:X J�HX��:k&ڂ�4�yn�x?��(u����)����˖-��p-�G*����(�'���	�W��jZ�FN��y�n�B9G��4��RMC��2�.MSݲf����R�g=�����ֳ/�T1G;��s���������}��{�̅!���������S��R�0E�9�yrf˱���i��c��0��633�Ʀ&��-�Wפ�λ2/�j	�..K2kb��NLL����w/�̈́�+2W�,Z�((�oV�/��O���;D�Z<,AضZ� �K�﻾'�[���6�5�꘿l�t�{W�zBĂe���}[8-���Ƴ�y_m�o4~�>�q�X*��:��ڼy���~衇�纾gP�>U�i��:d'S~��b,C8��ر�?677B}%���.wJ��橧�:�������O[��T�c�Y���X��̦������M�g���i�,L&hYk�.(������V�ZR#J�K}�|��� 
�=�MPl�ܶm�^��O���7�<���Y�jU�w�QpmD�+��G�����FvK������XS���6#X�?kĤ F0�7�=	,bpĢǫi���L"dY��K��@�@�SF�, ��%�j�TQg���t ������m�Y�w�0���%j��.��0�h4�NLL�5�*USK+:�\~T(F���U;=0G���E��ס�oi��e���0���h�Hm5��T��ι%5���_??5G-�u���D7GS�㔝e����u�˨a�V��'@&b��C���G�h/�wú�uy'��}7�3o���fP.i���fE��<�+�+�qF{���2��Ǵ���q�E�S;���n�*�;bQez���uy����>mg 7��xn6a�_�aۆ#�ܲ��"�Ѻ����>7;?��i��B�{�|.o��Gܹ�����U�h�K����.��g�YĵMb�*�o��{�����%���o}�p/��~�u���-����wM߼�_*����m�E_����h�}߹�C��WW�{����u�e#� �2O2��Ojda����Z��_��vCC�q�����( W]��XV+�=���<n?�1V�0���fs)d����.~�П;wV](ǒ@���	b��ɸf*���Ț�k����JRHC��U�P;}),\Lp���ꪫ�<x�[�n�,�=s�L�2��������{G�b�,�;�#���)�B�����s��#�}��bP���:&O2��F�\�?DR�|��G��"s����d��eM4jI�I/�	oRE�X�kzB�F* s��w�+�>滜���ꬠ���|��o!s����.f�;NQ[�ʖ�����K3�[QS�2�Ja��V9��&hYC�[�)��d�"�8�f�pƥ�ːhlZM� �3�X�M��C}�ґ_=N#�~��s��z֨u�����Ao����>���I�y�&j��YX�e�t��BQ���l��)�}ш���T�w�._C�����-�X��&�h�����=��h, X�%y����2��O��2�qUɼ��>w�ŒC�i�y�m>����Fh���I�i�[������オ��U�o�E�P���$��%h�l�I+��ѿ��9o��U�����w���v�K52|ߵ�r�uҗM��E���Ҽ���~�^s�y�$��k��Z�g�*������"�,�j3[�lyc���o1��	�Q�2
�U@�%1C��˿��խ��}�S��bQ��Dx*Ҷ����섐�X���gH���[X� B2Cf3V^,
�+�1a�@y5{�z�=A���Y��1����<�k׮��1mb����t�$��Y��*�{����T&�!G��5���w2���GLE����G0�L�^��L�"�����7.z��զ����Fi����L��8�\��k��~#�J����X�$����\߭�b|؇��o��Bf>(2x���1/���'ܸ���x�f&3�������eܙ�9��]
g@9QM�e��
y�,U|�T8N��9���P"�B|o�7m��*�fW}�̳���ߣ���[����XM�r��}�zᗏC]w�m7���Hj��s�43>Nu���	� >�����[Dt�����Z��|!� qC̫��$�LZ���\�Y�����Z����wpp�	s�2�=���M��zLѢ¹�~��Kg~���%2��oXV�S{��Ŋ�ի�Ρ�m>���*��j}���y�ԥ���K�/�C��m��[�t�K��b`�R����_�֕׎d���o��V���^��Y[[[��۷�|-���?���`�?��O�5�p� C�k��^WO0H�����_)�*�ˎ�`NOO�;v����o�槇j�&&Q�܈������ե�O������b> �"MtKK33��NՎ��u��~ɴf�
�"%ZzI �'�A�o�O�Lv�����n��M�6�V+!^C"��\X��Q��u#��ML �~3��������gϞ�oy�&�^G0�`�E�  <"4$�T���y�]L�+��R���$�}�d�1��0��0�q��;���Ina=���u�)(�qЀj�b����A����g�S����Q]]ZMOOͩ^�U���v�wY� �"�]+���q�<}��F�T[�LTxBLJ�C��sT��0ff���o�E�����R\�54��P�>M�v�T+Z���ʕ��C�3�ާ�b��n�B+���x=��{�+�|\N�����Fe	�����3���ܟ����|����ONL�8�����-�Tfrju4N�h�[�w�y��g���f	2L��;T�eooo-�dy��!�~���Z!<;tQ�g����,�BU��b�t޵�������1��~w�yq[�rş�b���,V6������*�����&m`�^^j��R�Q��f�vCծm���EPV��oi��'�K��Đ_y�z�[|��^��$.BY +�ӂ+�ݻw��_��(_{��J) W]��u�ԩ�����v���� I��C��e.��:ͤP��칳P�t��p���ܩ�)57;G�T�-�a�9������Mͤc��&ͩ�L����>s�����m۶�oX����J<~W@��"����a�:cb�{��/AFCw�ξ���ϝ;���T�2��b��$B�J�Y�L�R<��V���`�a7�^��z��ۈy��m�0G���bi�?���>s}<�4~��+uޤ�_���u��Z"�y�.�����J� Z�+�����6�)d\�y ��D�m׫dKJ����7�@'F��j��R:���(�-�
�C���?j�l�jJ�;GEF�ϖfjlh�T]-��&��>E���?�s�|D���v��B=�+�{ެ^>r��x�!w��U��.m�y%�d@v~���_�eMͪ�����xt���I9��J�T*���Ln��~�,߳�<��o�|�X+�3߿���>Vi��`�Al)��fnV˶��yBr5 U�rU��bQE�wd�\��%��۶۷��k��2�]�
-X�O�Yl��6g�XI��"�.���.f�~,����.a��궸���M^����R�cmo+��w=��2~(~ ��:�}��������H�n���0����m1�UP<x���۷��|�� ��k� \tY��;v����_n�¦Ўg39*�`�Kcc�G���<irb~T4qRp��	�l&KƍIa����P�'@&���Pe��吙X�ϙ�я~t���o��Uo�2����4$Y�|�.Y`U�
DV�`m@_�����������`�����F`Ł�Y�'�,��HXEcI�%c���3��X���6++�^�%`@���V�\#`�1��"ׇ�ދ�I�..��\�;�w	���hDKU9];�E�m�|��k����L6M�L� z�N�B�S���*�Qm��r�e��|��Q�&␤6��T��(���SCM��GU�)�{_��M;n���������g?��.L�о�W�U�{���k�yuPy�5z~Ρ��,��f�>w`dH�2���jkYV����w�Ǘ+�#!��TReg�x,��~��v�p�gY ��#�s{���f��Qv���"غ����`���Z�lj�MT�Ҵ��?���>�?���n�g�!��mKH�f��@��R�W�4��g\��-Ծ�>{��_�>϶����|��
��
�kP��ݷ��o?_�=�P_}J�8y�� mWܻ�������h^��X P��������#P@C�j�*Դz����M�t���) W]6��`�;�s�?��?��裏6��A�Ti�R4B,fiW�t�^�Ck�@��L�?$���K�GZ(���Z ���B��u�$A��)0*/���.�Ba;�miiy��{�}���~fϞ=��R�3��ɓ'�����ٳgu��ݲV���?oI��҉�[���CCC�����p||<m �^� �@ U�H�qd���7q*�⪼b�:�O�m��Q�w˥G@���6�Z��,Z����}*���|�e�ˌ '��-�!��X��;,�#}n��v�3	:�|�-gJ!�o���X�^�(|��  �&`��AE�9UCW��Y��Eʺ�Tt�ZI����ǒ���T��Pm:B�(,d��Jt����w'������M����_<H�����+3�5�ԭ��S��i:��4�����<m��jii%(`.Q��R�'���	��%�@%��6� )����l��]��&�|?������X������GFF��b��D�MQ0H�2��98��[ЭK,E>�❷`UQ/5z q�c�����N %�(`,�j}_��h�1|����r��6U���}��_ �ʎӪ�(��7�X��X�ߋ��J�7�<��}����,x;<ĳFx>x���MVI�w��rͰZ�Mp���S۶m;����_2�k�5P ����h!U__ߞW_}���|���B��P�ʁ�(V�RWW����"�pÚ��,k���p�;`&8B3��������A�r�=�d�}
m���VE�]w�w�q�#�>!��eB�׵v�Z���YL�n�d� E����Za�c��ltt�:��-�],�9<��	 � ᾊ�`ssP�#a4E�=M#><���2��yA;iL�> ?�X�ĕ㝀U	s>�L*�*��\Cpm���b�'uU$�&U\ˀ'��0�$qOk�c ��6�Q9_\m�S�@a{�߹SC�:c`�ϩs����t2��ġ��s�U�P	Be�b(��*�)��')���s�n}1��+(�eh�Ń�X����i�u7��bu�XM�:�䣔*��=W�SKr]۽�J|�^~�z$�Єr�]�^��-o�Q��ީ݊�	�����JTH�Ec:�\*�By�yUӅ������>����i�/N ��>�ϱ����?�wr�����J�K�� ��-,�\ͣ��a�ϼs�`̷�2���m��7�=��:�S��P�;G@ռltUڹ��K[{,׹j	,m� ���8pUV�?�������-:gh��O�������X���-�3Q�Z���Lfc| � y�Q�)�I \RP�0��nݺ�����O��9
�k� \t9P���؏^}��<��ӑ|��#��4,���f.]�|�
�����rNA9�����Z�
z�M���&�_�&�lv�L&T��,�JRe����gS�^y��7�t��}��}�_V9̙q:�.H"c��߷2�a�^��0�E��So��9s�>�W�`FxN�<�;�X4���*�iw�\>�x����)���,\{�4��=�ی���8��*�Y���`.��7泤Sᙣ�1��X�����C_� �@ ����%��+]נ���L+!��@�@���=\}��
��;}���t}=�nH���Y5����P}CZ%jRK�PM2�S��9]a��#4UN�k��D
a���T��N8U�2�QE7���TüB���ܨԾ�i�6A����>G}�St��1��r�{�jKc;z��>7��G�h˾]��UOQ����D��5�T��#���y��2��b����k�驌;�;�:���iC� E�a��௅�����737�/���^q�ܹ��e���1��F��ʠ�ҵ������Y�g��<���#���2���)� �'����"&װ�X���h�k��|��'���(�.�6���c�Q��/髯��w+�����e��Y}�g5�����T� ��M2�Eh^vD[���U{�Үx#�}�~	��s�X+�^˳��jr/�����P���\�q.��?w@}�)&����C�v�z���0��Q ��F	.W��<�Α����U�q*aiv��pD��lY���ڦ���@?�?�KsHA���6jM��
"��$�P��Q�5�(i�+�T�Pq]�f͚��s�K���?��.;�����m&H���4��7o0x��닐��o�p�(܆9�@�U>��&0�jxA�(�Xt<���_w��km�h)��L̔�EW=�-%n ]�$QP����U�w@[��'H���c�1(ȼ�X+$�@�q���	$�A��dmm���h\Ml���c$�G���&P�J��VV�HT�c|o�zPd�,X����>�#&�7���Z��d"����0��J��(���F�� ��*:R8�>M�nu#�u4�SϽ�FNW�|�Z��C�֯q���4H��J;��˽��
Ka#6b#(���$�)���F�Ox���LLwOx�������'����vG��cy�-9$�Mj#)q	 @�@��ZU�}����K��{n���n���`2+3߻����;�|���X6����izi~������][�P�-��T���p�)VKs򖊉��9�;qZ30��;���ܺ����x*�K��G1��1�\D����a���N�O|srb�����_�Xm�R|pnXP�8e�cb�Y�(�(�,Lu�,+#�'P�C���z��F@"��(��1�l�@f5� "c��=�'�˺Ɔ�j�����]�=v�����.}�v�܈m�Dr��ꊀҰ�F'S���_u�l�bo
�S� 3�&�\a ��u��?�rn��s� ��c]qVޮ]��0�Uj&���&�j�ϭ�PH���?~��S������w��q�$=��Ʈ�N��󈱚���Ņ-t�||[{��ɤ�:A��pG�	�\�(�͂�� 0�Pj!� P~���yW'֯_��2z�n��*�O�8{K���3���O��|�
�����a~�3W�@�X�F�Uʸ`(ì����W����**��ļI,|�\�s{ʴ��A�TV<�Lnc� V,���v��C<�y�xq���\�4��\�p`<�ox���*�H<��_��������Hb����@A=fGUor$5e{<��Ī���X����޻� �W[&�������q{յR�/勪V������T�|���mt,Ӫ>��KT��C:�ww��z��=K__��~~��ZV1n��j�6l&���f'��Ս�z[Z��M���#4��m����A�
>N��r�]�������՞��kI�=����3��I�(�+��?�����������<�ϸL�o�D��X����;*�V0�Y��7b��>����2�h���o�m[�lk��D֬#c]��BQ h[\B$�m�1^Q�����8X�z+�kp=~t|��'�Z �7�~T�n=�:vE��U@lؾ��a�vrwa���K�,pv���KL���C��������w��dC�_G1�\.3���޻w�ٮ����|�ݖ&�j�ϥ��qY.��M������u�d�U
H(���Vr�֬�yr��!q S�X
2�Q��j|�}�6��`�֍k��'��ʦ��
3�q'Њ1�����3�ǜ��>`���M�Ni\}�`��mS������`mP�"�àb����S��?��5���zv\ ��ɝ�"������m-�-�,؀���@��X�po�Շ���
J��,�&�P�{J����ɳ�z��Q�/���(����q׏��522�c����81�3�~	��ɋ%;���2|�B��wƵO���'����b�^�� �K,r?|��7p�Q��VD3 
n�q~��5����*�F=�S�#K���D[������W�s����Y�k`����Ok�����	:��Oijv���'Ԛ{(��M~ѣ|���s���asU<M�K<�{T"SK�ONn��/P<��jo���]k����l��� �ǧ&��������fc�5n_�w�d��zB�C�`Ɏ�i�^��T"Ro�K�96b���b]�Ҭ}L�U�(ب}@Q 5�`��sC��	߅�gY�B9'R}ަ�����V�H	ۗ�7@{�5����¢e[� +x�1��(nܲ���)��Z@5_{N�rW�u�(lbMNN�7�|S�mC�bm21�6�}�����sϏY�_n��}i��f��g�TZ��Ǐ��_���Ǐ��~	jk(��`����.whh��!���
��0���>����@�Uz7�'^Fa�LIA�8(�`�B�	
@׆����_�k_��WN=�䓷��eD�,D;��۔F.+�XM���E,V333\�)/VC���b.��%���?���X,e!�D���U�(�3�_a�ĜH��Qp����o 5����C�8�V* "�g���Cf�]��6����.�l��&���K(=�.�H*lz��R�P��3��)�>(��I�Vc��V8�^9Ǹ5�L|ʠo�F��v�Tx�kP�Xn0T�+���e�/3�r*bJ�e�o�6��-�7"OG��P/�?G�r��޵���R2�%��z������p��v�?@�M~4��T}��]G�j�/�=�
�����ylr�˾����tj�r>��d<��fZ�Sw�/i����[���F���\���9�2)�Ē�#����)�QK��;j�o3��Y��Y��9��z��Ê"��
���_��1�ʺ ,;~G�ÊwkIؾ�l�c,R��M��-�nR��c�8���D�[�>Y#��%�%
��F��Z��-3`����i���8/�B�^�m�I���Ľ���i/$>uꔎÆ��.�:==�2�*8p�Ԗ-[~�U�P���K\5�gZ��^��������♧�v���*Q���4�~���߯��I���и�(aF�}�!�(�85de�ZR���{)�#O�q�u�ݳgOyǎVcw�u�����h�W)�"�P�Y��������0�o͝+��y��ѡ�W�~gbbb;.b.�{��� ���z\��Q��E���es.v(\wh=��*���7��� Y�
��7/�� @"�b��+a�D:�r	Va����r�����<����D�rI[u�3 .l�����K�?�����t�/��
�c�����p���[0�h��RQ?���@������@aV�4��v������Y���W�k���_`ŢR
���x@�Jl���o�s�s*��lV|����t���;E)7Ew�Q��td���M�/���tKu����u[TkWU�r��Uc
u�j������iϦU��E��483=�@���,�r|�N�i��N�o^�fG��#<��~}�waq:�o)��a�
x,V)u�_��d+���5 �+��"
,Y��@k~��+�e�j��w�M��
��E �uZ֒�*q	��jԾ�f�Z���b_C��\C�`\>)�JE��kP�ZߢV�qa�W�z�C����@�|0��/9ζX����cYg1Nj6@�+gϞ�^x���c�O�[���sg:t��{�}����[W���J\5�g]�־��_=���>�Jale�d
��ģ$����ҙ�VGGGu,�>��Mqi�UK��!| P$NE� �o���BjbA�P�Y�K�ڵ����Z�˗/�o|���[X1��+��c����+a-��X�^\&�5�ӥ���Z@^�Ơ����A��z����-�`��'�z�I,������B��P\�0?ŕN|�� ?��m����X_�o�.̐��Rer��D�����t@ˋ��M�q�Z�
����������� R��R*n�I�C�),�}}}��UX���jճƇ� 0C� Q�]Л'���_~�3Z	ܢ�!�������1�}��݁��u�1ȋU+1`���5�&<Uu*�:�K�}����&����Cz��	Z�i_e��J�#=-j��st�����_�&�۾��3�����uV`���r�f���U��Q�� ��y�J�����nW�3�Lj�/{���:�.�����\zxrrr��C$�։��B&�*���$��ʱ�T�Ӑ|�>ƶ�����GW��GA�l~�@-��]��C���l�	�=���?"}����[��]�Y���l (�?�Ju���%� $���L���IY�5Yv?ɚ����_�U��u�ֱ7��')<��ʀ�pNAvXa���ѣ���OCCC�#��2_����>�+]�������LJ\5�gZx�\s��s����?�bb2��	h�@w�+���O��x�"��L�!�������O�p�$md���+�+��]�Vev�`	Hmٲſ뮻|�'�B�������1�>�J�p���]\ڲȡD"#�}�;�,��������٧�o���bAc���5�UK6t��|�BA�-+�(t2m�jZ������8�PBAV0�X�L<��s����$�I���f[k�f��v<78ƀ1��J�Vh�˸���[(��yzzJ[� ��v/�--z<pn͐UḤl��)��ӣ�Az��?��R�>�>�q��.�8+Y�WJ�jT*���bJ��ÿWݘ_�ajA:�\��|�5��P�,�*%i��kWw?�8���u�Fo�|�
��o���2q�j_�^�Lo<�4�#?���ar��)��à�\,Q���tTK*�i��9�[Z�Ӊ���̮a��po__1ٚ~���"5�OU���������E��n�9��|��"ϭ�1nWB�p�rӤ�Q�)�j�5�:6t���k�[_[�V(���Q�����җH]!�{��q�[�b�j�-��H�W�5&�2װ"DE�K��� ���m5��8�ڈ����"��n��`��w�1 ^u��fh(S�ͧN�pޅ���㐡���@���v�1��>޶m�s,��4��gW��Y>���{�������?}����B)�SP`�c��o�@�h�E��n�����e�eknnV�'�P2�}�����bޯ��ڰ���k�&�o���|�ԩ�O<��C��`��L�~�AɆ����(��h�|*�
��M*���Xq�gP��Y��G��E>(� ,Z 17�&������ 
�1)�^g@����\�梸

���O|��#����J����פ!д� +(���N��b�X�/�D�m$9�
������RP��r�<%�T��cЦ�P��j�.��8�&k!S��t�L���ZT2g���S���+">�Ġ-���m�W����|9�R��^��|\�\�����`�B�U�%>N�]�C'*�	|�~����٬���Hu��M�߯�^�N����Ryy��������}��z�şыՂ���O��w�$�����Y�����ު�f��)����*Ų�THU������[�[��֭�d:	�x��9�>MI��z���?�g�2��n�%��nk�v��X���, ��Y߯P���ڜ��{�m��R3�1ʰ֊�ۯչ��Y�D�X�8� ٰA��cų)�ú�MT�h���w;�X��%���ʔ:� 빀Lk\�$�{�]��w��vc�I����4�m6N۶�c�Nc�<}���k���=�|�\y?�_5�.`���7a�V�W� =�/�N�5Gz8�}H�kO���p�&X%<��/7��	Pi��qA���]S2���?'&����΄n�J��	xݯ�wvv4KҘ�����s�{�N��>/z>��_��:藢*���`?�|��:\�uttUTT�f�e�b��᳕�]v�VWY�ײJ����~){��5����	B��/�0��0��lw!{{��
�����@@~j�?h���{xSS�e�p����f��:А^���=�i760?�;L�9�E_M����&��%��@Q��6j��Ҋ����}�guR�\�	o�@�)C�L��U�A-{�ǖ;𽯝���hZ�u�'�\��'�0�wM�X�~�ĤN�*i�8a;�cc�"0�l>z�����AhR�����8*1Ҭ�M���hO�-ƍh��y���̕�ЅĘ�g�;o������z,��P���A��8����e�o
B�L�V3��?*�X���Jo�~�\�6=�Z�?�]�Ŗ�m��꫞8�j�/���.5��p�[�<t�9���S#=�E���D���$�֖��Z�#U�)ɩk���Zr>�`�x��~b���m�l��3�!Vy��������X��N��!�	�7ET�Ǫ�V ǳ���o��I�d�>c1�9�c�_�'�FY�hx�Mv&�H���A.��G��g�-�Z�_�ϥV��	V_�������J�O�� �F-�3EB���T�Ȟz!��7;��Ez�f̱n���m�Q�WV��cI��I�|c7�@�,�)��M��e0��pm��./�ˎ�n���t󲓔��?�׶=���?�e�mg���,����z�5&������(�����cՄr�!��u>%HN���x-\�vJQ,��`��C��L㽟!Z>�|?� �'�uoO~��pA���-0�P34Q��K}��hG7����AV��-y�}� /�j<gc�y�qo�Ś�o�L��	N�(�.��� ��`�
��sJc�U`|�{@�`��f-C��k	�ч��`C�`�(f�ی���.��L8�����C)���8 �N�a R�C�hKv,��SG���ư���Q�����'�$ySG튒��1���qo����������C��7�E7�ƕ��ܥ؇��$��h~���R�{���(�1�h�ʢVȳ�5��ҕ2�6��vD|�7s���e|�3�jEo�T�]�����������6U���%)�g�M��/`�Vvj�5�Gw\�~f����m)�RG̰�D{
I��R\9?+��]��W���5���[�	Ѣ:�������M��������oQ�:�(J|K��|�ge{Є%�ؾ��q���*V�����d�l��26��ZkJrE�/�3�&,d�^{�*��6^��M߂��&2
�.��6��f�U������" ii���6FsY��f������7�NDq��s�D�G�@ZPwHf�۴��T��l:���'~��?L�����~3��c�B�~�8L�H���ѫ��.��S���;!�y�,/+kd���AK)E�Q��[X�B���T7Ud�0��Ê}C`�TJ Ya�֩a���#���_+�S�h�����n�-JK��6{�/Q�'��%�x�&z�lw9��5��>a�E�u��Ĺ�����r$}4���,�eLR�&4�����1�T�(�MV�\VSFy���XI�J޳�	
���ו��4D�x`�y�B�*�y���8������y�	�����W	�R	lg�"ѱV�>?����t$_��O��C�U�� �Lu��+�k��"� ���f�g�Qvӆ+�!�Qf�i�V���3�d����A/�t�|���99�n��8�����GQ~�HbB��:�s}�$F�+�V>.�#�n�d�`{�Ɛ���6��� ��b�d�*�h�$�J�u��}u���K(��k��������G�v�tR�"[5�f�Ѫ��a����0گ�W��j2x�g�:������A]�,����/�Ɖ,�n�-0/RRm�Q}�����34<�s��������D`�nRe����Pk,�Q��	_ؓ �#)�X-��+=b�v�G���b������5��������F�h]��k@J����W�h?ļ���8��j�t���0&.}�R�]V[?���oB q��n���@н�A�{XS���Msf%�h����	2X�	�'���(�Q?�:�Ŀ����s9�����/8�}���*8�W��$>Ok>O㟶�Q����Ѿ��L<��
��V?���B�TP�����g�=����,�~&| s�,�z��pb)��y=]��m��@��t=�u�
o��8ڕ8���!�>�	AmCb���>j�f٧!��6/k��P��Dp�<]��&�T���E� x'
RHdp��A7�O)��_8�����=�@�Q1����Ԉ��B�����CkW[����U��]��/)1I��]�f]MAy ���bI��.p_����<twP9341]���e�m�wFA7�w�$Z'��}���+C�#�{d}�mD$؜b����1�*�E�d�J�N�O����bޙ�e���K��`�/��18:��/F,j��`51۴*�����TZ��o�]�s�bz��62׈�~�D������J0u��H�)_<m)\
���-g�ŕ]Q�jA����٥��Is������2�LT��*�琐����K$�6�3/�j�q������σ� V��-{Z�������(<S�������!;S���~�![�w	�y�0.}/6@j���>ӝ�6�U��|���t�+��pvk�M�������$[z�)6Bw�Q9���K�֍_e4�_eO���ꅸ�a]���E}���i�xQ��L��͍�(������P�]�+A���A ���x$jz>ۿ%�EW��ʾ�
|�z��Kl���ce#�)���T���Q�L�����79���d�ί��8�h$ֈ�<RB}��dj��
�&ߏZuě����:4E�K4�����Q�����?��.K6;ܬL�Z���90{�A�����������`�5+��55]7�J��x2��J}H7�Y�<��n�x��ĉ�&���~�TӴ����5*�� ��X��<����$/��fB��0�@��i!$��b`� ^�]�e�Yʨ*�s�K�)Dq�&\B�� ��c�Vj�{��#"�{xo���mCnU/�����iM�D�`��.U�ǻGT�	�@4%�`��"�!v!G	��!�����$n�Ů�89+�#-�TD\Q97\�e�t}����7@e���]�5K��7��R,���ϩ��4G��Q���|ټDYm��6�BE@�g����;d��ܙ�MQu6)^��R�{[���V�3�
֟v/n�����4ͱ?��j�[�^'���S �`����}���0+��0JJ��v��X�޳��B��:�����4����� w��<��/g2:�߰ ً!�[�<�l�7+�S��|��榪����0�:��M��(�/J�7��,lV�+���g�[��`�������*�H��=���lQ�%M&��AP����c�M�+�tq()\B����EA�p-Q�my��횇����T+�c��|�>XNg�-U��uv���3%O7�ϗ,�0\�(ԃwܽ�������/�'�E8�ï(ێ���������7����c��J������|CA��T��ٵt�&E�����(����F��C�k��Af�AR�����n���7\�vm��@� ���ds�$m���Z̼g��)������i��-�Osğ����I$'�;4'$�[�^1�#������)y�����y�\�M�wy�Q״�.��2�*�.��p���8v(�G%�iy� ��'��4���7�Jl�yr�� �)T��v��pwz �G6�39V+���l����4,��A�E���r�"�'���l�\v=����He�e�1������Ќ]{+���j������An��,GC�k��W#���Lr�Q�~Y���DC�{IOR4����� �=8������2�E��7�щx��y}�vlJ�$Q"v~�L���p�u�Ku} w����b�Tf�y+�8�f0��A�lۦx[��6�_|诣�,t�(���+{b���P-�Cl]�����e�C�*�x2��ꎊ�&�9��GW:����#��o�^�� ҋ5��G8Reh�����f%D�D�{fډįo�RFfҘ�RX�8��>XV������@���7KT۫��&<�WZ��ٝ��-�%6=�M���5{Β`�e��&�I5��P�Ѝ�l�f����׾�:�
�Pqss3�N��^�I��d8d���ۭ��CW�� �q��W��׳��@�Ev����ڔ�\�������M.�[)���[�`_)�$�E]]��2v���/DO��<�v')t�N�񸣤n�w�����~��y���s��G�<g��Qo������0c�H��01q� Zk��	>L�t������A�U� �V����EВ�UQ�9�G劐P�&�Q�=3Xf
!g�0�A��wZl<�B�:$t��F	����A`b�r�=��ы}.A��h���!�CqN���?����w\)ȉ~���軎��c��MQ����?���{�=Ow�b�')%$%g��O� ՞�ͭ��t����p+� ����X�"��$��?Z:e)�Քp���U'��.#���1 j�� �����]RԷ��;��ֳ�%��%hc��4KI�s��˫��a�^f�n0S�h��o;�:WW�7�h�������p����K�Z����M�x�~�T�_pX���7G ��;~���}}�M���O:]��*�mk���#�������G� �m��m�9��D2=��;�'��\��iSs����f�%/0�qH?D�W��7&6q(�
T��`�3b�n�D����jq7��ij����|~üt�lN�{E���E�W?�~+1�8 n�̿uj������y�="c��[�m���r�b�aDn{��p�)qڡ���c��yg��r�v���C�{�96���G��y�4+=x�X����q)�z���r��4�	�\N�|Η��]q�&�����6��JII	���r����u��u�8����Ze���y�ӓ���GD:����&����������W��_��V�t5P�i�jZKG��� 8p
�5��<�)��FZ�wg��|�?y���xXO�|*�������TF�u���|�)�w����:TjƎ�F��z��c%f��~p��H��ZDD�~������.cͩGr�0�^�j�����E����p̟KnIx��Dr��+N��=�a}��D�Y��p��BuۣM���Fp�M�QS�ӣ�@������֤J氶P���%��S(��| ���r�z�Џ�1I�\
�_ vr��G��ZVF�r1��LWE@B��M΢*�_����3v �-O�����wt6J�s��Թ��r��m�:}wLܤF�F��J������ۥ��s��ƹϚ�I�#���*�t�A릮�v���{c+y�����@[A[��ە�Tlx+DC�%Uд)*f��\ry��y*U5M�VI��;��ƨh���ҽ����[�`=�~G��7JC���:���Z:t��D+�Z��(�{�>�CH7y�f/u�\���gAղ�Y����5[�8���c~F޻7�Vn��Ӥ��p�:0��=�f���{�ʦ�&����aqO�,�������Y�f�F4F�M髥w+�����8\B�]�#���1"X�Ě����)���ˆ���Ӈ���� �_!!R:D�JqtãO	�L���B�s�3Е��k!�\�gE�̋3}4���� ��1���5c� �q���oÎ���l�������U٠��t���}�穁��?�Ì/j~z'(�)6xW�U��������kO�|-4L�m3��*Ki�	T,�3" zZZ`:/��a�q��P0� >�.��k��~��!� Uovw�/U(�����X`�ND���4����v@����r
c�_%;pnn*�^�گ�ߦflڝxYXP��,h�z#�IUз�2'm���q��'v�>�͖Y0�B�51�yQR%ЌC�	 x�����#�*P E˖��c[�ԧ�{�&�?!I��o�ePZ 5&�0�#� 0( ��������d��#m���_�/�=ʣ���ζ���-�.@��k\,�U��, �k7WWWHY�x�?2���/�ʈFk�ܒ��F�fE$+U.���7V�4�U���ԫXTKU��Ł�9�]��߱��jú7�g��7���Z��{�Y��3_�-�*�Bo?���DeIYnuݶ��nxu��K8��$���m�J��+�E�G��=�(��������,���7��u/���%z�7V^�V���p'��=���Z����={�m��v��l�]���-FH{L+[���p���8���^���}����nA�V%_f���ͩx��ϒ�F/ZѺ��Adc�I��{�Pp���W!��n�e�iVVlx�6o"��W����k�Z��x��h˵�C��8H}6?c`.�G���@���md��S6��4jd:q���W���6�����â��6�Է���xS3˯�쫶�짥j]��۶�/����}������{���ݧ����^*��������#ȠQ�-Wj������l0��H=�$�B�!�@�L��ɞ��B�U*h�Z��r��z�_к|n�h��G/��G�p���dff�ˠe�\;0�$�U>jA|�wCX��	�<,���r}�`�g�����@�/�@��+�P�ֆ� ��c<�=O���M3{n(z;L��)y*Ew8d���z3��Cڲ��]R���V�;H8�@��~`�S��3�gN�|�t!�PT@�����o��I�sĕ�v�3g���F��Ѵ� X(���(A5�;���
#���i���V��@�m�Ӭݛp�Q��W�f�^�C�9�ʈ�,_���W��-�6
�s_y�Mc2S�AB���&�j)N��m,�4�E9�ƇeYefks�K���"-�e�`Y�M��C���������~����̷�;�v����o=U�*L�^�պ�J��<.5v%��O�_*u��Ǔ�Sg+�)�kO��jY����ѱ��MM&�f�0ߔy�&�=6�Dh֐j���]�����d��s��/^�:�ɮy��d�H�|�yZ�Qe��\U8zd�o����#�ϡ+�u:�OKLJ�f�d9����������*�+�E3�ցw�v��:Wc?��@R��&�t:�x;w�C۶�df�-gMUQ)ER�)�����W��s���U�BM}�WY
��7�B��f�T��]��!�%�2��ly���Eɍ�q�cd����ϩ��6�OsY�h��?������}9�����f�ڃa;�����**ƍM���e��iP�Or�C�Y>�w�k�L��$)���`��`q
0��L�l���m7C[�<~<E`Z��Jw��\sج�xʺ�>�-���:�\� ���5Mģ#5D�UD�?�g�������8i�2����B��8�r���!�~|�Eh��2��֡����~����$t�ǃ�؏�9g&A�&�����t �S|"����:4��KR�1���G��������K�+�(�FS���7�����Y�}6�^�l!ǘ(����
�m��S���>c�	\�\��mE4+2J퐹m%j)�(3ע#$�Di̷��1���+ZqvuD	X����L�&\T�"'q�%��"��J�ӭO�@��Ȼ���,�{Śӟ�a��.|���e��:�e^�Y�{-��E:Sz�yO4"S��M�y��p7�����K��G<�)���	m�9���U�TΠ��Ј���`�}S��cec�ȹ�p���jh��G%�?o��#b� ȥ��8'�jg�U��D/j�݌���d3�↿|Y�5Æf`�E��J�"8�|n����0:&
 izЈvm�6�Tɢ��. ���g1�r�Q��~Eo��ӵh�}�Z 8��u�,��Oq�+�2p隋��B�Xcq�?�$���2tZ��s��5�/0=��M@E����g,W��=_)7r���V~n�@	a�[O|����S��24c�3���!<>a��ew�i�Y��`����ǝ]����`����F�5�@�Oђ$2�(�(U/���]gL�������z-���;�0�S4��.6��q>�jΚ���e��OA��3$B��&G�@�w��r/O�K+�2�����%�&�h�P�Qv�_���N�K��!p�� ��r�����}e�4�!�H� ����.@���Y]=������*wq6���},L��|rb�<�׏�bT	�Ā�	#�j����)���+�]�yT>�vlޤu3o�	�A�Q�~m��93h�R�TI������]:��N�����/��o�*�i{�7H@Q��	��8mG{��@-��ۇ_�MI9�F��;#%
��Au��C5�myVZ�͆|mC��:�'S��F[�g�MA�b2
����u�V�v�~�=��L��_�ǃ/V3�g!A�9S��<ŀ�a_���ְZv� P���Ƃ��^Ab�Ek�(����>ǈޡө��'�� }]�po�NE�	��s��������'����&̪�J.�\I�1s`��C��D��@�l�&p�*.���/�1=eQڅz�]�_�ڍ_�ڷG}��r u]"�
9��?
���d]��E'ژj�~�#!\�|8ض.��'J�����d@�LEN��c=�*���YK�4B�_h}��)�yO�t�{8��C�p������x�X��\�+`��*��Z�i�? ~��E�����<~���
O9|^����џБH�}�!�8� ��|���_�ֲt^Cܹ�	E����֯ɑF���?[��M��#s��Ï����������$�[<��8���-��t9��a�t�����>
 ��J�2�o�$a����Ô޸���������4��G�$a{� �R(�U���TJ���HeNJ���*�+À�1����Y2�`R �V����ƾ�g�gk��,?� �Ap#��]�o� ���Ӱ��0xrb<�o|O��|��g�Ǝl���	1E�6� �<>���	.%K��tWgR�{q�:�_���3Z��0FJ���ݖ�Y���s׮�6J�@Gx�|@D��I`a�x����P�8�ЬY�XӤ��NY�J)��P�Uf�\z���tiY�I���a�:Y��s��.�t�H:_�\yVl�\Cq�v�a�\� �g�ZV�N�9��,���J��ɺP�zI��~O�w`��ӾR~���iX^�pysXjـhc�p����4�~�aUBnc���uȗ��-B��G��s
�/����Q�S���.&�C�����il�=�I��@V:�Ƅ��]�H�X��RR������S����xP��e|�H�`�ɵtSv<�I���1��ے�Q�l����mR�ԃ����]Mq�%Ə6E��_��p�O]��&�Tvn�� �{�7��U'�] ���K�4���z��NPϾ˞O�W�K������m��������&���7�|4��Tt,�
~�9��) ���e������V�_7h5~Ī����y���p�M��k{M@& ؛
"2X0���t�&|��b��S�<و��j��ԏI�� ��T5�B�oy�tPI��X��+�H�K���X�=�y��T<?Ko##� t�[�#,��Ҙ�f�$�<�Aݦu����I�]q0ώp^��o�t�ah9�F�ݒwo�-��K>Y��+�L�L�1�x���
)Աa�����+n��'g@Ɨ�pW� U�o|�L_,��|@����Շ������ ~~U��f��;�)�F������K�A̺P W��m(�征
��L�l�6������Y5���nJ����vE�C�zH�;��W���2*RT�(t���+qI��=�xxk[!BZu��W�7�p1[�t�P�ޙ=ޯģ�� n9�[�;B�ѭ�n��d�+d��+�F�+�+�T yD0���^�ht��Ę��\��:6q�Y���~��A�t5l\����fC�3�F�i �Jr�x}ؿ��"���H���W@v��)��A�y�r}~wFkL���qq���E$��B�fn,2���
���S�_Ֆ|	g��)�z�#.�������^�Uc�.��^��_kH�#���P>��6�h�̍���խ��+���~��H�|�`QD�Rt��v�^�0�?�]�����R�3i"�J�P*كo���_�?�w,>��5�K�ڊ���<���+t?�F���0�DI�0�/���+	,��-��2���k�|��
E���Lٿ�^��ԭԆA���g�y��}��]7�0d�ș ��|Ϡ ��'��6��N����\��L�4���v�  �3Kp�+k�����$!.A����'� ��@�SjU����c8�D]�����æ薨�؍��A�j������,G�Ӣe�K'�J�0���bv�Z�3��E�`Rx�$���Uo:��_���˭iH'�n`�$%uKg�S�������,����>O�(H6��t���+���F@��˙��9��w���F�H����
�L�:�VQs�d�9�8��c��WhZ��n�0.�1�<5)��8O5@��:��̩����V4�=am�?-BEJ�I�����@U�q<�4'�"�J�fU��베H��7�W�푼��ڰe�-lĘ��e:�S���YMZ����4�k�V��`<�%'�U�%�u���m��[u���c�cȮ#}b�\K��GZ��*�$��������yOzv�E]�j2��=L�٘e��˨&��6G�^����|A{���:����;&�-��
�����f]a��P��1�X��� I�����*�����t���f�Բ���m�d��GKo����D��Ɋ�:��
�fN^W�b��B�#���7p�;��������"���"-J�!�J�Y��=��b����Z�'�����Ѯ�a�/�������D�+W��f��J���t�B�c��޶��S'5� ��#H��C�`�N�Gz�˭a����
,��~��Gj�%P
���Xi[�#��%2WV��;��m^v ��vJ���ȩh��t�>ď=�a+����F�^�׾��	�y�ݶ�v���Ȑ� v�%�B�I!�����x}�9-��6C��'*��Jfe(�ɒ���=TW�����*���iŉ���E>��р����Lޅ��ㆦ�R�����C�y}�z�	r�n�5g6K&;{ѴP �����/tf����Ϝ_&B-9�|3J�O+5��>d�"��R�Q]�c�?o�S�I/�F���MJ�k����Y��p�T�I�#l��u;�<��=C�(2�LJ<'�C]]��V���p|�$S"�VsF���N 긺����o m��|����oz�RU���M<�6�2�B�m��KRGW�)[�i���?�%��?\�]熺}_a�9*vǝO5��)�
:.�l�2�ʂc��U�U5w�НZ5Ƙ�d��*��37�-�����N--<�ZA>�U�V`e$�u~NGp��N4���#u�k��f��*��lD���<:-�4l��Ի� �&���d�)�5�gZz����P�B��)?0%pV1�͔�Io��5�vV�7	��e
�q�f5�J�c4ќ���M}�+��p5 �L�4&�ӆ���9��;Ó��-�>���T��;���+=	�	�c�����v�o�S���?��Y��y`n��M`�A�K�4�x�m{��9�T5��L���F���x���f�53���#�j�x���`�}���E8K|�K���q~r"e� ���:�wo���;t�&,��[��1I%���z#�t�R-8���X���PT� #_��?Dqi�>`5������'��t����~���2}{�pܭ+��
����v.�z=�պY��Q��i���y\ؿ���9e�JE#����l�����+-"���#tMp��1�v�z�V�{n�	��V'���y�b�$2G��k��'��!����|�G����Z�
J�SOTW�����O��2x�w2wL��u�}�L��	��;��w��� V���A���k#�N�?����>j�e��&GQ^��]�jV���B?����*�z4�4���/��?�m�F(�
m3��#V����i9��}4�xږ��oVU��b��s��;����Ŷ�m�Մ�~^s�VN�	���ňBor���+����@��.q��22�N�]��xy:�|������n>ݵPg'tݪo�Y����!�ԧ��x]�j:�=n~{�,Q��d25����Y]3ý����9�t{i���v��l^Nʈg���3r���D� �%����c1���|�;^��g�h�z�aUm�������y�G1X?�|{Wr��bM�С+��o��䀐#�1��ԄM(xھ��o/�i�C�����	zh����ܳ��=0gޡ�Z/��k��cP��#�1��(nB�Q	�>CR��z8[��F�����:�o���7G��æ�;��QQ+b4��˴�g��N�������aq%h(���{�R�4���u�KJ�1�HD ss�� �hfY �	��I����˵�d�׷��U\(�һ#�ܟ90�Jǥ!j�˝}�ݏMN��fW«����%�~�ǁ�)���w:�u�Z�[��,o��:�����,�X�غ���ZJ��j����V��U���Z�M튞��}7 �wa�'��4a�薁��(ؽV#O(�x+֎��=8}/�B~rIH? bxS_�D@9�4y��=�h�_���?b��C@6��=��z@a.ʗbUx)��d�����Z���k�S��������nt�Ru�Ԇ�f F��dD齄���𔸡/]��H��w�|�<`��7C�j�V�4j��4���_1V�PA���~�s`�V5Rdga:ݰ5KfL�K�����#��U��~+W��=�W*���8Ӆx8��{�}�]����D�Q�4I�f��2�|��>TkS�Q����/��g�)؛tL>m|�-�;~��Pؽ�N^�_��=���~���]����=i#Mh���F��;�K#}�ҍ�{)�U�2���1RʳWUӧ�6g�3o�?n�C�N���BkE6���I��I�?��d�L�O����A2�F]#�g��_���k�����ؓ�'�i�����%����b��ퟨ�,VV�Y%���7U���.�{V��j��D^�\V��퍛%X����c����O�3|.���'�ظ���:��nuz\�Kq��p�u]2�O��3H=JE���w�Tݟ�~w�<��ε3�@xa� ]����4���FgWߘ^6����F�$^j������A׆&����&q�f��&�����l^�D�ĵ���
��aDNT��[�X��
"�	��o4���) �����z�&y�����tk"�{{
1
���G@*�U�V_i4]�Tgi�����W��G��,�ՠ>�&�a� �F&�E.��_ˡ
�����(���.���� �?y�Z�W  My����f!�4C���=��*��3�Ъ�pFD@� had�L�6Ԕ� 3��Aw�2L��{�:{&rn�d�f�.�4�ib�ڡ�͊:F�9�k���.�56>��ꍘ��b�-�ӈ���t��(z�1)�����Q@�@~ Y�Q�x���$��+��d�L��!9�:�A�-V��)�He���"S#�R�&��,���r��.��q��ID��"��ދP�3ꪳF~�]��z����u���Φ��y��Ԓl\�n��T���tDIɡ'c�T��t#j����}Խ=7���N��U[{� ��������͊��4�,%c��4F�X�]��Mo`�X_�>T���\4������5�˩���V%���9���1�3Ҵ�܉%���jD�Iy}�r�^@�t���o.+���S[�a��u���;af� ����[x��)��b�LoY������n�L��M�� �&����"G�D�4*��H����Z��6~���"2" ����-�w<�׳�`>��)������)���X�z?�|oɈ}�1���ٹ3;���ByWW�r�1+�2˸����a�	�R��c�(썔�J���A�V�G�����%��S¹��,"]e�C�δ�cR��nӳ����
�YBE`8��t������@	>��� ��H��6I�m싍M��XFuL��Mr��nJy��Mt���>K�#*U�G�I��"�b�)�El����Fxr����Q��>8�@�V���n��_s�1\BJ�ɺ�:ȔYx<��i�6#�o���{/�0����f�!�+ ����'hiN�{�و�ܻl��jt�4�F .Y�2��Mx `�u+�Ζ�8�EggUt3MVZ�<�#o�"1.a�^��1�^� u_��*�O�hm���Ũ������l��/��T�U0�������Z�pc�MʈF��-������RJ��<7T��!��2��IQ���F�#��B��#�	�M��˕c���7�.�1��=�'1�_ݏDb!h|O�g�C����r�?�U+F���U	/.ʀ�J��PzJS�#E����UY�����X^�񍯱*��h�%�+���ԕ�����h�$:��a���ǰ��_!�@մX�qWMNU@�!<�2%C�fY�々��C+��zj�PS�~��?Bk� Xf���1�m���^Wg��u6#Q�� 3��e	���*���tv�K@�i��.�2{V���S�Io�Z��]��-��W9⇅��>�G(rƷ��ϱ�Z�������f��d[��A���g?g�q���`R��&�Ӹ�z���_�����)�m"��e����x��8�\���EF�M����}�R'AJ͋���8�uk�����{�K�K��W�P��\3%�%���Xq�w��t
��:y[��<o�~}d��w�v鎙#l�C7�;�A�Xea'�[�ƛ�ʶ$�Y�?�N�d��x>�>���BC�s�Mը1�I y:�榗J �^\������F�0�I�`|uXG��|P���US52�N|��1f,�-��%��􈻾|��d�R�?���̽Md�%%��<�r:T
�=���L�Q�����kߒv1��hN��p@4{Qi$�E��u�:�����.��<���@!%~a{x��B?j��K�cy�4b-�c$�Dc��"�x�h�x}ƓL_�"�H�I:l���;��6\�>Z���7��v��"�����]L:�t��
�%�e��;��M~�����g������������R��H�r�~��Y��:�����3TC�[��]Շ��n��.��Q类���M�Q�K��m�nB\B�.sO�v9A�!}����Ȟ�'$]��z�̱NE�AvԂ�|v��L��֥��ې�8�4�mǯ���������1��#�q���g~A,�)M��=P�~n�'P!hl���w�q�b7�:�����������]������Ng�w>iX�.�MX��(�0t0�U�C�aI�.��&J���^WW�я�������r�lw� �>�����<�;s��&���a��hw��Lmut�wr!�`��\Rf��3I��l�J�\廉��� �Kꦇ�9r�A��V!Լ�O���I4�#,\C��Ն��x������AX �%��N�w�
}��ws��q)���|]�^�(�)'?^�I[�?�zjW��+�p��~���} {Ra��,�U��,���FX�d��#�+-��i���*r�Wh[����
�����!M?[� �?�(�A���t0�Z���f�a��u�n~G��g���/ov�Gb@
^n�$Z�h���J�T��X���-�t���7|�S��}��~�� ��ו2�*�F��8I�;C#e>�!H�JP`�6�$3 <��h"��\�@��><<*�9h�S�`��M)����{(-֣����+���V�H^�]�d��n��*���t�F����zUjM֩�� �@�@�\��jYX��e��c�tiv�.�z����(��C�DF%S.�hvf�G�@���v��rՒ~~��.����d�x�Z����1֫[�汿+����,�����wa� �����x]��HY��B��CuJ�lVVuq]���%%T������\goN0�r.���87��u E���*�,�:�����A�(6H�A�E�n2EƩ����V����+�w�u��sa��7�O�zW�F�i�o���ɚ�IJ���m+M�i$~T����֭[p��z��g����>����}��8�����\�-���,7/Mp�,��@�e��_<��3�;w�g��F6qe�9���2Fn+^p����^�B�*���e�|I����`����wi�ct��%y9&]5�g����c��w���O<q�����${<~�����bE�,�Y�d���I��mT`�cL08;{��+��<���O�c�"�]K@^a\}����ŉ�B��(�XCĝO�Q�����j��c���E�ӈ�p1\M��E�R-to���E���"�>�����H��Z0���ׇ2@"���p��1� ��f.�i
tBKm9�K�\�9����dRS��]kqU# b�Ūv��IE@`!����wcs�Ip���C�Z�M��jx�@	��0��k���Ȕ���1\d�5��)Vs�=�N�d�ܹ�3x��U�q�U*1p����b���qo�8����x����OMN�������$�'jX3Ծ��Z�c~jm�ʿyB]|�-�.O���vӃ���r��]��M[�m��O��a�Y���T�=��"�TX)�vv$*�|el4�Җ����a�c�������א������㳳�;X6��6i\�������b��QZ�BNU�#���d���˟y�g[ɷ>��Z�sº� r-80�v�A����p9fA<>0�m�
��Z@�N����1�8�������f)���\�j�7U��C�+�,e�J6��v��F v�9c�ߴ�6��@ڊ~:���+ H� �������M'��a� V;w��XyǏ�W_}�eYX���U�w�|���� ���B�r[�&�j�O,��;�����+��W'N�Ș]��X4�P�����^����W�jF@QXK���8�L��ɿ�"J[�)��!Q)�����w�jm�re��t�"�?��f���%�Bq�_��b���vkX���?|��o�۳��k�.8w��
�������}�zLl�B�*˽A߫�۷���|�����.���S߾2r������<������
�.�(��|GW���x�x#�Y�$4�v�V��j.��x�Ø�5!�r$v��b}�6g0�
��aP��@��aR��҆K>,,�pI�皘%�W�n�~Ww�J����{��1Z\��JE�E�%XW��|��D1��K�!>������Ƃ�O�T�� +�3�����A�X�G2`좃ءR*�L?�s�̤p`lg�M)L2�`�A"7���넨<|0��dR��֖<(�U�E�Z2�z�^\y4��IBM2��vV�F�ě��g���0p��b'��<n�E��
%��+���"�\���J0��&R�Y�)�� �����e��Z����x��{��������U,^���u�zm���IS�R]CĒ�F�={�Z�F讂O�*)�YXTo�9I�}j�|Pź���Pw��2
�r�J�gX!�2��K</���~�w2P���G�8}n��<��J�ʟN�L�]��s ��U0/%ۡ�bLVn"SVX.d#����qtJyG�0����d��Q��qӳ�}�O��O"��J8z�;�P_?�@�O��c&�v�T$V�_a<a�b^G�Y��L�؀̶x���)3^���_b����LQK�Ō*dJuɍ#֦:���o����Ϻ�V5�!Z��Y������k����-s��Mb�1c��?bV�9�s��I��g���~��w�<����z�Ķm�^b�6�4	,n��W�rӂ�����}�������PY��C�`y(TP*�l٢s��32�#.J!T\^iR�`�����	IN�UG}�mG}h���+W�(�9�H�+QU�_8�Ȁ.oܸ��׾���k��ݧȐ9�)��2�y��b�݁~�q>�������nmm������W��7�{pdt��3�S[ʕ�ʳ»���s/��&F�X�[��C�IM\3\��$���
���t���͈���{�0J��oQ�W5=�a%2 @[p�^	,�(�ɍ�%�z���$��g����|MH\,�:	��a<#�f|��)9���B� s�5���DR--.i+�5 �$�E�ĝc*yY�M��N����=��P��2c��DR62B�3/�kdUv��L�5Ў�Y�?o�z��L���MPb��E����Q�l�_F�9\�1��&xP�FE�WB���DJE�q��8�u��]e0<O��i�3Xn��V7I��Tf��w�6�L��깳>���Aժ�eR4>=���몐�Ӿ���5��pi��b ����K����xx�8뫈�k�>��c{z�{O������Qb97J�'&''�����NOO��$�)B�@�քzW���(����^����d�?>T����SgMY�*f���J��f�M�n�n����+)���o����\�VXO"�Fd�ڰ��z�"1V�>�` �k6�6��$j^E^�v-r|�����'ο���W�}���Q���?�l=$M�lkk6� O7mڤX��###��_���~���={��j���֭�	��M`u{�&�j�O*����?�顳g�z�t�5�zynn.%T�������I���*f���!�<<�e�d,׮Q�ۏ��ZRX����m+�U1y���D��j�@���;v��k׮w��f�֥.����y�����"s�;�G�K#�>߃��@����(�-^�=m�y��K�.}���R�܂y���`%��y 7@P��L"e��%��u-w>�,6��h�X	9����mG�yTE���A�ԍ�&^,�$�����n8G\A�,�b]�9�Lݸ^\�Xg$~
��ᢗIg�Ԧ&gu��<Kq��6��ifN��������"��*0�	����iNX��C��*d����v�j(��43���&i0)��$)6�u�!�O������۶ ��2s"ܡ��8��K�c<s���P ���׃��/8�m"�H}D_
��k��c9U��}���%��0U�j��rS*�������ޮ�S�)���x�����h ���I{�T��~�7������KUj��js��0�M�|�L hq\/�v�^Qn��v���Lwo�=�t���-��i���2Q��߿~}�뗯\�47;�XQ@}����� �Ѷ��@Ŷ�����%�n����zc+�!ez8VLN#Kɍ�o )�+r�I�^ U~=;��ۊ�&��"z��wQ�_\��o귁j4�X程����(	�7�9��"_l��}����A�4�}��:e���%`����fiY���{ǹ��ʌ���j=r�m��
���ΐ9B�yy����_F>Fu��N=��C�ݻ����qej�۲4�U��ZXp�(u�<yr����ײPp��Q �R����a�1�V��P��"d����#(wP�q@�hrA<��׀�.\��CQ��}�_���NJ	A��O3�{�СCϱ:u����ۉ�-a��"���B����{0��b�n����{�^�z������笠�n����{�EqW|��I�k�"����o������R��J,q<�
\��t8�e$fJ�#qK�ذ���}$	F}�b	3&�-�K��\@@�2$�
X@ᗼVB��w�966��C	���������a��g�M�亮3��7_��Wa+� �����HsHJ"iɴ���e{BўqLx"���t�1ѿ�pG��1��VO{ƖL�-R�(B�DJ"E��;PXjߗ\_���߭�^e�C�(�."�Y�����{�{�����h�,84 �j�u<},4��c�-5X�W�1�\,,�=O��[xX;sbR�3&WB(Er~��� �49�t��>D>dM@/�fy�%�'�>p����`�D��Z���B���4�y��3�:]UkZ��YU�k����M�fjB��X�j5��t�9R��z�E�AO�2U�S���]�jiS���%r!���kU�y�K)�nU�UK��\��)_;�=!���^fT�b���ٱY��T�{��B������uXcT$W4ef#��0K���S��Y잳�'����_*nv7��T\C<���|2�QG�JЁA�V�i����<�I�È���糔�o������﷦&�0���p�TW�_n�����ktb1�|MӼOY�oGS8O[��4o�XǇ�[�$���1MR�����>h\����~�Dڮ���Z�Q^������M�@\s�ر�w��� .�<�Hx�Сo�|���uժU�����`�FIK�j)5M��D�����v|�k_����W�Z(#hba�c�,z����ɓ'5���DlP6�8� �`���(,X>l׃>V<��>Fв�!�B�hT@ٙ'�|�G�=��ɕ+W�2 �v��>|X�>}�c�X�m0�}x���ү�"|�$��h7"_�@������vddd�̛n�h;1g`Z �<��7	.i�N��=����F�b6� 27s~V���I%I �g#��p���) ��1�.�e�F�F)h��AC'�����g� ������A��Q��
�[�8B]0^'J AG�� +ԍ�'���3s�a5P��Ɋ�R;_�M6?�XZbM��*��`m��#�L%�'ء�yx��`&�D3\�`���4�(G ���"�	|�,�v���B�@Ȁiy���i-#�`�S��t�Z[�ݐ���P���lS�6)��M���6QV����ɟ�T��1�ݟQ�]��\A�:��:ֵR���w�_]�Q��n̪�kS����ܔ���:�*b����ii)v���~G���������^�>���wG�Z����Ȟ����=�A�U����$X���L��g�g*�[����<,�%~�>x�k=�f��<M�LcΪ�n�a������/?	�|���#O[������1��k��D>lrxlYm?Ĵl������F����e1-t��f�{�mf�w��O�|�}���>R�~3Zv��ᳵP02�r/��w��tM�������+�_|1x���w�1��C�;p����w���%`�˝���RZ,!�՝���7>{�ȑ^��@�Bpѹ��{�ƍ�'N@�7���A�â�!�X�L!��X<�V�2*u��O�:eNحY}Tb~Vrk	�p�(���[n�姷�v�I�gF]�	vڗ.]
R�]{�Mo�h�M���3�<�I�q��z���Ge<!o p�f�a>��"�s�9U�O�l{4�@�X����eN�9��O$M�(j1,�nԗ�p������), ��!�Ch'�BDI^����Ĵ!��Ɯ��u6��Lc)���f ��ظ���*�7�L e�3jtdL���ڰa����;@�6sj�ȼ���Oc��`D0�I�����0|W��@
b|� B� O ���I��W��6����&���,�!Y �sn�m�X0��@]�SaǈI�>�?��P��@��8-�� QX�00�D_���y�Vm�=��eʯ���2���aK�� �ւ��5V��ٲ �bFeY��eUG[���*�3f���+�T��e��8ޜ��-+���:���{�:�nS�{
ᖛv�HNFgBr���j���괍��?0�oio;(t�����~S�sY��V��LM<1>>y����J�+�+���������*���fǅ攁W1S�f��7o�AC�U��Ͽ�^~����<��d�ƃ&�.�-��=m]*a��	��Shzu^��I�y �0��& �ii����h�9!~`��~��h:�~}��6��+`��Ͽ&��)�M:����֘y��o�)4��QV�w��`��E� )fw�ޭ�9`��o* ����מx����w���z���%��%`�˟���RZ�pB)BJg__��/���ݲ�T��@�Y�fMx�w����~[�9s�~���N}�7�~�)�$g�g5V&N�A'�<�Gb}\�N_{
F�9o�Ҷm�޸����.���N顡�����X��
��Od�Ν5y}bm���� ��1�e�lņ��35=�A$��@ٸ��}�pA̓���FX���B/%���SG�@�瀽1�;��,���`�|�lGm�� P'fg)�T92[~ �Ўj@a�\���a��ħ�1T�z�����~��|�
�A�&�>om�P? ��U�� �y�f�tX��m�A�J�Рm��&�)�y?��i�F�^� 0��܆�i��f����O������r� ��p֌1"܉�"��Uss�&h�-��\^��Ⱦ�F]kQӥ��1э�-_&����رi�tJ��@@����j@����+z����BQ�,�Hυ���}q�*��w�jͷK�R:,UU U,���"d��`Z���������񸀫SV{�3ʬ�~�9=>�����܄�x�#�|S�&iQ�+_#� `1!$ZǴ\.���^=�si�-=�TBsA ��O):�Ri�}`�	���H��z����v��b�,Q�`��?���3����)q����A���i�� ��)�oj�d2	���5KEc���k����S��>Sp�`�V4	��=�QX`���U�wӦM`S6�: \��+�޿뮻�-��(�I���>��ZJ�RA�u�?���˗/��E����nS7n4�ɑ#Gj�Ν,��q���9��0���l�X�����#�� m>R��8@��n�X�Ȃ6s��w�`ǎ�K^�x��i��s�ԩ�ٳg[��ySb�Jڅ����l�����F@�'���vual�;|/BmVu�t����!�#��|d j:`#��6#�bTQ 7&qi���~����,�ѸNO���hMƬ������ƪ�>{���j��9�)�#��#l1>������+W�/�-xʘ	�o<{��6�E���	
,:}ʨEB{iV�~C����i!4ϑ��6����-� �$� �Q+D��YuG_L�@�IX:ux�/���8���a>����}�{���J@�P`>eL-�1�@E~X�,Y��1k���T5�R����5�jxd4��Uu{�rY���A�jTuI���Z�&f�TK�[uuv���q��]�sE�'�08���еQݽb���W?:��޺Q�l٣���2TA$h�_�zNTL��G3R������==����hi��??PB�~����/~^ �r�5{vl�|�F^4���Ԥش@�a?'�VN��	'����f�I�@��/X7�"�qbϤ̯�>�|G��_8�}�h]� ���>e>�⚐�p�V�&����Ǧ�>�N%4�^��6o��C����q��`i���!gF�C�vY&Y>z������]q����}���x�'^޵k���N��?��Ǔ���R�%���I��#/���Fh��~�j߾}�68E�?����n�VH5 I�;��	� ? afc���@`�� �`A��	�Ci*��������9h�����o��ۇzS�����&�S�~N���SkҰ�B���q�/�M#6�\_R��$uM�\Y�������2���1@耶utvg��s��a��X@c�jY`:��l�_�2+: F `7R3��D�)��B���[�$GJa}t(h: a	-��P(ec��͏���T������Y�׈�.�u�y�bD� �Q��%o�/�y� ������s�LUD.[ލ�^���0����Sv&�`�"�Oj,��ja��I`�Ou�,�	�W���g�j���`0���@$_ۚ���֏��[N3��� �0(��x��e��=��a.������s6���w�������
�1<gx���G���|N�~=g���ٱ=[��q�Z[�2ʁ4(�7l�)��ty`P����X�/^V-�A���V�,kW}��W�ԩ
�\ػj�V��6U��(R�d���%4��8tʞ9}f� ��;��"��@7���I�I��z�oO�;w��ŋ��Y�x;�Zh��4!K
�����dy�bqs?����a�1��~��%�V"O
��ǎGD�ʆn:#=/2���><艙
�|7ዙ�|
�ό��7���9\49M����wx�ؿ>��Ưa�g���P�/?��b{���۵�7awf�,~��W?_;�Tsmh����|`3�C"����\��<x�&ך�@��A���@�ݲeK�~�zC��Bt���+5��j���ѝ;w~S~;�l�R�n��ZJɄ���;�����C��� � }�����7n���kjr�=�T끥]7u
5��~�i��;����"�±]�r72k�E���������ݿ�ulO�5���F�[�'�X�sb�q��*�<�δ�`lT��!NƼC�u�̯?Av��7iW��`��!�4性�q�}��x�J��~+��눀3�F�yh�H�J�;}�i���yLA��,�+�3f*�<1�e,u�0]4����5��5�5� (B]�&�Ȓ$�����k���N�M�p��
� Eb1�u��h�9����s�2$�0b�Ϩ��q`tX�Q�%# ;��2��������xXa�0h�o�Դ�7�	�SX�?���k>�?����3�|�h
	3�[;v�o T�����G��gL�;T�%������j-���b�J��1�l	�&�s�*yWlN�i�,�)�TKg��toVӅN5��z��8YV]#�a�U�����k%��w�RC��tQ s�E�ڕ��6��-�����RМ6ٙ�\088����&e��S?;�+N�����/�vrj2P*}ع����c#��"ث��AS�8O��څF�jQ턯�J M�׿��g�.-P����5��J�
W~d�D^M�ת�u���-��)(M���|�����1A�oA�=��~L��,'�V��~]s��d�*���+�"/h?˷�q 21W���C�0�暍�g�?���۷��]���5��o�a̟X��gϞ����ޖ��R����ZJ.�b�!��|���g�}j�<N���,�3�h��F�S��H�X�����X���7�D�2�
�R��ӟ���G����߆ 	�f1�g��Y���̎ �xF����g����K]�[s@&�v:z��.�6��%78���m��w?Z�b�����sB}�����[6���\��i�7]d��Ϡ��!k�ߠ�;[�RCACOS1�]�#��%��I�ީ��I.���e
f�Ք�S`W�э{�B��ژn ҇ZðF�H��@���f�L�?����"p�1���4��gAgh����dGG{d�W�83R{�j��p�O�IzrR�C��Nk��9���������>�y��aL�5�E�!�~d=| i����8� R���h�h�l}��9 �0i���/_n�I�~�8��UN�2S.	�PaK��7�٨Z�2N�*�s���SiU5��8嗮���ԧUF˚�ڥZ�E53�Ps+ת�U�*s~Z.�����f��҅s�̛o��5�nU-]�"�jnbV�\::���nX+5y~���X�W�B���+h��m���gd>$���E���h��V1S2� �hn��.��QxS��k���A-��jRo�5��F5������@�\�����nH4�=�@�H��� �ë�b�g�%�5)�k��t5��h����5N�G��ߙ�{�q���G)?Y�M����� ͏�u���?5�QA�_)�]i�@�h�u�,�</���(Ⱦ`hHs`�k�#G������O����^��y�eV-��.-�������̦cǎ����>q�Dv�Ν�=�ܣaZ���Э{,Y2�Y�6#pB�!{Ow��4+�Ί�4!��%�ܓO>�Z�*���
�90	�I�*/�"�0x�T@u���'��ΩT��w�1j��n�8�2V�����-�I��{�zI�{L}B��m���>00�%iӃ�]��.lf���n�*�*���f�n�Ϧ��~P���4�fNQ�B�5
`<ťF��qM�����4�{���^��l�H��\��v�
(�V��/��Y��v��$c���b�B�K���8M�0ٸZ�~�{�R`[{�1�
����ѣ� �6u�F�+�T�,#�I~sV�HVA�P&�o�dBj�(ty���L��C��̑p-��S3�y�a�3n0�C� x���@�EK}�|Ͱ�����1���ñ@���z�	����Ȩ	�w&u��4 ��U�ah���|��5>ѯg�gUKN�k6��Ț�̄S�Y]h+���v�m_���+U�w��̨��O����j��ӝ��G�S��w���z��-�.S|R�'����<�ʗgfdtd����M7m��)���~�b#+��Oo�~���/_^i}16�p<�T���=Ag����$c<��$}rb>E������}*2�2�q߉���F-�s���1�f���H��V� ��Q^�uw`$ >mx��������d/��/�Z�P�>0M<��:?t�be,��r�zZ��b&��z�H_^��Mc���J�A�μК��>b������2Æ8�9w�1W6�B��F����_�};���
����~������qY-��2-���D�z}���M/���W_}5�w�^}�����_�uТ��J�a2�Q!�X���Jp�$a�,<ʽ�+��`y����y`�ƍ[����7���N���`E�@��h"�)����pTٲ�}ꩧ��,To�n��*(�?�Z���|~(0�6��`��ݣ===`Q�D�uS���N�~]ڵ	�����>i_ ��#��J%�9�G�`��	��{=�@_��L���Ob����@��K��T��x����A��M` u�u�q��ҦF�86��G
q��4���4W	��B{{+���6l�вX�#H)�<���0�!�'��L�0 ��w}�D�_��u@���6-�IN��	��7�WVHC�_��z��?=&����F�b�c�1�Zu�k:�-�$#"K�i(�����zN#��G��o�O���8�gf����eԪ�k�Aui���뻬�LNe
y=71��d|T��Z���n4i���P��JM��~�{i�vu�^Vӵ�����>=:�:^'�v�t�N����d�ҁZ�r]��y]���́���3�,�Ǐ���^�wϮ]�����5��E�GFGG?/}��G�/��/�&����j>��/�'������$L�R�@���wr�3����Eh�x蒢O��w�p	ȼ9��O����6�)h8�|%L��R	S5�~��$g�׏�js@;$�Xj$@�b�7�-�~߼���k�Xެ��ʧ��WW���u*��7�9O��5�)�.�_�^E&�ʘ3��fƷ�zk���7o��5Y�F�R�n��ZJHiE+>��������7oٲ%رcN�Y�ik{��̯��@[��X��`[�����,<?!�'_��'�~��M�6u�8qb�/�P�÷�T�$�'�F����
rښ��u�]Gn���[�nH� I�� BO@?$�/PÍ�
�ڪU�&{��'�Μ9�S6��^���d~���iv���w8�7Kk�=��� �h;y�VC�Ƌf4��Ig��}E��y{��1�Y�,ǀG�M�P&� ꄃ�(��׭Xl�a=e��(�Y?-�h�2"�V4'2�A�E`�	��#5���΀/�\����0"Ο�����$Vj�< x�٦C;�*�?N؇V�g��'���(Dҧ�B1�b�d
�0�Ë&��}��;~�F��&�����b�[�0hP  ��IDAT?P%�����~�?�E0�Y�v��r^��P)�#C0O0�Us.���.6*rߌ*�����\_�Ud�"�V&ЍْJ�J���K�wn��ΨcC}z��C�LWT06�������{U-US_��p�k�^�իzN�+�@Ō�D�AX���'W�tv߳aݺ��o��Ila�T�[��~S@���
��ʙ˪H5���W�����'_#�D���}�Ѵ��@�X������<��p��s�S��h*<��5)Fy��痟J�&A@B#�LM�3�|���k�I]�qA\+��0I��_#'I�ïcr���������v,b�����Y����;_�n�̡1m�Q����2�9?��� fư���
��G��"��n��桇~��M7����?�>��K�����RB��_��曏�X�"��
��E �I��⒲&<�7Ęjٓ���g� �5GDX�����/�˗���/ NV�/7�`=|�ܹK.�gGyZ�!��~WR޸ޯ?����۷oP��ر>�	������}m�=5�H�Tҝ�+������� �V��d��̫�.\�-��e<�a��ୖ��� �X�0'`� ���9�
� 4�õ�(��y�]kB�����ģVwo��p�-���� :���v�e��̉ ^g,�0�&�8WN�{`"���l�#�j�lhU,�3}c��V�@��zgT3O,s�5`�3��y��g������^�ql<͟3�!�B��9�c�Z�JS.@%��0����3�����|h�c� C�aI1��)�"��R\��'���3ʅ�ϲ���eeMʤՅK@='@)�:�Zu�a��U��y�\V��/�U5W*���������j�2aG{��ݼI��xV�HNI&�����[��m���32�/�wBM��ӝ׫bk����qZS3��/17;�z����e�8&s��㙓|�|Z� A��q�E�l<�R����c�������]��E��-���������7�VٗZ���	�n}�5F�eڿ0���O�	����3��f����9�Z��>Y@��8Z@F�X��xw�v�z&���My��j/�䷦�7��_r.ڵX[R.ߊ���'k��+W��j˖-{��?��C}��q0f|��oo߾��eM}o	X]�i	\��	�l�Ex�-;="` b)�?�֟��[a�iM ���U�����x�xxL�����DP������L:t�"����c�&��o�����lo(�Ar�Y7۩��`ӦM�����S7�I`F�����vB�$���ZD퍦/��Í7V֯_�I飼��M�=&���̏<����2>1k���{:H��1�kĴK��A#V�m�'ac���31�*����0�� ���{H�O�V�����tAC�~�i+� 5\ #��wFU6S0B=�q��Ţ����;�q�b�f{�و4��79
w�d`�ǆN�I\�z@{�WŁ/���V���`#��h_�D��#���B���QW�?[wS&�E��~��7f|�}�w�A�`�N�H+�iIp@sl��R�0�j T1��3�ʡ���4��:8���v��I5�ު:�2r5;3�&�&T!�)]��t���
�5_�2ITM@t8Y��(`1-B�tSw:+௪�G�uG1�nX���ޣf�&Մ����+��1�}	����m+�ȩ��J�8f�[]�����ma#lm���ܶK}�Vo޼���S�$�d6I�P�y��
hBk�̍��j�]�"p�%\[���=�h�b�#K��������������9���C�]sK��L�˶c�.�5�� ��7!��U��q�l�ʲ���QwuK�%��=�W+����R��檚����4��̀��Q�p�VX��j����qTm۶-C � �w�yGɳ8��㏟D,+YSޑ,�{⭥��n�d�J6����eCm���a�v��>
�<�ÂCᗪs+XV����x�������O��گ������/�����o���9�Ƃ�:#�����|a�q�Zavt���?�pN��'��i�!��H��cO�+Vce�Z $F��?L�f�UU��d5V龾+�O�:��F�F7ת���V0ګuw�:�: ����J�AG����h��yö[V='�S@I� LL��<�I+B75��
���jj��[Z��Pw7� 0p�= Xhm�jbb���ղ�e�T�SSs*�-J��,�Aǌ�Q�G�jx�	���=��H�t``а"����]���!��ժ"߇
q�ж�bD�P.E�\��óG�>���J7B�����`���|͠�6��ӂy&��}dB���@̂'������9g�c G�;���`��(����|!�3Y��'F���)��UF�2 _��J�U[{1��s��d,dnZDjB�H&�S�]8F�����h��ϤTI�zv��gg��&SY�s��.�q�b�j�{f��F1����Q�]��[���ݸԧ�GGaC���lyZ}������媷�5#�Z�UU���1WR�R��L:��j4��D�@N�:��WҎ-҇�����\-���ql�]cq��d�$s�,9��,�=	 ������3ooD��P/� � �܏=�Ƅ�H^�ۊn���F�Bh�*䙩σ��T䓥j��l�ɫ��k������s�o*n�8��o��g�^�����Ǎ�>����P���k����m��UM�]`�H�*��D>��}`�>�ܵʾF�/�x�R��+k�C ����x#�s�M!��
� Rz͚5
2ԏ~�#��ԧ>���ݻ�"��&Y�� ��7|ZW7h��n�,�����w���NPc��fL(��e���υ�t͸V^Y�B� ��'���)B�?>��cG�o�>��3�� лﾛ9|�pA��2yea�E��o�@��ײe˾�裏�x����F�FY�d�:`J'}��n�Y{
g~�N���À�vvv�TIo�o�]�|yù�{H�7_��SSQ�!�vٜ��GPT�2�8���3������"�#-�/2`&&�a2erƼ&�CS�lY��A7�أk	0�[Z��ʆ1B}KK+��g@���_QA:cWM����K��\[�7��eb+�q��&�Bᰂ>c  U��*k4Z(�>�x�A�|�c>��F�,��l�TX,��ҙS{���{2�h�=�A�#A�@��c�l�j�S ��֙�Z?M�X�,3�6������H\/ 2�?d��|��S ����%\�r�#L!� �ֶ��oK�a�jz�h,1?��8==gxL�M�?�j�;�&
�J˵9� �Ml�b㓖N�� �}ʐ��&f��dT��E�]�Z�mݪΌ���<�Cg�葑QU�hS]�VL����̫ڲ�*	h���*kf��*�|b,�ut ӕ��PJ��puI�����7��cIYj
�*!�6KIpA��Z��Y�O���dP�䮊�3(���%c�m�w��E���	=Zu�AJ�|�)X�AEB�ִ������M?O
�ɾ�L%�׺�|�!����#�XdLc�����,-�\���I�h
�7�;�UW�f�cAt�wT���7G�똦Y1����#`@�ڂ������GL>��ïmݺ�Y)ﰼ�RK��IK���MY��� ��0X��]D�������|��Z�4��3%�>�l~r�	Y@�˾}�~�{��?��?�+8|��'?�z���˽�aJ_*h^�ɳz����V��g�4�|������޽{GS�y�`&���w�I���n��A0��ݜ��|$j'D?+��J���\}�b���?$�b��>�lmm�0���Z���8G����i��0S�����Ey�d��e��ȍ���EbK�B�~�N�����\I��|:�8��=���	NExs�m@�� ���ᴍ.�)��n��N���  }&�S#4���D��وe��&�o�k�<��'�Os���B?���)�g�Ê�����Tk�S���L��A��������ɘ	x�q��`-�� �O���T�P$�nW�\� ��91&�� �@~�4!H3{`
�u�4��cD�h7��7#�O�Pٮ��?�#�g���ksz�
�ժj)d�U��t�m�
�&�Bk�U���TWOw�K�}���bAw�r��� �ˤ̬�N�J�R���Xpy����ŋ)�Zk$���-�'������a
��cr\�V�e�j$�QSKBnƔ��O&�T�w����S �	�f"���W��u����\������ ���v���ۤ��/Z���Z1�r�u����[��h}�!�O�}���>9қf��� e{��cf��}�;w�M>v��a_s�m�&M8����i��I햧�Ҝ/���|�	ʰN�Y�uv��A���jŊ��	�
�w�O}�SC��~��+k���RK~V7TZW7X���l��O�:��~��[�}��^�֗�~+��o�O���;A&�@���TD����������. VHo������GH����T���B��4� hY <)`�ROOϙ�n��5Y�.�O��ǝ L��׋����U��QN�v3������5�6l�пnݺw�}�qj&u�������^+e��Ajd\�4I�l7T��1�����Q�j@TQw>9H��������3e�| @B���M��:��IϬД?7;�)���L����:�IB�+�7��ԠX�A#��nbbҘ���t�w������=P>�`��"�G6�1@ b�+:S�j�q�0��i���Q@��U�� �i�g�`��i�B��
,��O��"�� eyx�q�pH����g�Kz|�BC���4 ��������`��:V*5�=�a�ӆ����������>�X���kP�74�=� �S2X��o�5(d[��޴���3J�si�����fu!�W+�{��m��h*P��'ՙ�A�#��������Ʌ����M�:{u�-�J㳪2's9L������8��O��&��o���@V���ӧOZ���R�ه�# �oJ4p5MB���O��z��@���x�)���Ƶ�|_���\KS�&vH�<��c���χu���,��+�3�s���c>w�٠�Ԯ��~�}�.���'�]����H���ڃ^Ӧq��ԍIr��y��r�6O�e.F ���Z�~ws}a��EQs�9s��:t�;���{A�{]��n���n��!���w���7�x��7S�?�#�� S=����J��c�qjcO�y"Z�������ҟ�ɟ���z�]'O��_�-�l��u`M ���#�U�I��<���;���֭[�i�r����e����y�������nR!�<�l������ݾ}���5k���w�YJۥK��`���J�"�h  C��&��{�M�jܦg65��x��X�����Z�<f+���j����^0�x����a���(����Q9���Ǌ���R7��n��|A�H8�@��;�a��?`|��;�>�O[�#�H~F����`�`�2�,�x��
#�ނ�02�4L�d�sf58�%�5odsd�b=Ok�Jj��f��Q�CLh�&��B�0fv>� øfw `��G�9��خ\�2��Z9�12$�D�����,����1�u�l��(���}���u� ���}��R��ZyN7mL8u.�3tUC��ʷ�H]ת��Kjj�ʰo�_�Vf�*�+�Yu���}}z�D^�Z�a�{��d��Zp�>D#�K����(2��)#}�^��;����I�7~� ?d��y���oJ�L��@s�k�@I)�@C�����2��g� j�D�,AE-�W�>?�o0g�|y`:�|mS��(C�@�����	8[@v�ip���8s�$�i��U�߻7��b;���?בD>��ɕiנ�fyA���ZZ�F����a���*��}�,��qu1��칁]�����VXb�k�.�q��o�:��R����1���A����#��S�W�[�<��!܊Pa
�0�/6\ZJ`u����t�|�da���_�������,�������~뫯��[��Ԭ�)f7�~���0�m��Хn��aÆ�������={&ԍ���3g������)T��<�͌�,ҧYY�k�*�V���T\�2�~����~��2�Z!��x�P�x B-��Q����?�NG?��B�v'��'I�@�ﵚX,��c�#X5���n��mmE�U�b����єcUxmށ�������m1���aFڌ������뙙Y�������\Z�GE	�ڐ-Dڪ����2 .����k���t��ڪ����>�N���L7���H$� �H"H��K�US  ��>�VKb���,�&O��v������u���0��^J���!4�$� @�FYh&!,5"����5q���n�����jb�}�F�2$�9�P�E ]�Y���'�ٰ��L K`{�jlؠ�'�ԩS�Բ�!��ڢ:�9�;0�.�[Q��@����|���T�V���u��tub�5b�.hå��K�=y�ܹ��=���?ם)��=�x%5�k1ߙ&ګEY0�����M�s|�ń���u�5���}0��M����A�~ے��d�a�w��^[�,}|��N�m�E�5:ɼ}�W����o�����O��X�Y��`��69�	o��5��5^�ٟ�Wj�M��>Yf���ʮm,_{ڮ��G���=�+�S���o~q�������<,׍��pk)%���qR��ɓ>����w~綾^
�s�E�:��g�q�|W��\#ݺ!5��EH�,B�s_���#�����J�A�رc�����ʟ�"@� �pl�Y{�M�i$�{�o	�)�/����D �"�����++ ��I%���2~A�!Y#�3vV��������G�>(�����Y'�h+�ؼ�E�V��PgK����S�\�Le�Q�FdOS=jF��kDf�1� �b���C��ĜG=��t*�!����ii��Fh� d���H��~W��hD&'�L&h��1M(�gf"����ۼict*nC �o�}tZ2�F�$c�泚�"�� �'P��;i�GA��f�~���3�3�&Hmx� �3m^�}c_3P�=�1�E���`�6p����yF��!�����^ Z�/ )�ї�B~�[u���0�H��Xf�[j��ߗ��Pc��0)��� ���81���M)|z��>W�jIU�5�L���{#�i�G��N�F�E�n\6�8qE��t&\1<��֧UW��o��\��8uAO�v���^ S2�������R�207�~��T��hbbb߅~S��v=x0���
�#�z,�6��~Q�h��怱{��v#�hz�y�y�4A��d�h/��^hB�:��@���KhS��cA|��&o�7����51*�t �c��Ly�&�APB�M��FkQ�W�y5�>x�4�Vq�@�����fjo�����K������1}�X���S������b�u����x���ׯ�馛^�=�YY#��>��RZ<-���<Aȕ��>�`���?������<~�x�>�/�σ54��HT����XAvR����E٤�����g���pQ`���o~s����d����́�Vh�ݜI
��B>ϭ[���={>صkW5u�� Ȣ��Y� �o�4���k�����X��,��T a�{�w��enm��H&htvvM���ÓXj��je��EZ�H�������1�HX�I(m��[�4Ѐ�c�9���X!���) ���nh�xB�EG3ӳjzjF���P.�i2��.��̘���+W�4y3n�Q 7<� Q V�p����N3���`�qd
\`A'�%��8T�i�E����&iJ������D���s�`�AlMG[M�E���[<������'MP�N���xU��0׃ D:��q�FS�k���0~�@7��ȸ���w��P������W�i5���sgg�d�Nҙ]C#h�^�����iz�1�9��'�<ٶ}d&`������@�4�`l�uU��R9)�M뵀+u��Ju��E��L�>���^�ծ�e�jxhJM��r�CU�U�mNg�e
,�������V�}}}��={��d^��6��Fa��%>��ci��4����GW�'v���:א`z�,ЈH#�����!�X�80?
�~�|M,��f(5O�4=k,��~���!_�e���������y�6�<L��b��O���ER�,Oy`�����k�?7|}@��7���-呔0O�����O���pg�u�X�,k<����=��ݻ��իW�$kN����������u��ȃ�#�>V����}�K'N�0=u5N'q"n�����:��y8Q�k+��L����=�����~��g�����Ѣ��˿���_��_o��� ��ӷО�ؘ��% -������ܡC��߈�J�ܑ#G�5n"֑ٜ*���Q���5������;�����ͷ���￿������̣m2���$���1�0�����
�Dh"�H�'
���
1�����e�66��T�H=�7q�u|O�jZ���Ӕ�t���-+���2ׅ�Bݝj��`���/s@<? � ;]]�F��s��͛\v�� �.�ܙqA���œT�H�Bh�h��B!o4h�vllԜ֣�vB���l�#�و�k��Oj����G38;F�>OXt�*��\��D؍	��Rs����D0�����	1d�Z<�.�U_X�._�l��-[L��'��6�6ǆ	ޔ6���	X��140���/N���l���&AMR��/4Հ�( �	�����Hz5��V��QUʅ����֭Vr�t:�z䕒�z� ��V���S���Td��*]�SEY�S�F8:<�׮���l.]����ɓ���}�>;5��O	���1>&���.b�mIM��D��w������|�}0bf��	��u��0�)�G+�f�u����i-�_~B�d�O_���Tl�����:�!W��_�E�'���Zf҉pz&�8�>�IL�l�b��}������8�C��>J�w@��˯;���1��<��8G|��;�:�7�:QS���Isi�V{L��Ț3���ye���_��9YO�@��n�����d7Ҷ����|���_~��-?��7��ls�֜�`�&a���F(5Lt �P�㩴�hM��o|�s��/��������~���/�ˏ���9ڳ� E��<��a�FR�����[n��Ȇ~�f͚1u�%�쫯��꥗^�Z����ܤ�M����/��smmm'���(-;v���~E6��2w��yEW'6)���p���m����Z ��d2i�8N���'�eY{y���6f\X�	�"��`?&܇�Sh�2HY�9�LG�?�WM�`�'��|�h��M&6�+�(��
�o���_�	����xTD`)p��^0o�u��)��9�7}�R�b>���_-�r
=�?M�X��(�Y�zMC�	+ڲR�'xA��{OOML����3��T�h�`�P� �[ ����7�/^�j�i��p�
��ֳ��Ɉp���Q�sقb���醌�� �!�Z�p��e Y�o;��m�#	I#rpw�e��BaӴS��\�`V�
L�6PC��R�J�aiX�U{�jikQ];��~����QU��-��Tw5P�$�3� �����ZR�4Wk�%��o�>��FR�ݱ����8�����e�x,!K�oL�6��f')iJ�o�SB�u )�o3��D���fb�R�eL�B?�X�����_W_��4�T��*�S�tx�h��1�W9�D����}�E����Vy�V����}�>N�g�I�2�iђ�,x�w�B@;�xع���GP��9�N֛k��"A��d���߯>���%h�Q�oV֖ ��Dg6o���e��6�����ҍ����u��.^��_���ۿ��C���]�J#�9��)4��%����֔$.��J�,�5٘_}衇���G=.��|���ٟ��r���'����T��� ?g-k�C�<��) �d{�Gy�駟�6�"��D�\-@��ѣG�,C~���y�����,��;v��oٲ��hc(�}����p�� ��<T�"Hײ�|@s�n^N�����".����RY|C��s������� �SIjT���2��;+��N��O�L�R�B�
�����AmJ�T!~��bS���\o�����`��'��(�@�<�/KON0�(,�~��	̋9-C���(��%m��}��� ��M�JA����$�T��z�~�snR�c�;�&�Mݰ���!Y'�"�jٸ�ZP�u�,��Ԕ�>���`k�bM
͉3�������d��`������A�dh�Ѷ��e��hMp舾�xB���� ��: O˂j�k�U	� fVEU�7Ra-l��n����s�r����v�i�^uz|R���Q+�u�]�~m=Ы���ZW?k�@g�zte�$㐝~��Ǫ��wԝy�#(;���v\�4��_�z��
���i5`��>�у>=axE`�B{,ƓR1s�8�����,2m�6R���� �F�D)D��� 5?v��~Lq �p�s��]F���'K���i�Hc���m,��������2�!���/�����Կ)�0�pSp�_ϱ�@�N��X��߯�o���v��.�>����oMs��$̀䌱��7�	k�`�e��Up����;�v���_��;�����˩�R���%pu%���í"�?��/<��K/���[oa��1Y� _,J�B��Hڲ�YtR��=����I����<�L�Zu��W�������$�I�Py�Z�@�%hό2h� ߽�=�|���Gn4`eFw�-鷛ȆD�n��Ihh��FZ�ҭ��:�gϞ���ʞ8qb___�g��w��u	�������|/�	s�:�|�~{|S�td�b~C ��Z��8�� A��H�o;�@Ҷ�6v46��\�LF�ɟ���#�Յ ����ٳ"țߌ6m[�l�*e�"���p�`�����AC�����ؔ�9����#�A��Y�G��͞�{xAˌvXut���Ȕ��4v� 2{����썧��p��~�A�HQO o�=�-��{�1.F�� ���f��0PE�/���>@?a�A�ߋ/�q������4Y��/n�l�߭@�U�xF�Ve���EP�qG��'��F����Є&�� ���/c�B�Vhgaj�K�� � &��/3%����FM�K�J>�0��:ȳ��Wm�)<�__�����L�\]�v[Fr�J��tE�xR5=S.���C�?�(W:�`Z�*�&k���?#�u����jv��i��B��y�G|�'�/���}_`������w!�? �k�����e*�;��V,�d~��8��I�����k�T"_�]������y���b.5��� ���?����{&���P��b�'�O�""�| ��q��_\9 �Є��4�����?�}�7^%��;Vښ7�gܮ�&_���k�Eq;�5��s�j|˖-�l޼�Y�~.{�R��IK��:J"�v���;;�}��_9|��!p@�`�q�Nas� ������xQ��i-�q�O�������o��o�|���Kת� +-��z������ X���� �p����36��=)��{����w�=�n�$�*��/n}��u�Ĝf#�I1왲X�N�����˟۰a���]Oh�N�:���d<"�򑑑v�%yp�U�����6g�2(�DJ9F.e�Y�u��A�s/��V�A�.M4c�`:0s#�.�0��3�|��?�9����,ʅ?�%\�50�R��oc6��q�P/l� "M`46�!���y�sl�j{{�ɏ~>4���`�D��eU.�UA&p,~!%��E���P[����\õ !�<R;d�VI�A�	_3�xT��R�[�r#� P�0��T�ew1��0����O�	|gL3�o\k}���i��a./ +Ȫz0��YR�k��@?FZ�H[�J�����;�y������;5V� ��?�J>��\�5�l`�l�ԯUʪҨ�@#�<W��S��ҹ@��Z��׬SS��j�^'�5�*u�)�&]{��E5�������կ>�k��;� (�m"N��͔���;u����p��@�@��9�L&hj6��T5XJň��6���>Z���<�5��i����̛Ԙ���u|&�h��m9�V���"��<�o*nff����7����ye�xt��!C�'���r�����Z�'5Uʮ�I �8��=����I\�xHc�*f����!�������-?������[M �1�55�����I�Qڳgωm۶�cww�ے���ZJɴ���$��������7��m�LmڴIÔ�B#��+W��`����V��F�`�G���޽��"�T��}뭷>#��o�b��.�F�O�갏�k�9 ��0�8x��YY�&S7��Jڟp�y����cǎ��6:vr��OC��1�^�q{����cW�N����ŋ���;$�^�E�L��Ν�8E����Em�g���-V͚v@���ˍ�ܚ����9 X�?�� �hLw�	�� p�gfhhP���Q������{{{�� ��S,F��#R��;�@I�1B X@>����Z�q'0hCҀG%�mM���G����?��YJӜ�i� oS:��f�ׁ
3d��Q�GDfʷ�"��p=4yx�34F$�`ic������#0a^0/-�5�@.����HPm��09�|A�b^ �&`q��M�X�8�@@�y՚�Ƥ��i>e"A+�϶���LE�uX�/�BF�U�F���+�tNƩ�j�5N�Fg�joi�:-SCR�K�e�F�)U���FJ�ȩ����?�Y�䣟U;w���Y}g�V]���[G��;.^��]�d*J��\�|R��&�����w^hM
Ʞίc&M@U��Ʈ+�����Ůѩ����'�!��F{a������9�i���5ȯ/�4t��^?�t�1pe
����6[��y^3��6{�'�K�v��X%Ƒ�ŀR��&I7��?���2�&@���o����}��#X��I�!3�ӱ��}���{^��5{6k����;v�طo߳���� �K�j)-HK��:H� dD�^%���~������N�T�&�]��j`` M�̩�=&���IP��={��d׮]sתϑ#G:��/�b����Bv�u K>Y�	���j��H� ��߿��|�k�^���1���}��у���R�[�&g��^�֤>L V�֭[�߹s�)�1��Z ߾�D�}̀"xXM�?�s��c$�v�c<5�ʭFL8�F��a~"y 3����-eYϔ�S�v���g��r�_l�6�1W�].�\ `Ш�����&���f���W�Bq���Y�5- W���l����� s�B0�=ж�{
�ּ��)2?�Z��f�M�ȿZ52uT��>C������L��yjC���u��,S3�1����=�aO�������v 5e5���E3B�4c|p=�*\k��"����? �͊+�v���Q��l��cE5��ߋ&�04�`C�� �3I�G;8�6|�!���I��?�����*B^Z�H�7[���@�TFǯR]U�J2��.�5��%}3��1��%=<6����զ����wޭ�u���ZQ�V�Ʈ\n9���n�nmѕ��^���法��Y|*23E����{5mWL���8ͳ�烶�z=����:��wy�恗�1ID�]�5?1m������Cj �ړXYl�_'��^����#�@��6I���ʌ�cD%�jLz����&���ÿ���mfO��7�.���B�BZ�x��Y�1�%�>ǔ��p��6Ⱦ_��5k֌����"G=/�-���XZW�GZ.�ʆ��	Ʀ&Ymmm�Z0������5���"�|#�����X���=�бg�yf�Z�B���|���Ç��o�
!��pX�
S��B\ �%B���C�^>p��;[�l�!)M/_�|����x�ĉ6 �!ɚ��	]Y"k-���ݻw�ݷo�Ǫ� �r�����ǿ(���̧"4*� `0��������AY��}��٘%�pB9� R��̘�etL��N�ԩ�ScMP�zq�`˔o�(��B;�c��B���e���+�o�T�
���<	>:Q���d V�#��y i L�1����Ckk�����j�:_��`�?JMT��h�L@�1�tl\)�����=Ј	Xx����3ɴ}��UQ���i�,�0�CSK
B�[�G �&7 s@� 1�p�j�,#�)� �\���l!�;�� +�lVg M9�x`l�;m��j�����'�=Ae���۾P3�T#�
2��\A͍���ɩ�������Y^��y���+ɸ��V����JW몫[@���k霖UؕW�<�@�c��ok��Rٙz=?;=�~��E=1>.����V����!}]���N�	��i�B�j���4c�K��?VRc�<PF`o�)<V�$�1N�DR��B偧&��i�	�/���ɁV���1�x8��ǁG߼��g.�~nx��z��ľ����'_s�����^���Լ�y6�IG���,c��Ƴi�ǃ%���߆5���
ǖ�+ϯ�ϵj��K]�z!j̺!�{E�����@ ���֭[__�j�r�����U���%N�@�J�)�P��p׾�V���L��|F����tx�<��]P�L���@MLͅ�i)F��ͬP�X^��5�Z�v��P��s�=��������&~X���,e+�h+�1v�������[n9�cǎ�ԍi�~���[�f����":�M�R�1��!,�D(+�U��/�ϟڵk���?��ϝ;w����Sӳ3��&��S�S���=\�z�.�< �2@�ӊ �
�m�O>�3�@�	$l7}�"�* �8�G���j�3������EX.Ut���^P���p:���Qh?�%i1��(L �����9���}`���R����7��UK�ܖE�S�-�aw�*C� *�Z&yZ��e�g��3Ɣ���C���:�"@rBSB�Jղ���r�r��F)����`�7. ��Y"|O�9�8�����>*�"6�S<�>Z6N
#���$��q��o�jB�g� ���@GZo�%���x�l4Y�pll��PY_NR0�-���"9	gjWטKyq��"�e|l\��S繁i#�Ζ�T*-}V,�h
� �К����*&ż���c�-�2t�"��7�f "�F�� ��4}��q�w6@�9�2l��ҘΥ�.	6���\ReC��c�L�Z��.K���TC���̴��U1E��	({#7�ۤ��z#������?�����a#/cZ���+�ԙ3zxd��*t��0q����g,S³�S��QS����@ۙ�e�\hXA�aMv���^�d�Ј Q��� s`�?<��/�'�`�v�(��4���_#4ʪ�QfS���։(_����3�c����Ӝ� �?4wv��6� M+��|M}ÒS4��y���|�o}���D[t�l��3I.��e/�f�d�%�߫sS0m�/f��T\���L?/����w�s8.X�h
�ZT���y�n�/���ŋV�Xq���_������q��RZJ�HK��8M*՞������uX����ٹښB1h�̪��{զu�*��p�����=\�i����A����D�� �6��엾�������k�����ַ~������B$��
�eYk2'Ѭu� (nڴiT�yc���}�������@ᕗ_�>s�\gdj�8Նc��	p�� O$�a�T[[��Ν;^ټy��F���kϥ+W>761�?NNN�F\��0��EKTQ	ML�{�ȟ.�n���ݘ.�'�M $VXS�]�����j�"!׀&׀��D�k#�k�/�T4�V`�<'S��ZP���`M���YA7Vs# ��:;:5>h��3�S����m�p���L�`��e�b����(�H9 ���PS�2��a�
�����!q^iZH�E��ۆ�4���.$�S<t�>�N�H�g�̀m	HL�X�bރ�l���C�C0�ߘ��h�
��{�7ʠ���E�	˕� ���d� 4Y3f�񚝉	a,#2����-���X,@�o�� � `���K���;p����O�E�@
��O|�9CJ�f�2E]/�\�vsa�Z�U��˿4fv*0�Ւ��95;'���l��P�i��ɜ�Uy�v���]�{��:�R��Z9;91��ϟW��cЊfU���k��
�ݠ`	�x4e%Þ��Z�P%L���5n��� Fq̎�9��B4�����7��.}G �g��b`d|�����M{MM�R�� �i����$�Om��vQ�&�;$�\y���D�Ml�M6?jjv�5�_-b1v�$�c[|so���R��>_�6lpt���6)�Cc�19�$Y���ɾvy��ݯ-[��EYN����>BZW�d�ű�˖�#]S�m̖*_��f���p��)U:u2XYo��z{��aibJ�� ��k���;�fJ�l$�X� `D1`��K`�[�jZ&��ߵk��5������VO�����p%�����[��njw�y���瞿۱cǔ���A׉����_~'�"t\=��K:Qף_��;^Y�l�niI��.�y����[��ctl�Ω����b�:;��}@ �<i�S�6;y�hO']�$
� @��d]���fS,͕�6)�5�0�K��	��_C��H�R&p�zј�Ҭ�j[B߇	}�?$\@CC��W�I^��F3�әP�����2��q���`���>vC�� PR�m�4w�
�@e�����{>��5�3�hkk���	�2"�$����$��(���1^��'Ż5ًL#�<wB�S�Sa�aF+�z�>��I�5t��4M3:��}�,弹s �	��xm�1�=>1n#�9�)4Ɲ�NtD7�o��&��� |�m��	�Y47�h�K�*�"��������c��>�3c�ߖ���z~Ng�F�Ze^kY� !�d�9P6cр?��TJ�=�U��v�?8������+V�5��cS��������0�H��9���Yz���6~��{!9!�
� ��v$ߘ��F(H{�E��צ��3Im��/�ɔ�'�p>N~�(��yK���O3P奅����J���U�?{e��%c����W-_y��Xh�����i�Wk�U~K�v-��f/4��cl�	�Jg��,��#�2�;Й+|�m�q����y��D���u��Zֈ�j)-������/I�%��Lezzs86���T��R�Pp����N��V��jCG�Z.yP����C�%UK�&VU.�! ��U��@h���:b75���I���.�r�-�?���}0|��g�}���?x����AH��F&@���2.�V��r��ٳ�w�q��Tꆌk%��ĚW_y�ߝ=snu:�0>'�jn��D$��l�v���'ׯ_uz�ڵ���z�;Ｓbhp聉����	y��4,hi) ��$��&*dx�&Fa���B	A�I��TA�=7[6�D���Gk[���fgg���R�
�0�vtt���0E�f�Q��<�!���Ǹ�����c0=+�b��7uB��FZ�offZ�$	D�JM�̎�|�%��Xn��!:��Y�Q]ͦ�Gc6��U�2Q��l� �Ն����oVc�����.O��/BI�A�5�t� Q��u%�=����mTV���]����T���I�@JV����4�`��L���hKBb���З *h@2�p�s���M!���&K����4K8B�GS>�,}�B�[j����������;�@�+E>!0o�+υ�0;u;~5�x3Ɣ�%�UY��l��v�[}��Ԯ�n��ѳ�r802�ﻀ��F�
�
%Ϡ�
3��$��֓��}A�`06��O
���kt9]�����F[洎kg�_����? ڕ1���g�Y��q����pA��DZ@0��/���r�ߤlx�w_�o�j�����w~ҋ�'��	���|6c!4kR��w1�8�ܒ�:��� N�G=�\� VXχ��j��No۶��5kּ(��I)����R��i	\}]�U��Q�y�e|4W�<�������ܥ~�j�>�imؾ�=g������J�"<�w�gd�x��`:/�pK;Ova����J�w��{ز$WdA�ʯ���7��4H��:���R�Y���N,$E� 	��"Q�@�Z(ɖ���m�1�����	k~M�DG��D���1�#Yc�fSVS\$Q�DQ�)�;H� 
{P��{�˗s���u�U�Z2��T�
�o�����=�����[��z^�s�ԩ��{�饗n��r�n��l�;��K }�<`��+0��߿���\s����B����m�?���0WO<���x���j�����%gc���5s�>{���?����1+$:th������f����Y�X�˖���ϼ���,z�������0nVFW�y״�2.XG^P=|2�ø� d6� ��"< ŸX,4�%Y�$��!nD�eE]�;�����q2�AWW�c��R)����^�F��{vt���b���b����Iu(�?����U�OcVYí����H\چg.Ƥ�Q�hFI�5j�����/r��"Jݤp�Ju[�Dl��y�p�P�>D�K�.#�� �y�s#�c�X�bkq�My�9���h���׭[g��Ċ�-��ԡ5�J ����ͺ��r�(sJ�� .�[�),�V�D$�?I��~��J�S��d�C�Y/���ۇ6��7�_�*�t�@z9��\6�t�~��_S{o�)H���B>8q�>;tVe��ʴ�WX[/|�j��K�.��K)�����y�����;^��KC�Q�iʬ{����,�=r�;%�P��ќ�f�q��+�a�ٳ׉�>�1��M��"��y�����g��M>{_��k�����Yb���u�L�<7a��c=0��ڰ�X�k�cޥ��6|ժUo�_��߯X��5�xCb�,��ep�/��C��5���VȂ�������g�}�7Ϧ���nP�	V��Ҿ�jե�|�o�����������L�ܚ]��}�z����ٳ��
Y�mdD�݌u���F5P�
����-��.ϓ�9�:-e�cR{�'���ʫ866�y|�6PI�ȸƫU�w�ɳCׯ�	��޽{u�u׽ua�-�=�ȏ�$;/��b��dK���B� �_\�V(3^�ә���~ֳ��ݏ���bo��F����g��71>�l�+����шK����b'��U�`D	��X�5�g�1���jIf�9�2\����`�&�	�,2�@Y:ݦc�J	{�d��P2^���A�Y��`vf^�$ӈ�	f��_�6��ީ�t�uqp0��92�����"��B1�w���¸)��x'V�������B5߲70�C��tv���V0`�:�	��K!�*���[��r�؅m�)�G�F��f��>���b�����'��l�H�B覩l와6����L�u1o� BL�3G�ݔ��V��`^����C��� �c(Z���eVD
��y��;w��3��U����-.��0Vn��Xqu�+}.J�n�R/d�	�Aa���]O��Vt�T`!�ί��U �j�Du.p
�f��je��~�>u�5{U��K�OOC�#����*?�S)\�H^��s�w� �RF�[\�b��S���v�f٧E d�Q.�����of��3�,b���&s|#$F�k��=��)�^�ߋdƣ�&�^�ߪI��ד:Gq����n="������G�~��**�ސ_�s�������̍�]��!ʡ`e�ɛ�A�V́p�c���ll,�y��_^z�ѱ����Z.���ep�/�`զj�֠5��/d*��:F��y��w�g�N�{ϜRy�%H����R��c/���d�|qN����W����~�K�7^}MgM J@���/Y9x��g��/�|�7��@SU�	(�7+2,0�8��3'~�����0��W�>��/�9q�DG8	y Tq,��6�+4Hk��ǀ7$cd伶{�����7�]��TZϞy��~|���P_&i����E �Qv��V����L�s[6l��t>V�p,ZG������/�����%����I$�ųiu1R]�'�Zb�+��b�cLK!qV�ǻ�-)%IxE4@b������<�<���ji3�^-ZņR��
�ş����=>�y�[�T�=+B��a�T��U�P�sa�J�Q��;l���N����.X$���� @[�ԙJ�X���9~_ؽ��,�&-,\����^aK���p�K>��q_�#��q�sw�-3���{m ���� ��9�	 Ed�Q���	-`д%0mц���u yx.�EK8���#,\q|���J�qo��B]ww��A�!)LN4�$8���O+�-�͓&
�q)��~���#��j���n(�I��f.��qr��Wd�*�ͳ0������x���m��޾������Ԍ:3Ħk+����u�(ISj���N�#��M]�\�	CЌjjXG�/���HY�"�K2�a${���0�|�����<q`�\VV�+���5��l.�E���\�'���rMi��?
�(�=�m����X�	��]K\���9�y�t��� ��V����U�z��˼ �N�a�Ll�2�8VhG�����޲�c6�y�GR�ɭ[�~ݺu���d������2��0�ݪ�2�T�X<=���#��11x,U<q2��J&Ʀ�E�J�M�L���J�����~5��\�V8��:<֝|���;��y�ө�U3��Uɂ��+��B��P�Sq5W����;�ةE.�#�p2�L�&��P	|����y\����Z��y��g����N��.}U���0Ƭ�ݏ�U�+��]w��_���s�BV�_ɣG�n��Oz����e dx�0��KV���p��X@`���	�����ǯ����^{�Ƕ��O���ܹsW�a{'���4^� ɂ�V�����x�[PYŨ7F�e:".�vQaq��Xe�`Ly�Dzh��8#�>�7\�p�,�	��r����(�Pǃ�ϒ�t-a|����n�-ɺ���cYx�	2�e 3�z�JV��(�aՇ���
�`T�5�q�ښ��t��O��1���A��bIn��k�hH�Ľ���@D����L�b\ݬ��cD�oA�]�حR=�n��n7`����%��q0PPg�/ꂾ��he6�����v@����JH �1��;����h�[��,�$�P8_�(Α>�uWEa�$���# �u_����+j p��7��=���(�jr�%��D��i����	 R��M9��~�z��_V��}����U-���������ٜJ��	�U��!?D?�:�CA@�j���f�h��%@C�Z @���bDGY&(>[Pt�����uRb�� �.�r 9.g��[|�W��&ʲ|��h(��y���y:��E���ֵ	~��/Q�+�콮�pN����e��rǑ���o6dxnW_U=U�������Ʈ]�~100�k:nһp7|��G,���wX̤���ȵ���oN��n���w[&�9��~f(�ύ���\�CՃ�]"㠒���1/YmO��j���<?���7|�����jǵx鍎�x/���[�3]����O��2&0X�q�SF�m�&����իW�7������>z��'�W����O2��/$"& B���7)A�d\������_?�.�`M��ַ�:|���>���yv0$<]5�{�Bg����Q�bQ)�Z���7|v��k�){S����ÇgΜ�O�޷�0�N�#����}>@-A��#�Ģ �K�$�$}*1d�� 2��a��׀�"A����予���n�Ũi��P�`�2�=�60ia����,�E��0L؁�������F�*�*�ԦX��@������4:�|lnwu��+:�,�T+5]��b�¢pg��l�|Kx�`� ߎ�����T�ڄ"i�]w;%q>���\W-ր1��
�k��M���f� ]wO�%�������B#1+
�d����� �p10�k�1�����@\Qo�x�` �z�3��M����$��Bʸ0�9�sF:�I���`�E�b���2L1�qy��9�����b)9��� �mP	ÆbA��?���_�z�%���s��e
8i�����*�~ٰvm�{_�=}�mw����Y�r|J;qLO�O�d���Q��Hרc�U!Ȉ'��3��r��'���f�Y�av�+d��W��鸰6e��LcC/p�����\��슛qݸ; �AE�ܯ��N�_�ɲ�G@Z4�2mn�sx�s���I�esش��yn<�jV�9�m�����sc�؉'���gŉ,�� B�����s�LD,G��8���^�a���41�VR]����[`%�c�}�?�i��Pt(�s��K���7n��U���惱e`�\>J�T�+z�j^��bӧ*�����Vb�L��������?�!���~O$yb��t�kU
���}C�Lz`��T�'�n���L�䱣�&N��_��̻Gu��A�:1�:h�� c���+ʚ���&C����!��3-q�湳oONN_���}�����3ަMn~����`��ࠚ=7BVC1�C60,��DU�$'����7�(:622�\V��?|��tY�P�v�J������p�B��0f�:��bŞY2D��_�����Uua�������臷�:u��@K	
؎������]+�3*��C���������v<�e˖�M!.����r������#������K���k�,�b��b�� b�^H����b� q.�ۭ!k�] ����υ1;ع���x���v�=�:��ݮ���-Xd�Ë/a����Y��	F�/�/����Y�/�u������$����P���HG�.2�4rrMNNq����L��	�$/�u����nM���}hc��g��=͊[�Q�]\>π-1rf�@"�{3a�䐁4��8&
 	�8��ƿE��2|�I��}�6�;v��C�_K���!~�`�����m���R�K�a�n�����n�+;��?k�%�1�F�x��D�޳Z��'���X��m���Ƒ����?���$��3�\	|�B�B1��*��j��= h7�*ԹR(�Nޭ�ުn�e�ڰq=��`||B�<sZ�����ZS�8�Uz��7[�NP�!�y�t��*"L �����M���~.q����'\�Q!0��c�O(�� �A��#1Nnq��!���}REs�"�dk��kR�����G�� L�^�e����n�w���k:Ϭ���y�.Pr��p������a��ݿ�k
��6D�Ki�N�bI������*Ǹ��l��g`�q���O��6��iӦ�i.�c/T�d�|L�S���<1�:{j����������k߫�l~�+���+V��B�Z,F�l�z�`��y�t[-��$��UW����dG�l����Z"�O1U~��)0-���3�E�X��Q�.ߙ�*\����:71������~K�O�����㩹l��\M�dZU�FFB�旓�׷B�[�j�V�����3��,�Սk/�������?u�=_>���P�N�N���Jɋ{�/C�U��*V��MLp|{Ϟ=���/�����|��eG�����9��a��Dx�K7ƪ��:���(��7uս{�>E�x�����@�������կ~}�m0$j~���݄�X$]&�s�� ,��kּ�������[֟�>F������������M��I�W�^�z{zU*ù����Ҍ���z�Υ�J��T���k@�����;��$��_�R�͡� �ߊt��Ђ��J0�a��;�)G9���L�A�H�A��=�H��//�H�
P��ݥV����
l�SFF��m����㷐�)��kg!߯�	�g�� `���K�M3�V��8�������vm C`d�-�r��	�r�l����5�ס�.�_ ��Gag���$���P(G�� ���c ~�t?��ILV`r�����"�eO��P��
�l�I_�#�JH�3��L�B�,i���h��� �s��9y���^ �$��^H�5q��~.˪T��������T��T�?X�P"�H`�E��������[.ڢ�T�קN�V���0����C��oTE�H�7����������`|���킩F6�	�r��F�k�Ћ���F��[-���Q\��EY�[3�<Z"��=�C�|
��;�P\q�_�,$��:�:��b����0�{��5�y	 ~�8��ؐ�ܿeNr�m��|���*�,E9`#�"���Q$��&�a���0��c�W��I�x����V�X�l#�\��G,�*pE/PRO�{����|��玝��U:Zc:���/�j��M��$�'��؁4�b��.8mAk[�nk��D��U�7��������=ݫ�t|���N�^x![�j��uv�}E��<�X-@�I���^<��͜8�d�]���+K�{����O��[WSzz:�15����H�˓u�4f�Ytu*�ۣ�� �f+d�&G��䫳cjtf����?����ڷ߻=K�Ս���N��.Ŋ}�p����$F���Lr�"Mh�=�P���Pp�С�O~��uo�}d�O�*'�Ej[Nފ�0���.�	22j�k�xz׮]��*qJB��Ç�=��#;��0N����,t�������s!�
�"DP ��+v]�ë��i�@�ǲ�v��������8??�itt4	�U�A^�:�y� XqG���_@�u�1.�	ַ� ��)���oq��h�����j��"���P0������C���-c���?�˥z f	��kkk��mnn�#�Ո�cl���!k�%�T���	,ti�����[v����%$��Vr4�l(�����֩�8�i��ϫ��	����.� N>�*$�qO1l!��|�$��*}b�73¸�и�Ibg6|�CF�����x�%\ � Qa��|L��@�V�X���s�(�A�dAi }
@�z��������`������$�#mv��)`)�*��&L��Z�Uw�=R _��*:�K׀7��*Jܖ���q�1�̽����J�T�B>�sy�TD�������Ls����n��}����ݻT.1^�΍����{uO#)5��~�xCF~��F�0�kH������$I�]6��.sy��!��/{m����;N�E ¹?W_H�1��߬]n��D�ǒjy��4b8�bQ����ԝD��#�^�n_�@Q��k�v��כ�F��t��Ϣ	�nzC�-��F���ifƙ�dEK�H�´�}^Dyd]�m\���\������پ}��i~��˪�\>��Wd������O?��W�س�Z�t�B��y��unvN��IM˂*�;�	 �%*W�jM�I���ڣ����i%Gv�ѸVCmm׵f�o {WUH�P��nճr���ɀ�8W����+W�aЮ���rSjndBe�����l<93�b��ZA�`[M2���d�Ų���J��l���2-�\L�Q� ���C��\\���]��k���W����8��=vY���R�������S?�
�V>@X+����D?y2lf�Ä�������~���� �P���P���e�.�F�'�t��7nذ�2���, �����_�������_��Ғ�Ć<��h��0��Y���Ȼ!qNxN[�l~r�%�>�g?�>$@������[��Q__�Z�f�7��V���NG ��,�P,�'Wa��x�]��"��!����S����S,�`BW���F�2��ų����ٍ'!^�z�ŉ�	+���M�=�a ��JUb���p���UU��<'�����jU�����N�c�wE!��
�@kes$ќd�8q]7�	��kzg+®�FV�,$��]�,��wƎUW�"�W�Fff�1�>d#�$��xc%9m�,R�QQ
S�> ����eǳ�#��Z��}5�"J*�~#��0� g�D4cIr����āY�	nZ `&�<_�5F��e�<
���K2��9Ʃ$�.�:S����y\��%����HmF��{�W}�k_׻w������ӳ�~�_%[S,MT��+���aׅ�	�*��!�̈́� LqY�E,Mh�线xh0��B�ה~e$ǽK�50S��Vu9o؈�-.Ů�����b�?�j���>Z�w�$�K�i��d�a|&b?���Iۚ��}���~��^��W���L�R�_��tc�,{%�t�R6-�a��@�5��^P(�a<X��B�$f������Moٲ�Y��">�}�9"�˅[>5��_���%�\��LvvC�RȤiݝ+eUR�hq�A9�$-jmm
��9Z��u����%�T�"h�K �O���nz��1Oײ����T�dL�4�$���P�vZ�k~P��5��b�r϶g�a�+�+��|M�";ʏ�j&^����[R���EǃB2�� y��T�-��+����3�	ZH�t����pՍ7<y��w�\���S�;wNl9�k"�G���>��u��O�W��1�&����/;^4I�i"�&�sI!����Mo�������Gpq=4�c͓v�X	\��%��+j�����{�y�[n� w��$>����_L uE��ρ��փ*�*P���q===�@�0Aq��o|�K��ܲo�G����o'ɰ�1==}7����ŋ�%<v1c�$Xp�]7Ƒv��p���;qn>,#IE���`Y�c+�P�����Pss3�qLBp�c)t�4A�T�)'�2'Fs�^�l��k����`ꮮN�|vd�7Z���g� ���F`@kzfJ�f�z�9��[S��"�v�`iu�|��a����)������ؠ~���>�O
��6W�cp��1l��_���I�$.o& \�%��
E% � Vf��p��ccc\G�I�!����g�?�.�[�<�7�,K|�l@�9v���EqU�#�z�%�_��Qg|&��o�21<E5P�1F\C�y��b��.��+��T.1S�Z.��/�\ݼ�f��<r�lN�3�O���J������ǎ���Ls�5�+kF�C����I]�àEO��E�M�uQsݽ���0���U�X�V"��*q�Í��\�@[?�o�m�et��D���Dۦ� R�5S���u�N�-��9�R��(��n�����b���#R��?
|�ϵ��N�����@I��̨����1#��<'�lz�ZY|>_6����|n���4���z�ֹ���-���q�O�2/-��W���z��w!�B����/����Nu���-z����U!�� <s攞��T��Y��|AM�Usgϱ�D�I����F�)���>�'�BA ��
s�*�b:S��'@Q��BIװq�]T��C�3~U����Z��15ْ��dYU�(ȓq6B��؈9�fj���\����l������7\~͓_�K?������b�l�{�X�-V���|��a[�5�Y ;��3F��qZ���60.������?���j�S�g��-�CZc�\�r=ݝy�l۶��0z��َ_��W�}��]bV�]�@��m����n�߿�A���Uq�1$�M�V�\1�����;��?j}�L_z�~�ϟӂs�}0�*X�T���>8'n�t}���݅��� 瘜E8G���	 �\�CF�o1<�]����p������ܼ��2d��`� ȑ]u�L�e�.r�ev3yі���0* <a{CC��� ��5o6��/j��GW���L�����2��0� ӱ'F=��R�wc�0��D�1k�����Z��8����d�&��B�8.��C��80yd$����@�0<,�b\�d�U�1 Q԰AdrPq_������6�y�	ӜWu0xb��}�����C������j����H�Hs;A��(��Zb6L쇭#ލ�Eepn���\�K�@��U5O�R)�RA��}_�Yv}������-�oa� ��5i��1��sQ���Bi�8C��@@#fX�z�Y�1W8��ClK�2Mn&C~���Z�c��24^l�+bC̖{<ޱ��[`<p������X�@��Q�gJXY<��&�����s�y�/ �ݔ���pĀ���ɹG�2`��.���_5).�sب��T��ȴ��	�Ujq^14�}�"�m`<��x���!l�C����*H����z�������5k�<E��	:�#���e���S��$+J��+�>��׵m߭j���)V٫fUU�T�=�R�N������+�B��|���
�~���|3x�?�'���U��:�J&x�F��
:Ƞ#�P`�_���.�b5d�4���kO������z/N�1rtĂ�����\��[��/~��!�)24��Z0G��KR,v�Z(��������p��}��E��˃zd�����[[ɕ�d5��'d�~�^kU�ą4!�q��K/�>����$��w�I>��㝯��:����d�	��q㲻��kW�Vܶ}�]�v߹s璉�?�L"�D�I|�����������&%�� ����k4(����������R9�窫~s�W�>�:y���o6���궇 VI�W�^���I1��qM�˜�Ǝg�0F`D
Xr�e�2�F��A2���p��js��H� w;W0�%�%4x�A{Gv����8�1:�g\��@{tt� zݺuA(��e���x"��:s�[�B&����3|�ٹY5==k�Cqj1�d�'4⨠���Xѫzz���^=hbฤ ��wwwҵ<2JȩD"L>�h{!��eK5��,
�hd�q��%�EYK ���ۥ��Y��k���u9�� 0f�l>*Ĵ���M�T�����Q���aJL��S�&��A�Xhx&x��qc�
�9I\��3 P"���1m�Z�����_�@y�R����%���D:�4������kvud�ϩ��W����I�����N�:���O0�~��3z�b !^�PC�]�6�!�B��zhA�n�6lR���k�\p5Λ�1Q[��\7
�"`D��2޵��4�����X��6nd�Y��,�����~Qy/�� �h6�7���B���S3��'�q�:5$AnVh��o�Vy&f���9�~��1�P��M�g�1隆��]64�u��ܼ��p��U���]z�+4�hU.���6m�?hNx�.�����^>-અV���z�/����x[��?�f���+�z�}B^�L�G��`J�p��˾n`���u{T����(���%�re�ڑRU"���;G��K����^E J�W��gUa.��d��i1]��_m�~�Z�{��ܺIOT�ݱqu�����ǆ�kٙ�@��C�8�W��j0��Ͼ�o�����t��W�����?|�>�����x�G��g�2:��O�&5�&�MDq�,����Α�5D��"Vixx�屷������JY��t-`��H�����[J]����GL�$�([ڱ�3��{�?���Ǽ�~���̜9sf�~����z�;!m�2	��E�kW�aVFǆ��*0�!��O$=��$vw�=�vmW��`��똙��ev~����ɕ�B>�E����]�5�C�,��uU���"F��$�!��p�������́(���Y�&��d�0��U����w9L��'��Z;u'��b)��ۺ�5
���B���jI�UKB�δʴ�x�q��˥*�P��v�f� '��%�᫖dZ%tZŽ<��IO��W�Pa0���y�&@W�&yNY�v��*T"�6u�YM:�&��2K�K`H�	?90-f�8��_�1�#̊�W�˺��a�.&aQ�H=�i`�+�� H"���Uh7���"y����
s���	@���d���'������i[�t�=���A�W��fT6J�+>&��زF��y0���L=���11b^=���Ju��r ��1՚�	�q���*?P{�0֢�:��:PU³U��q�J��k_���Ւ�1���/�#D'ⵂִ�Ŭ�>�[�RVkW�V��?T����+��;7�O�<�r�,'�;*ުجq�NO��'`�
��'Aą��c>�ޘ�H��1:b
2>\cY��踑�]�s�C����]w��z,fc=+�s܎��̇q���Eboĝ֊���l6l.���'ni
%�@r��
�2V�qҿ�0����9��>��J��n�81�.��gN|��AC2W�U���[\ke�6s������98���L�[w\�̑Ma�w?%�;5��\����m��A߱c�6l�Ugg�o���a�\���.�p%�f=:�i��(�2��U%�è��$��1����v%��L<	�}���گ���>��KUgk-�Z�&���4-x�B�X�2��RIM�'���sC���� *�ܹs���!o��dh���\�Y��ܸq���~s��[o��ꪫ>�,h�T*�|��T)%�1м�)��n`&�N����7�zCy�'ּ��<9=q$t9�^{I�i�7VK~(p�A ?����4}7�gϞ�o�ᆧ7o�|�ɜȜ<yr�w�����_�z7 IQ�{�D�c`K��i����(���
J�:�LU��r��{��}q���	\���+�s��g��?711�(Bn	qCe>��(�)fjd��#�`h�*jJY	)�J��50"'l�<f���!cYd��?0��47�c���9OW.@����� ���$ؾ�P�J����T*��L�!J���D/�**K2m\�X��^�0��RȠN�X�b�ڵp�DN+�a������� ��-��p=�'`�$����+���㮂 ��q�qWr�<'aQ$7����Kӂ>�BA��H�k���K ��1>M***�Y�<3k��m�8*�:F�<�/h<ǖ�T�Op���]]a�*�[MMNi���桁U��.O����Jl��H��
tl?���>ԍp@j��$�i����B�V�j	X��K �b|$���=b�jtl��
2�Z����R t����W�l.��K�Bϡ��jժ,.:O����U��_����;x\�N�>p��<��y�y�E+���
߅Ůp2�``C��y�t����_E���������;��{���z)f�	j���������T�2ټ��p�N���ֹ������^ObR���舂X��3�jQ,�6��I����6�W�# ����o�܉��*5J��M��gn�9�ٍ7�۲�'uى��s��۰��1GќTڴi������]btX-���iWX��Ћ�Sw|����Ԡ�؂1 �[��'y9��Γrͣ��-���c�J����<��hQM�v�.�
��j��)5|nD�������O�9���SS���f��T�w�^g鞣�_~��d8��s�Ωo~�����=:hRj�IPC�=�S X&ET1�զ���������y���/ӵzႄI��dt�L̲'�lȰ&���M7���֭[/(��^g�'1666�裏��ӟ��v�,@�g��
~I��v�ڥ֯_�8qB|׍;2d��y��o<x�}��}ر�G������k�f�NMO�%�������\7q�0�U�8��Bij'�_��\e0��
C��L�Ő��N$���kqo���c@B�������{���ty.����WH����L�I�[�Z�
Ʊ��
㻨.�A�D�*��#1nA����W"�X*��PuKq���8��U���U
+��'�x^↵�8h��]X۟`�8�Q=nX��d�قs����u˔�x�2jqAuv�y��	ToH�+�uU��\���Œ��/�'n}�> ���
�%�"���ܕb�O�����B}E�s�c�+p\=�s�� ���h�)�>��}ed��(;;�@���!�w�^V�gޓ����@�'�5O�tvf���j~��XY{-�������m�6�E�{%��6i��y�>�urܻ�7)Jm�g�4ȏ�q�:j7G�uf�p�}��`�f*��@G���!d�i� �zD��Ia�gb��P��~&m�ܳY�(q�sE)�/�n\5��EI�|��ߤ?d�]�Vw"����w@Ԣ�y��8�n��Y�pY�H�I�\��]3a�MV�+-��+�=f���ys��q�47�+W�|�K.y������au���Y.���iW=�s�\D/���*�6g�:^\��q\���{��;�ġ�0-�+��8p�>�M �s�����J͓a��+��'N�����Ԥ����bE�Z�r�y2,ߤ	���`>t�W�# Rطo��Gw��Kx	j[�mMF9��
 ���ihx�'�;::���_~9A��
�2tX2,�C�{�v�e���������pV^�Ξ=��@՟��?��]�)�pM���84Ƹ޼y3���S�Nf��6��8�����o���G���f��{tl��R����wr�]]],�����Hr[]Ŭ럀q��I��4���[Hˆ"�����
�r�q�a- A����l�I-�/��YB��x,�E.Y�����VܫV}����	���$[Z���]�tuuk\�΢�8m�(�����	Be�T7�+X�6����B{�7�!��a�W8�^ ���ڏk������A��b� ��L �Q�k�YC��0TV���1����o�.D�\��P�BH��X��x�`�$Q/���%l'���`�	� hA�	Ȳļ����6ͨ���M�,��
�ˑ�W����`P�9���hb����E$fJX|W���Q=�3����������߼#x/�[(�ɪ�U��v��w�u�F.��.����D�?�hIdo�W��� m BqVq2f}��s��pஉ26]�E�w�<#ao��6N�am,��mb	vaD�uF%z�˴8�Â�0� ���ݾq��vK ۆ"�M ��{)�����ė5��̽.M��R���p����R���N������t�"�n�V��5j�ߕ�?�l�6K�	��`�1���S����lݺ�g���ޫq:�#��.��r��W��ӂ�j||�rz�ziAM������D
P@FF��pƍ�	'n&[1}�LvF�L���f�R��bd�e�������/���}�295���3���̔��S�#T������xE�N�}uŊ��ecϞ=�o�����^�4i�G)ddİ@��a�����#�Q�*H?�dh�۴i�aR�w��ݖ�����#��F�+7�@�6��[��X2��ܹ��ڵk/4�*FFҺ��և~��7�|s&{6������n�:�]k��믿�k���x�400p�ꫯ~���)~��x�S����LOM}qbbr���� \���WĨ�X!�xp%���D �J���&1�%r��HrJ��>'�e0�E�ɼ�!Q�0sf�� 1a�_�xf����Px�����{0�j�={N#ff�m�|���l�f�H�ZU��nPk׮���lܸ�U!DAF=7�$0�2���^���H �{Y��>��U�X^�.o�{[7��)c�@m�#�
R�9E�0|f�֊0�K����D��E�ØID��/@]�ĭ�n�����z��;� \@"!`[ ��,�}ذA���K�b�]�.`� ��q�"#ov���p,�-�+�TEmb�켌�K������J�ރ�z�<��dW���g�}�,���F�!�[������4V46��$ָy�\�e�^� ~n��V����:�q{��V�D���Žy�"�@��fG3a��c��^�>s���y݈F�O����a2�;c�9�@WI���<�(o�"	p���.���b�#.��wmb��y�a#ՙ/���\�M�lf帻�W���t��s����.칀���;*����w������� ,�vs;ĕ�a���yLƑ�OXɳb�b���K�SSS�{�l�'֯_��gG��T�\~�����h1�=|��'�x�b�bQ����@_�Zm߾]oذƜ>y�$/�0����3#��;�������Ӻ����c���䤞�����V=53���,\F���ʉu������ٳ�ʣ�7l�[R�A=��o}�����|矯��[����F�R �]�P�t�ȑ�W^y���>���=��P�^����2p�,qQ0���L��U'زe˙;v]����m��1�:x��W~���������+Ļ�0��o  ���*  @�נg_q�]��X|峟��ԏ���n!��⩙�ۇ��n�E'��a%'��!��f�X�n�#!@X@7ei����C�A�Bd��1nR���c� `���0ld���s�` ���v���rb��404`U�� ���s9�,,ۮ����u�0�-���p��Ԥ�O�$�e�AH�c)G�89-����$�H���1ܬL���ʞU��'Oڝ�и���3��!��9|�k��	1�WE�qj�fG{�%N���5�T)y����g�/16p���R�m@!^J�e�$�����\�U��X�f� ��~�����r� L�
t�����
xE1�>W1��%TA� ��D(z�X�a�k	�j-�q+��*6&��������Sůp�d&�Q�b^e�Y�����+�{!�*�������+_�����X�����ٳ|(�w���j"q�٫�pK[��Dcp�$�s��RI-�Q�¹�Q����vŹ��5����{}9IƷ��Y�G�I�Yp��l���D�$�]��Y�����ƶDҒV@J�ܺ��l7���g��%�� �.}�:n��/:�k9�]E��tsmm��+��vC��f��in����`^Inݺ�ٵk��-�o�9\��r�ݔO:�j'pu��o�}�C=����/$3��� `�B9�%�q���'#np02Y��(d��Ci�8�ҋꏞQu���"�ܹ�`z����a�i��'�ܿ*ղ_�T������֧���x�K��;zӭ��%Cg�^������v�Ó|-��w(t�+�X�����������9��ȀJ?���_���:a V#)���W7�
�b�0��s�������g���`E���cǎ���#��F@u & ����4� @+���)����ȖF�b���]t������㬼����=d��515u-�/#�� �+�׫0/T����Uf�3.v7YX-��s�]E��s��1ސ�H�	\O�Hx
 �]Q�u�w:ْҙȩ �0�z[U�`~n^�+%㢗T�j��UP��ή ��Pn�[*U�n���BsB+/�X�!��J�뮆1�x�<�a엸���/1� E#m���0�l�����j0�`�F]O7&Euܘ���zbN���L�����3�D3 ��'\N��U����4?�� ,�n�h�UH�#N����5?�[�3���ųb��Q��CH�2+��c�F�Js*�V�d�ZMR`n��)�N�:4c���J��� �S�q�}SY� �X�.BT� ml�c�C��e]CR3�$���CwO�2��Qi�`uٲ�<@�.��2WW]u�3 RH���З�����s�TsV�<�{1!18�r�ۼo���1�]@%��k`���z9W52!1ejA�m��S�[�x�RƱ���1��������2�0��ֽ'{�nr����b�b�����+[�C���v��پu�}.�(T�y�VmY
�y.�.`�}�-0��6��8+�-c7�O�܎��4� t�4�Y��iӦ�h�=B�(���\>L�ă+Z��|zz�"Z��X��D���D%�w��:�� %�[U���h���;���Z�<NWR���%���-�%v���|6xa�R[&3�c�g�n�]e[���aq],�;ww	A���݃/���wwMB���]oΝ0��ꪚ~�*�g��e'�������)�WU}�0�����Y2A~@	����D�����Z��H�R5�˃��5�1/~�#>���\X�6����!���$��P�����9L�/��x*��C�:�[W|��Ŵ��ڧ��P��?���Uޏ{iX�xi9�O"++>w��g|�~g4D�%�t������v�OQC<�����f�E����6��=s��H��o_��F�u�Q��mA��~�PTk�;��O:L98e��"*�˥�#C����	@$���|�H��.�H�t�[�&Ts���Ƞ3���cI<4�߀l#�77�FA�d��/znږt 4p��r���0u����A��S�v���l�נ4Y�����6���ڤ�ts:>Jx�`v��ީ�b��H�L����ֵ�3Χ�nD�s�	i��Kr���ڜ%೺v��	���f��}W�����{0�-�U�\�7��N��=E��.��RnyXe��E�x�[�P_З�`a�zA*�����]G�cxG�����𵔏;Ȝ��/C��g��(e�������azDA9��H@.C���.��U�8-]���S���Up׀|9"���ll��[��-N����w��+��N�飕N��\�	�X#2d�?�FH��~1}\B�I5u�θhS��P	o����V)�~`�l�<5U�6@#A9��w��-h���;�/�Fz����E�ݴ���3������'ܩ�ؕ��*	Q$Le���p������������:�κ�����K�12Q��p�pYᇰ>��s��b�h6�$rG%�B3Z�()�h!�W��AU�#����4$r��� ���������U�a�[�ٖ�ָ��8�=�~Ifb�ާ�3�jYBȍi��P�ﰸ[����d��� ��	-�Ʀ�F4h��j��E��<��7���ѣ{�X~Peͼ������g�U�����3.��2t_6�޼��]�u���Cy�O(���񴅤_
 �jee�ޕ!���f��g��Ȝ��7Zcj�>Y�����N�����HC�Y�S�H:�;�BT0�����B0��O0�U��60�V��a����Хf�Ai ���O�١�������3�m�k����A� ��9�@9#���&R�����ښ~v�W��X��I�'�GsPɊd	�/�OY5���8 (���H�d�`\s�AH5�!�+B	q�b;j6���C�3���� �TP#I=�4�vwk�v�t)���t$��㾽����Ӧ2��L唰6r�jv�I|R{*<w�e-�;/�^���ҋ�뻔蛝�E>���E΀����ϩ@�OC�������~��#&3�c[U6�B�N��|��a�ԑ	��
p��C$vGV�Z�(ެ��F�e&I�AC-E=��pW��q���Z���i���X�Ys��C�٢�W����9D�l2��xS���p��SP��*���+ڳ�x;!�����S�w�B7&׳"Lѝ������)�mR��Y�ш'����$��MfdE�m2�9�F�}�&߾�ƅH?o�i������t�����"hG�]�Of=ٽ��3����4��C�
�	9�#ؔI��I�#��s�JOs�e������:�{�9��QN~�<�#����y͚��=i���:IG��N[��m<��*�ړ�{^������H��=33÷
h@��c�?�!���d���������L����6�6��uiBuFv��ڏ?���M�=�M��?M�w�&CXVZ�tZ�>�_������|�Ɓ���'iH]~i��Kz[��G�Ԗo�w�R��!�;ԟ�bC9�f`��@(���?�<���|���[w��!�ʮ5K������8��J��_�h,O8 �_��Θ} %%�l]���}p\e���e��O�"�^�Խ+>�ǀUV#m�#�;P��Zj��&l�ԭ�E��PF271��Ӎ�=*�wF[�,&f�Ԛ������/��H����Pq�y��Q�l��!����A�u�K��=M�N�.��b]��p">�k���jj8��MT��ti�c8�Sr����C���75���b���La�2�W�a�˦O[m��~�O��qD�A���'_���#6��`^GG�R�鰉�@��R*�<ߎ0{H_��H0=�ōT�,@��C6ϥB��^��X?Ť� GČr���H���-Ҿ��Yr�8��C��m�g�r���l�D�g���>�|I��Ҷlz;��E�~�;|�s�6��C&�E��\f輆��������c�2��N������o���������Ƀ�w�P?ĩ����
��,��涨ܲb/�ʄ_�B����:�{�R=*yc飻�t(�>�?�_ȟh�8r���C����vlG
<�a�At��&��E0�w;F��,ų�8F��Vٜ��<o�{���0� ��v�ό?|6##]�K��Z���>��vȜ�rw0���%��o2��,�ƻ	b4�4�W C�R���%�_!�N7�^ڇ����u봎�(r�����]�{�Z�R���#����{9q��N�t��W�-Q6��ߩ����w�*�F��R6>f[@P�~4up�zC��C"�nu���8֟��>��B�n��� �f���?���z��
����Pxlhi1�'Ϯ����*�`\�h-��Hb:�8v�*:������,�L�h�g �Pr(���Q��e��Sз���7���nٺ���B`,�
��z{:��g _�������j��P��wF�?++;'�u��=��c����gUu=O�B}T������ԦG���{�f�gV�����=�| �e�8���I�~�k�hc?h��������n/1}7�0�6I�k2��ꄦ�  �k9���mU�G3F��a0.�2�_�x5�8�f�t�xUz���ඪ���w-P{y�x��isMYA��?HV�����t�Ҩ����o$�AقU5�re\���Y���F�d��԰JT���e����z�͗���g{���3�m:vZ u�8\�/3��	�H!0�!�~y%��'��n�iͅ��Ȫ����bT�Ĝ_~�F�����<}ݢ��/�4��
�"NE[L��(��-ިIB���Q!�˾��;�����k�Ͷ�/�
s02�
�>�(خ�]�W3(�m�Yg�yう��-d�Q�Y~��}ҋ�ܻ�2x�����}fͯ�!�#��o?���q`0�55���\ɨ�ې>'5'�>�8�~�%c�w���F��d}��O�7��R�|�ہ>wk7�Y���������̒'
�����1+"'�aT��.}��0U��;���)3�J|f�/ۑ�N��w���\4��&�{��VȊ9�>�U�N��~��gq#�D�~����P�AΉ��<J���GK��ay�� ��U��W@�)���u6�YE�u#q�]���oi���h�Sx�F~�{�����B��:�G:(;X��h�!�Y,(CC7~ �-��s6��x��(��3?���J]������@�������J�����L��q��;�~F�:�BGh�`�=*+[8[J�3c))c
P����]�;�ˑ�|���v��b�}�CDV���v[�3f����sW7�I0�����Xu�^X_3��<�AN��&�l�eH/=]��"�A����F��3�>���$^#�	�Ț�U�R8}�тB#�ɧ�p9�;&a�yg�����
%I�ݺ�W�>��a����U��t��1������AIq�����L��>Bv� \��7Z��_t��`�(�*dcBLs��@�ذ�?"'Ⱶs�F�}����H��A|+���`�3��Y?�Zu^���!�ͫ��.�,.�H,�H��@#�o�'`$X��`���V��+��i}�S�z��<DF�
D&X`c__�w�'<�$;����բ�M������a��m��L�L=�����/�}�]uM}z��r#��X�@_<��XK��
��)y�Y�b�έ��%+��a�{`���ߗ�� $�x213�BL%�Fd�uu�p����*�V�\�5�9mV�.����y��(�a��6V�Dm�w�9���~?�?����Wfo	�dk֎NB�d�HlM� F;o+���>����Ry�B�79�����L�	�q ���Xg4�.&��>���W��L4��a_�����t3V�b��t��-e���� �2�ܵ�g6d�ר}h�97�i�8�(q�L��Z�����=9�e(�pP��)4�%��鶴M��0���`#����$���8X�]	E{x�A�P�������a�y���쟎��n��L�x{�!�>,`{�J녈�'r '�� &s�w�>�؊�><,�L�/������Ȏ��72�����@���*N�Ȯ���@i���B�)�w9L0���5�2G�y��5,fR�T���2��>,
C�*�y/0��c0��(ߴZ�A�HVz��95r1s�;�^?Ms�^"�H�^ĭ|ㄡ�j%ɀ5�DB4��	b�m����<-3k��ꈀ@���6F�\��o��ݍ�OH���՟r�;��	n(�f��v�`s�xI}_��<�#~ nX�&�0*��m�����
%��W��H�ܻ`��0�k�%9�	9�i`�u�'�Qz>ud �*
R�7�$� ��@���,V�-wT`��.ut��6�7Ƣ��rH �B�J:-It y��|��Ҽ�"�))!,D4�aJ,�N�Uwl0�9?��=�R���@��gK��b�\%��
�3!���������g�+����Z��)�/��t���`x>��{�u.�Dw+�����KH�<�[�eh[9{�i�o�0��݀�W��`�]DGW���:ڵ>�����72�YK@E���y��'��TzS�2~�܆����`��!/#	���Aڬ��i1[���)��bx#�؆,E4R�[�}����DrH�'#���^�G$�B��Ab��#D�ӥK�ģk�����~i�8�11�[=I5���T�'��E�E
�4��ܒ\9���U�c���w:$z�����ߖ>yR�y6���Z�8#.���́���JPKEU��Q�c�	4����:;�G�����U���b�*�z�
߿�l���:A���`�kªo�B�~V�j��� ܎ҩ.������g��J3���g�p+�.�Οu��G�5���?ɮvC�ݸ�XmR� cX;�ޚzz�;h��V��;�U��e���9�Gj���QB�4�Ņ��ޜ���/K,L�a0Ƥ @;��n��g끎��2�O[Y�n�/2i81�M������M�juT1��F�v R|�=�P��)��;�}��L�	|�i �[hnA��TR~�rC	���vtǒ��Y���I]�!��m{O_��YⳀB�U�#CwhǛ-OGR�fpܝr)�>�&��ږ��0Ґd��#.������E�2����Ϲ`��G"C�՘U���Ug��yޛ �C&�s-do�^AO\J�T��g��|�<�������g���S�5�f�D�м~����v0�p�	�J�A�1�m�*bX������1Q��IF~#��3O�u�D���5�3|���w(�*�ްdl���γaыFy�{���tR�8�װ��r��L��N⢌��%�T	ҍm��y�"(!��;�xf�vb:�����;XXǾ�)�u�P<�,q�6C�h�A�}@����a,� m��ݲ�2V��tM}���l9��H�D��@�B�ڑC�C�<����z�3��>�	�:~��x�ۉ}���w�[YD���Y�$ȲY䁾;{�9ҍ�����!�M6�����{�o;���+owc�G��,�hڝs��������Z�f�Z'|j��H:���H�n�8�dd�(?%h��sK����G_5�T����i�XB|A+E:F��S��!�S��đ)�_�L�lo��9-a]�Jsxv�c̉[Pp����.:�������kZ	v�.�6A�A���"���<���zO`��@Ȏ$�;�Q.FP���k*� ��ֲ���c�4��|@��|3�� +���eT�H��
 ����aîg�}��lfE��e ���uR~��[%�őw��<��?��4���4[Z�'�JȷL�jȏi��9��s��-h�v��E�5�P��E��l��3M�=H�0�=+:q9a(�&�����������|��;L��3����[��k�U�Ӈ)ˏf˖��|3(^�R:�i����V¨��ÈN��ݫ�S��d,>1��As���"�@v$g��"���� ���R ��l��3��`��q���lH��:+�@-���.^��v�������9��#��$a�~cKv�{B��Q�!Կ��W>���|�/C>��)@kl����)�?u�=�nx�)�-�/Sr��a���-���C�d �~��`N��VE��b��w1_{�
N�&X33\/3���X�})�����XT��#@e�2:::õހ�$��̈́ZĿ���M�/pƊƱ��y��m&�e��>�߫d��b�+^�|B+B���B���on���:Z�1I�����\�N<\%�n>���) ི���������=��lg��k�E�3ᖂb h��걄��%FR��-4�'�6!9%q阁&5kuBN�<	�Q{��#9�����5--���Ee��?�|�hu�3#�~_���U�>\XGad��PB��	ׄ��%��e=�Gq�ڰ!h�v���ڏC�T ^[}���F��ϥD�[)�V-�@n�.j�04��W���m܉�zx�� �pr�]�#6@K�*��4_�5�ei�����{��#��Q�)����kCȜB�$̇�be��˱��[�h~��s��7����(�}?��a#DH�#1n�C4峈{jRc�I�x�����P��-20�s�w�!*I�
omK�w�$�$��rΝI���<; ��5����S�:[-
	aLU��))/��(.vOs�P�<�4h}J��T.7��͸�*�
�7ú|��p�Nʧ��Ov��u��ۚ��i�_��ِ>~�K�$�u.u����!�����_!�eT�PԪ��NB�u	`���\zx;�ْ��x�Yٕ��Z?$_7��?HgOndz���JLw��=�d��"��di�7�R]s!&�޿��ER
o�]�Z�9�:�=�J��+c�Ru�ZX�x�%�،��ð�0�g�K#,���Y�k�67XOE`JX��ҳZ��խ�{�-mB@;�W��\f��[�;�6�i�?ˡ��Ld�dgw<��uz����}1���8�4pKX6IJC,��E6��I�
����*/�);�J<��H�n�����|柭�Γ.�������P�����r�����	VJ��k�Cf3�Fڷ��KxD�7CȨ�U��cג�VH�Z�c���%zMb3*�Zֲܵ��J�c���������@�N�`�l���9ڬ�'�z�1��BW7���v�t^�\Z�,��̲�ksMFr�O�
f��+q�T�Ap�I���j����}G����Rڄ�T4�_^���|^��ڞH��E�u����L�r�J��V�ۛ���Jl��`�2[=��@���ǂ6�B՟����d3��U�)N!�&=D
YT��[f�X�3�*[E� �hRK���b�t `v���/��R��b����:]���|��̭6�6�T�}<��Lr�uQK)_���w�0A�чg]�??�R��j\�
�iFp3d=��ھ*Zh ؇���X�4�O᳏�>S�,�"���~fK��I�1�$̂����5��J�c��+�їB��'�'������ԜZ߹���77�o���q�5��"�j&w��Հ���i䲆�P唂y�����s����h��e3�zK�b��嘿	�\p}�p�y�����"�B���]�8R���0�v��%|�l3{A�џ�p��Y�O�R�!a�UH��R�M��r���l�[�n�3N���w��ѓ�c��|��0��:v���c�{�E<��2������j�&��|g�5qn�M(�r�[�� �²��ϙ5��]�mpiqzn1@�wY@SW?�?����I�b��*��m���[m'J��)Y���!��ۏ�^L�>�g��}�ɵ�֭���[��V4���'mx�������1������!����Ɇ� |J��nʞ[�ol� ��Q���`8o�<�8��o���m��WYMz(�0O������?��z��m����t夳�
0qn/�l��:��wG������C�y�'��.�uA�~�ׅI�귝$`4�F\��+���jF���Vh6i;zt�v�X�VS�SGVH/��+륝�u0�~P4��i�/���f�E������@��S�Knd�sɢ�bo�&�螺���9�XX"t%l��)�R�f�g���V���jD�dy��m����o'��=tP�@z9��o�24V6vc?��O���dD������':���#g��0��'�a����g���2�gX7,��w��&����<���v�����F�땶E�H����Ѵ#@0�����-^�p�
'����&��k��H����9;;���(���%J�ű�7�r����j�	�R�fT�$��JP��1u��v}A���7�`R��=��e�6_����swz*˫�e�Q%����F�i-�C������3z�)���#���#��ҟUbvk=�3�}��KI�J�H4&V�쑃m^�.z��������.v�����FB��i#���0�9��N�rI��j�9?�I�o��aE��b�q��0'�	Z~�K�Nf�煢�c��b�Dq��o��˸���_����"/ay�?%�)�B�0Ga����	�r<����X�ns�_ݩ����]����,�ˇ�R�~T摏Ƒ�NB�S��xR�����*�Rnt��ec��V��/�hV�W�_�M]M��vq��4v�ۑ����v��.I@ԧ�����K����`��\�l���}&Bi^�/\�ʧ�����`�Rͣ.�[Df�6�}�t*=Y,��,��5��
�.� �5��ȦG-�o��&��v�}fvǱ����������������~U�DYuS�ޗ�݃��z^TD�6��ʡS���>�@�)��Xv�~��
�yn��ם�E���v��uן��_��=~�·�>��\ϊ�<�̉p2���#��/҃�t�6i=n��j ����`��m� ?~|<��2�1c�>�3{��Ӯ�Ħ�yM&�Q�����"���s�\�G<�Xƪ��
V�.0('�q�-�?�-��'� k�2�d�%Fn���8�O�s��(T+!5�5��3%j�Q�A�1�GY{5=v ���i!}d�|��B�^e��c�'�	 "g�c �k#�JG�1D"� Y6��R�3~��&�C^�o�߁�{�6�, �ԏ6c;Ŷ��ܵ�X�|����T4O8���/� b��(��)�oC�[��H�b ���1O7���U����5�t	�>Lɀ�l�6��Y�@�ßf���?%]ˈ��n�4a@؄��_Y��ˆ�$%6���v
��,`��y[�}��6���0�)���f�|2�"m$��R�q��w� 4/��`)=l�a��t������ByWu���n��_�%�U�:(D?�������] o(���Ag�r�[̆��O��<�ᘌbܾ�V ��t��5���L��f��Mї"w�?�;@ʭ[�Ξ@}�t3���;-n �me�[n(R�^bo/<+�(�IbE�p��@[ƥ/Li�O��F�x,�cgX2G��'����x}є�H�/+�^��J�z�V:�ģ���}�P;uvn�w=��ŝW����i�?M�tf�� ������4v�֙*��h�
�S���UD#��􍗎��^��6��L���	��ɏ�*U�����S�����f�Et*k3�j���B'�싿R�A�nQp���j���w���(N�i��m����F���������82Q��8���������Kh[x}}Mqn�9F�A	Aq��s�?���鵸�"#0.$P�~���ܞ�����~H�K�v5��e�P��b�(��>���^{}����sHY����$=?C
��_/�����20��}�6cT��:8�P�~�('7d+�򫠽�Ų�Z�>*��y���R4%8�?.��C�ML8kB���@��1�e��ˮ@`�!Ȗ�q�%t�����t��	YJ�³L����lT��&V�<3��~`YG�n~A٦6@:��(Vd�HV��|�Ƙ� \n*�I��u�hZ]�m����Y%E��F�y�R*�r�Y�T?�)S�@!7�/[mϖ�����E�e2�ܰ�K����;]�ս���-���;P��^�BC�Y	�7��m�|.� ����@���R@���Et�`x�DX�!
�Gg���t�� ���[����A�iC^��?�1�>z��g�(�
�[���G�I��ò���U˾VŚ���E/��1�-����%�d�`�5�H�L/@����`2�I938j����k�^ူ��vX�v荧Y|��ԉl'�0�
�#�w��m��I
�5��o�Oo�n�,D��mTJ0�8d�������eT�����e�4O���m�V����L�|ʻ�#-�3=�a��nw'�8F7E��e B�J�^
sj�
��Q��^j|���$>|��"�"꿕\�U�ᇀ�E�=��k*��f|o�=��9�Ю��R��C�0w�r�o��/É�� ��º��c��o����Y����&��i4тܻ�?ld/�B���L2��X�J�ц�^��o���>m��Ն�C��|��Τ�~�;�,�;��#�	G`�/�NQTjSӝB�r�/��XW77��Y���E��%�8�^��U�j5Lӽ��ãq�/?67�	rt�	�kv�Kf���nV� 	�=R��C>V�)�,�Y��`UT\��0fu-�F#NH:�)��^�brOA�q"��̑��xA
�m4�#�����X�]YlZo���E퐈hr4��$�B�)�!��e�
j:󺯘4je�J����ܗ���#n����f������ߛ�p�3>�ק���@�WӞ�TK��O��k>Y]P�5���a��1�V���C1�4b%�E�7��̩Ƹ�­��A��B�#y�?�����u��9\hM�}���L_��)o��J��0�������@||.
D��fI(�g���M={�A:��]���h�U����������Q0��{��Z��:B�����b�4'�A�G�~�BZ�L�{!>�#oUL���?��Ɏ��T�WJՅ
=��Y���ո�E5M޽�k�l }�`�e�������=�
����dP�0"V*4#�ڡLs�k�߉���a�
�x�KH�uP�>���e�����2�hJ�:X��,o/�ot����$����I{da^�@tgu�=�e����'गq
}-YL5qC���epy���O��\��o�ܴ3@���j�S��:��(�BL�Wy7|;�U��	Xq8�\�%��r<��L�9r�hGF����;�Z���i
gC�W2BB�΀�7ҍ�߭������X���$�������E�C2�^�ЬQ4;MCFWs�:q�����~U�Г�7`HQ����w�$xֶ��Y���s��'���flk�I���x:�.�v;v�|�D������z7��C�a���3�_��q�n��=H<a�Wn^��bb���*���1:�G��+
J�o�IƏ諍��V[o6�"tG%��/�頚`��7��Yb�g0�C"
OU����I6��a��}�j>�·;BAC�2�嶾%,g*��<�V��iFRp�_�lS@{�I��f�	���%��0v%#[v� ZU����$<�@
�_Ț!����l�)��6� ����I,	! ���;)AI��\�3���D cv���=B�5a��PNR�
Q;��jB�y�y�Ǒ���=�%�bΦ��\�h�Jqt��ц�}��1.# ��P�h�h�m���N�%/��B�7����O��d&��ӗ�]�7��o���Ӽс��)y��+�x��u��,\0��:�`��Vz#��V/��4E���(������Q���`�p��:$āڸ��Xhn����7���]��`����=D �C@��}ͺ��-%@���֝�r�`�9f"�ӹ`���M��D�[D�hW �T����).s��峖�罙�'�~��O���SC"�H�$T?�|[iFKal\L$��E�^=EqNPW.�vr�[���!sXm����:�#ci
Ԭ�RA��Gf��e^	J��fG�y&���Y��n))��>nZ��J(t���;�q�wK�+-vY�i^���ΖCBB=��_����}����I�   �㡅򲲕��5���!�~�w����E_�\������v�X�ݺ��8��f�+��2��5�O8��{/@%�^%coT�gk�窾9Cx��!Ք�l�+�+c�b��,Lx�f�^�%��Ծ|TW �R�!W^9g>�*rIsMU���W�b�F�7ѐ㫤�*
����R�yM�l���`�X(��;Z�
�__����)=zܩA���ւՖߪp��_F����.c��-y8��_�<(>q,\5�� �I{\%T�&t �Q��h2��.s���3���������GF?���Y ̣L��$Q�V��y�ݰτs�E[9�����%;����W<wQ� �t�(A'�a @���q �2-���x������t�-�6���VK�+,~u&��|P*�S���WKf\���W
�O�E���A����ff|����
{�~��>g���)ub��$�� ��>	`d�`;�VMl FZN$�u��1�e��y��<,����	�H�bX~�a�TŪ���kme��,����� ���	�3�F� �Ӝ �y�hTNX�D;)t��k��h&N%���ғa�]"[Ɔgӑ���jW�x��3�����`fv�zg�;H���9BA�9Ǽ	����I��Wv$ܧ�a�&Ցy]?�(�kq�=lY��t|�:K�z9�U���������B�.#��<��P��z.�~ң�^K �?�	%��j�pm:��[x���k=Ϟ�ig�?��s��r��Z���n�?_�^�~�[1�J�ξW�/�	���K/%��.��8���oܟ.�y:,2s��c�������PaC�睴�{�wi�{?�����P�Z��#l��1���z���S��h�]ӏt��`RLY�+�0	��PK�G~�w\���eG���gG��(�Ҏ��0E6#�ڙ���*���^�O_��_��,�0�>�O�}��ds�iT�PM����a`.�v��sk��� ��A�ޱ���7����mH�$����
����K���aƥ"�v|�5���D�P6)��4��wb�ʡ�#KM��� �M���}{7E(��z�3��7C:l(��g�'Y?�&�E�Zz�/r)�}�e��W_!=�æ�Vq�g1�e��l~��P�^GP��>� �aS?yR�^O@�:� ��?e���:�G���=X\ՏWd�[�mcө�zH~���p�[i��;2BG�nX�9��}~���m^���#���G�#E	Z$\��G��k�����L��7=pA�����rv��0��V1�����"�5�U���fB���Fx������Z|�ҹ�RZ�kR7�M�ϥ�w��=�'�M�η�v6X�zA��ҴX���C��Ʃ|��;�܋�րT�8�l���'F��Ώj�!�6�ڔ �����W�rN5Y3�TB������	n�g�c0i�����J��o�ט���m���.��]�����L�����i��AUL���X�Fˍ���O�L�KB͂|��k�F«���8T;+�-v+���F%��v�GW�_��ٸ�?v	� 3أ�vgW�h��#�G�Z�y�w߷���[p��zW��3.e*9��xA�M&3����Ė�9�G/E��w��:|�T�GQ���
$���A��.����]�sl���u0Nh[�;������
P{��Ҥ$n��@%��
tfs#'Z� `.!d2��������85)k�����*&|��E�<����&Ļ 2"gdK�2fR����`q��r���\v���{y8:�#�n���_�}N����_7y��h+oygG�F[	5����`8��NEZ_�-d�Z��I;������-��G��]��|S�yZ���R��"(@O%�	��U��ǈ�M+��l���`���cA��B�����Ŕ�@�f�_�O��l�`�ғ���ǰ��hv�E��h��uY��V�f�s���zn��I�L{(���*�&
wkZSgþ~uE��)�c�o!!]]�ǥ����K[9���� �Μ�7Lx�0��X�LW Hj��#+|�G����D'p�\��~4���+���v�k\�p��U�(�1���p�J��b=�'�qƵεs���8�֟+
7�i
w%)��"�;6@}ϕ��
�fu]���|���m)�jdj���4�|���?�����O[kϞ, ����T�D�;GF�<|���7�v�i0F(��xx@=Ee[�>t��q�?6H!��b��7�-Y�� Hm���)�v��W����S�*�H���G0��5���8����8��/��<���Q���Ð��z��ٙ��"�x{\�?�j�]VG���q,_���wě���ʟ�݊I���w��"0��~�C���1�H6���"\tU���q�3�yn�h=�Y>؆_�ͫRG�7�/�[��<��%s�_��=I_H�y�s2-�7�}��j�

�
�����,�����i�0��~��p�|��\������-��\�N5�w���P���a�[SWWW��p؋�K�����z(����2�ŝ��K��sN�����a �lc~6Z8悱�̅��/�b�W`G� G��"V�+}���n�@��q1^һ�����R�o�!m2���j���dD�L�R�u�����32�l�며�� ����:8i��vc3G膊Jy��ɡ���r��	)ֶ�z$� O->��(�V9��x[E.�(��p�<7�2RZ����.����Q��$G�Q��{j��T�CM�d2����b���`��%�،��7�������9��-�8��pc��
I )4Ρ+�qͫ�H���E��l��¶&eM��sQ�:�:W�������H�F�H��1����PЁ�
�{'�v� _Nu�21oi�����Y�y�@9����e�h�4��G�s��*�
�_@�{��M�8n��)�KlO W�˰6.�N�MG�$$�S�A�=�[Ϛ�y�5E~-��%��d����`��;}SA0;�j��J�_v���]B�ɛ%����g��ئ�K���N�c\!-�l�~��|�z�{�{��덒�HN�5t�kќ^���.u34�S�: ���&�ק�ߵ���y�wO���~UM���!��a���u����*�,g��*Y�Z�wc��4O�.t[}��=lN�|/��|�����~��z(�gz$��b����UO��<�_ֽ��{�-[�:^l�vͷM��X��귕�!���n�mb�����=���"v��?��_罯��D��y��{�^ ^�Ͼ�k��ݦ��?�b����"���~���k�������~�o���G��a�HxZdNb_8�W��qh���=#W�H�O���R�"�3�j;F$�˞p��D��$H+�)��ݗ��ю-G2E�O�*���+l��֞���|�'�P��T�<��3c�#"<���$�X"�G�C��)�������Wv�O�b����{����"mx	�ݿl8.�����(&h�쬞�P�$�������/4�u��d�!�/���L��ś�7x��3��� V M�K��\; �A�%|�~�i��I�+Q�w9��.�.+���x>�Sߦ�4���(K��}2MS���8GU!L'52���c"5F母'�����Q71���0�`��6Y�2�h5�'�o�1��qy�_�*����� �ׂ����D-�����`���*�Q
%���E�d��/S՝[��o�j5�"�s�KmD,?�,�T�;��6ݦ7��. @�C�����q�i�A��� �@e��C��c�9�ƥ��.�{f��?kZ��gۀt���|X�0O���}c�����5��oA��ɵE^���kF N j�X�1����À}�9�0������Q���K/	2�Xs�A��`��Uw��ֽ�bŊo�����?�(�X�V��J\]��ONEo$-�裏6��\��[o%�or��]�lڴ�;���{���}���O$�u�J�ݼ�[�N���������	�x#w�?��咼��K>��'O�����o/���~�������ɟƞDP)���%���Kx�1��{�=��K/��}A��=�J`�+���H$|aӆ��m嚭��������?#�!������>_9r��׽:�EK�-���<���E�B�>��Z0�����KLCc���&R�X�C�̨�"���ϟt��TmR �`���4��`8��X}�W݅�q��:���"F�� (�ǅ<' [�$�)��P�} �E��d<�<��4��'\����Y�ފkZǬ����-������/���U*m%�Yi�;<"�C���\��`{� cT*%�hH�A=�p2.t)�QW0*��EuE^��t��@a�*c�F����E*�h_Ě�eKe����f�80c`��E3��/�\T�_
�Q�/�+�bP��	��Բ��T[�三��(�n��2Yw,�Ę������;S�����1g����7���֡�¢����ttd4������v~.p;��)L���X�ʷ��c��h�BI�t��Z�����tYU�i�Avn����9c;��xa�j�=fFw@��B��[�r��ǔE� ŰZ�,��OG���p��{����3�?չ0�������eY ���.���;���3ߙ���hx[�ޟ����Gn�q�ں��]B��n��z��۶0y�";i��-�I�[֟�D���u���1�y �0�lذ"\o͛7���-`�*�[i��+��{v�����{v�ލ�����n����ח��]"�c�$�l`.�c �8\iʝŮb�s���n������5_{���׮];��ȿi��.X]~R�;z��C����_�u�k���y߾}�y@u$]�d^��@��Q��O��o�݁�BL�9���g��x�ͷ�O�8+L��F�_�� �0Z�����{�gn�����+�^{�X�Ʀ)�V�u^700����o�@1V��6bhd8����}��qG1�f�<,�`7:�� S0.�n�f�̛7�]�xN\��{�\__�Eϐ%�Q����0α8�Wmj��p,� �NË�����WA�7C�.���x� �ύx!��3Ʊ'$�����E9觉�ಂ\X�=�zh\ KŊ�?l�%"ãrb�P����SL]�,0v���W����r�A;�T7@�cla���E���㥹d��*a�0�.dQ�z}* E	�e���-���C{%��qp%�Z�߈�嶒�)���P�R���u�
��s�����߈��
�,�ڪK�\h��(]�>��w*��R�#���N�27Q�p#`φ��1�ڧ�=� �G܄�1J^6*�x�w�/=��d͚5���H��:u*���P���� ��NY���Os�����2<����8#�� ��eTC|na��Ƿ��&ә~�4~�`9ǎ�X��X:�R#mJ��T��-3�L��\=c�.�`B�/������7Sߏa�fE�~������u�R�3>����a�2��f�db�$�d�cn���OL�n���7�����0o��˖-;w��W��~�~��f��Z�r,-pu�Fp+�}�����s�=�'1�3�X ���v��V�裏�[��X6�)��HԒ���$��S��7���ڵkh�޽�|�s���x��g��S�!���ɓ�O���{�7�������OŃ�?L�X|`lj�dtt�+�І�m�ܝwމ�صw?��OR���������Kr�����c�T��/�^������ݾ�͛7"E@S�/���|߇}��G�/��x`%1F04�x� �b%F��D���K��,���� +u�7��A�ǫ�뒛��Ã͹�4��`����OqW�?\�p���zLl���ɉǧK�.6��4�w|����	jux^���8�t� �J���=��I6D�c��i{B:uC��Z̿���`��s[iS¥�Xn��g���w��� ^�M10B�-2;��R��Y����4Z�����*�. .>c,
��`� Na��O��d9�|=� \� ��b��ٽ=�}����K�,�(��S�$o��Y�߂���)2����c#�0��9�c)*թ��M�+�%M슽�ɉ)�B��ڷ���Gl�i܂$��+I����abJ���`�-?Ϋ��8����=���Gv�]w�l:!wb��h�'�J8���]����i�ϻ���1-�(a"��ƼY�gZ�N�s��������{Ɯe��>]M<aF�m
����d����B���ȲC��iǏs���#�)��ب�\�w�w������\2C;_��4%�,h��ۍ�������s���:�ո���O��Խ��ux������K7n�s������nP�J�|ZJ\]��OrK=������߮<}���1�MNTKG��AP�@�����.\O��k�.���q5�I@�BWy���7�����o�9���?���O_�n�a;	t?�[��_��7����I~Ϟ=��������n9s���`�7q{��{U]���Aw#�����r~bO�;�<�䓉&��%0�p�z+���"�kwuu(W�o.X��o|�o~�_ܷz��O���r�C�v����ae��U�*06%��Rq��aw��S4F�ƻ�,J2`.��$�kIU��B�PQX�S�N��u��ǚ�� ����FkM�
]UX#�#^����ӼJ�8�Ÿ���ЁE��x^ 
<�&�M`��h?#�D������La�sF=���(�%�͝;7��Z�E�\	��Y%i4��z-5FI�g�@�N�e\�(��ϒbs'�Ɩe�bܐ���5a�*����bQ���X8L����V�\)���ä礫V�J�R	�6���d��{
�:k!w 0UQ�n�~!�9Ւh�À����8%�ED�F��`�Bp���}�<Vt�dY������J:2rU0_`�&�ӱ�	������+l6�@����z[����-[���Đ�;�&X+�1���n�X��8�혰._y01�a�% �uC��Bg�1ם��6ng��<�h�)4U���E�捦�_te����L��P
,f7bM�/)��� �ܚ�-�-�5m9M���SF�´��W�F�1� [��9WB�ӹL�����7�Y�̊!�7W#�6C��=���\P�%���B:T6{��Y������\zk׮�����m����j�˹���V�V��`�w�󝯼��[�@��	����iXPj��������Z�N��\�8$��j(�!�)��
"=�I?�[Fڈ1��o����^{��۷o����UW]�wk֬������|0�i�&XavŶ�_r�m�Rx���z��Z_߇��n�����ݻhIc��t��ɿ� ���t,Y�db�����\s���g>�.]����?p�W�m'��H����	���ԃ���bRz����>�ʝwn;��7���VF|�7�vzp�?yöl�o�
`ȶ��/���L��FH��PR_�c9N�����CC�$*}�9��r`̈́5^"r��n��`F[������$t��2�`o��=�`�C�}C���	s1D� x�Z����L>B���0�y=�0��d�, �Q���L�"I�<����@Q��F�U�$ijC]� ��mqw��ئ���������P&,�2E+!�"#�� MhK�7��I1V��,sV�ك�e�[�;T"��a���X�)�'ꖨ3��5q?��G�;����r��a� U��"���:���U�>��f�xpU�ڡll4����s�ߙ�L\ i!���mԸ�4 �bt!�H��A�J��B��R2U�
qh���Y����o�|-�.�#����E��Ow��1yfƚ)؋I��de�F&.,Q`�Xz�%���/�$�رT)4&�-�b��e+0�{�'��%غ��+�qg���ɂ�F� �gH����͔.Ŗ�R 0S,V<�*@�l;�v�T;g�v�k�뜭�i�4;� N|��ug����lsm��4��a�b�䟝u�'�������l@�c�����p�3�瘓~�����^��\�jĭ�*,-pu?���h�sϽ�Ӄ���*�s@��3���dR�$"5����{>J@I���-��N�>�ju��P��J t[;�	�"���<�*�F	;��KmZ/�N�8�����7�۳����u��������F�/_2��7�V�k~�m�xu��o�wuͮ_HΝ��x��ҥ�JP/�%����/��S�����h?~|����*?!o<u��J�Y�Ӽ��4R�<,�:���BQ,���`�y���v�*�0�6��Z�J\�~���:����[n��}0C��̗o/o����J�H��S�Ǯ�z�<�裯�t�=#�����3��x㍫>��ၣ��;?Ծh��t�ʕ���9��Y���,��So�9��k�V�E��ldA�� �J"��k5��]N�ƅ(�Yhk/%�	\�����%J&bH`�YPTÒ.xM�c x���U:�q	\��a�'Nd�"�V
������g��i�xxD�{`X���*E:�671Vu�'�stzCxK��5K"�1^<�v�ϝu��ABᒷ�{<8�흝��c!a-ƍ��i��YL�H
��H��1m(m ��TLT�o��N�Z"�[��01������e��m"ݞ�?.ɼLr,��m�i���8+|������)��1�LS "ε�u&�N'�h߾����˷M�V�+���B���}㾝gut#ӝ����{�J�9zL����}�%�0�=��(�1,�>��j�̓��&�_KŲ\�,ʗ��������$Ďu�6���F���=i��xh��`52 ��ڡ�����B���B�M"���9Q|�{�52|��y���׿��䮻���ӝ�p�}������q�²�=� ���i��(�e�#9w��0�k�,Q\ ���������F�8�Z�@��J%� ��b�(�l�7d����F)�*�(Fn;s_<�g�qlҁ�V��9�� ��-����U����APm��{#ۄ��:�8���أ�2�O7��� �&F2�|h��wB�6��]�b�"�č�g�)���{���I��t��f���&��8f�� ��|�x���sr�������^��5k�����~��7	/h�V�M���B
uoh�|�g�|ㇻ�����+�R���,��V��hY牉��獻	��A�!Sp'7?Q�E��ZCvǐ!�IBM���I�&Ђ?����[���?}��J�������]*WhTGF.L�_�a⥗~6��V�����(��;,��$�𳩌��U ��AU̓��Hx�\H&
F�y�<�QOEi\w0�, �<'bu�17�w߾���~�ɾ}���z��8N�}V��O�$��q�[E�Z}��;���-�����۷��5��t���������vX�`����X��)a1��#I��Nmf���IXw@1԰J�`�O`�����s0H��۔�7Mҽ*�K]X0i�5�e5����(� A����Ǫ=	lLQ��·��FKȕ#;���i��tx�1 SS�R����Jԙ3���
�.^� l�6�S^�T���㼦�p["�j�d�kх/)��QCf'�[�Ǘ�F���h�F��.Qtw������a���L�E�u�*Z!1A�IGٷC�0x��]H�.����e˥��>��R@�r ���1T� w�E3RU��3�0k�y�a����]A9&��0���b|���%�~q���@K�]�-�Pڔ�&ӧ�(�ߤ5������LGGF Kd�{}�Ġ����?}��\���nE^�Ŀ�~�v��aD���モ�����(��x�B��&����Z4��>����vN0��$��ٱ}��;�
��o`T���'�Y�ܵ��r/U,d�D��y�e�2ps>3�٦0L���-�Rh�aQ��`b��d�4�μKܥ�+��3�<�j�e��銏��~\}r�e�xY��o��v��97���"28�!�@g�+S�{�s�lذa���럙={�K�%`�*WHi��+�����AQ�;＿���v}���ޛ���.�]��.�f�5�
���RL��Ն������A9�0��5]Լ}��`7���_2k"U�"�BZU����(A� 0،Lө�w�y'����`��q�4��U4υ����a oN���Km)�S��F� ]BAU4�qMM�*	pC���?w;d_Ϝ9�����sy�WS`r{�ߒx���+�n���y��׶l�rh͚5ÿf�����3��{����}����JK�.�@�##�w1��t߉*RyÇ%�!���s'D~]D2�{�Ī�(�%9�h���%.U��Xﺐ��E�a!�J�ۂ�.>Su:1��*���< ��0��!�2��i�<�h,M�1>1�����B!J{wuw�g�� �-�+��&<?�%����h�4���km�̟˵��@�PE0aB`��Q�k��fZI8~)��s1~����l����˧����tݤ�a���7�F���!Z���U�1s8W��Reڨ�}�$�K�-���B (��<M-�,c V���i)���q���:��� ��%��M8�kP���>&O�A��)IT�6�F�+��>�`r�=��E�:?��
��2���Q���w,�0�(���5�9Ɗ�r�8��"`"Ð7��g��i�����_��q$NE)x��3lD���̒�ȀN�+f�b|Vj<�0��ЌqK�͛��cEI-�*8S��@4�'��M,����ུ����K�������zX���5�l����u�Ȼ�ub2䇓>�"G|o�=���tΕ��?��bŊ�=��?�?�����h�J��[����+z��������m����Ua^,8�� LP�Ɏ��	b�� xax��CF�v���Q��@4*�B&隲�SFi(�p�����ĝ*)EC*�`���n��Y�\v�q�0�N��\t�P§^e������� �yñvq�biJ� �$!��.���E����o��իWZ�z͋�ݾ��͛7�X�v���g��������Y��x�s�-*-[�,�rN�)�fz LW����)�M���4����<��x. QG�o4����}��?�^,��$�G(a"c�0S��.mM?~��C F����d�3��@x�:@�@���70��.�-���u0�3�4a�Dݬ*;��>���C�K�����U�sa�W�l�A e���P���w,ʚsW�;�IiS�!�3N��{\��Q7�r>%�Ѧ��?0`�@�Nd�����%�龜�D0�w}�d�0v��Jg�s4��	?��]$�}Q�1Q��g�K�N��s9����^���F�����Q(�T�Ե�Q�E�cs���Ӎg���᫢s���Hr��K�X\ >|X�5��j5�a0dv��0 K��������q/4%#j��ߺ`��ilR���`�j�{-ndq�[�}2�c�A��L[6�gZ��}�Z����L�n|6��2Q9�'c�u&���˞���4s��&3���	d���!�ogX��K]�3�����<�q������}Ɂ�j�2�Q̈�%(��Ǘ�6a�%���=�׻�6m��y�^����U�\I��.��y�ڽ�p�3�<�?���?���q��y�Ⅱ���=2�������;����w�kW0�\��8*�\Lh��&x��fr�x[T���`�'S�(.�ᯀ�r,L�H�*Ɗ��,z��O�i��$8T����/�!���N�����UA$F\�ƨ������<�����-�A�X��T0je��Çܾ���Y �,�6��y����VZ�m��R������&��uh�[����Q�Svm┭Q�_�,����� V��	�n����� @0r���Hj�1&��F\�]�����l���LAf���3�j��??�XT��Yp����)�`dH�g�-M����s���(��dvC�A�������g
Z��#��)��|^��n���n5����o���{������%9�\�/����hk _�fA9R���ڷϪh�0T6%g�LN�:%c.^�s�!8����]�i��h���.7Yd�A�՘��3c	�Z�ȶ)�n����)MJ�z�F����*���v;w�eE��%����͇�G�9׾ʰ�3�y@岮`�\��yӤ��[�Z�ތBu�.�_��e
��(80M8��
e$-8c��؍߳.�:�.��h�y~�3?�Hib�E]_�{IP�w�<^ƅ:̸q��=gZ��,b����P�Ц�7S�;�0�P����Jf�Y�l�w��<?��H7<�]��o.ڕ.�30X��v�wտ{5?G��X���Y�`�s��?��Su��*WPi��˻T���瞻׮]7�T��z�QY����ui(�ړ0�%'Q?A�m۶���7�<ϋ�����?���^�4q7�,TQZ��,R�m���#oJ'D�z�tS���� 0���^kц01��N��b��:��%��Nŀe���x^?���YHK�~�J���A�z��׮[�Ӎ7��c���n��֑�o�����ý�����<p��'���jɒ%%�  X��F�hw0�N�E�F��Q��!*���D���
������ɠ�:���v��� �=>�fut����/\8A
7)�����.��V1X�����RҠQL$��xV0Xd �D��?�P]]"�.�����0 8�@� 2a� :�C�w� .q/�F�	�Q�A�g���7�p����*!��0Q���� @�(�;���ˆs Pg��J{���?e9��%h�2�5��US@�F����&
ER�{
��X�J�<ܛ̖?q�d�c��d�Ж�Sf�9��p�娒���*O�K�J�ǀx�+�$קB#�@8'P]PW���U�T�*�*_��Wӯ~������b�A�����<;�#�_�HJ�f��)�x�9��g��Q�9,@��?-se��&AB�<&��8�4�R `F��uFJ�L�8W�p���z`�a��5��	<�s ���5,H�l�m�3��S� �Y��h ֥ ̴��<�g���8���x���g�����g�_�Y3�Z��L��9�6R��n�d���Z9}���=nG�<�qx��͛��ڵk_X�t����=�Zʀ�r�����_�{�x����o~����%RLN�aq	ٱ��^Pyn�bĄ�n޼��#�<���;���n��k�������z�ՇkP9��}V:22N�L�nC��i���4��Ju7Mt0�` J�������r�s�L։���X��$$,�!5$ Ş��a�ք��2ޠ+�0��3{������y�=�������u��B��_� X}������7��S�N]��
,���Mո�U�F�,��(1��Qbw�5���[��u2���|Aѽm����\��䆚=�׍'�GOӧ�~$.
�+��HČq�`��t޼B�bqF��vTR<�d9w�5	��>`K<8Kgw�I��L��𐛝a�ٳ{���� �>���������N��;��!�������M9F�2s�]��Nd��j�+ik��*C���0��=O���4d���a�W�;���N��W�QE�An� ��k���1G ����i̢��:�z��qEm��+i�6�0fm��Oxo0	��k7��&�AlTxכ�^AcHR� ��� �Ѣ�����*�tD�p��s�U��R[�@�ࡦ �m��ƣ����'��j�u�V�-����*f��:;�]��vvuÑ*����Η�/��� �3�B�p��@C�2W����\��c:�A���i�Z���L=��kY7P���]���2^��\]�شq�����>�u��bܨmO�N�~�u�����%�S|�<��_�m�����M֜����{�i�j~�#+�ԍR]eH���~��D]����uL�c����'�`WW�^�+�����q�*�r���K#�.|��w�|��?��;�-��v�]��Y�F^�)v�zCM�rR���'���o��֝w޹{����j;w�|�O~�O>�䬿�����J�{#o�TR��~�gI]T���46i�3�0v�!�9�N#�<�.lT*y�J*���C<lP���v��Ji����Iu��J"%5ʨUõ:;�&�;��WJ�����{�'�r���?��s�����睺6�������'N��ў��9|�F�HX�҄9v��4 Ȱ�s�? *��y]˒H;k<�,vp���M��&���.D8ׂq���T,��"��Äs�O
��� >]�$_�:��:��RA,N 7�:(F;��D0��C���9�~�_���%��9Μ=-u�� =A��$ʊ~�ϚՑx@ n_��k����"�
ǒ��=�rʝon$h�Z�$w��t�a�[7������o0T*4"1� Yh}��������fk�"���z�;���MQ�\�֊`�1K p
l���}]���wNO�����VH����M�l;���D��]tq�',i����9erR�-d\��!?U1���D�2��
lS� ����H���G�p�۰a�\���U���6���(c�C,I.��y�*�D���;M�C�=c�����V���Ȼ؅:��$g2�E�g�����\��ߎsK �g��+�ggx=�)���2�e�P�0�!/e�'� 瘚�� �c�!�r%��HE�]���-��7f��s��3{{/օ�'yv
��m�Tݘ�q�5�L��~�jS�H6.�=Z;{���[n�e�������3�Z�U���W�gi;|������������D7�� ��j�]s�k�=)6tu�������{ｻ��gw�v�m۶-�@�?��?������n/�C\mo�ּ���\��b���[��o�&�.��WQ��4ݓR5���t�AN��C�R"`O�5��a�Idx�T7�J��֞H.�J����:;g�x��/=���}��oS��Ţ���g��ݷ:4�92������m�1�:�w�k���%����2�l��t�A[�pE!��9``(���
�p�c���/)"��Ѵ0<"-�:�D=4�S��6�&�oll<��f�:;A�nD��<
����̖��a@A�``dx,=�x � ����ę$7ȑ+@+�8 T�%���dwu����

�Ĺ�
R��#k 1�TR`��s�G�xр��~Ӧ�j����.�Fz]ċmr  ��IDAT���n��74�ѿ�H� Cn�����c,�ly!��m�N�Ed�n~b���F�Z�R/2�d�@C;��hca����>���E�����Q���D�r��^�"�6��w��I��"-��=�%��5�i@��d�Gd+-#d���X ��Ƣ���9������f��T�\�
ƭ��b;��%�F�	Gpd@S#�b���X7�T�d�H�B:S[DV���2,i(�n�:�r#ĀzF$��*������˱:y��}��͙cg�����Y.Qf�N�>.�he�ͽ��a��c,�ʳ^�+*~D;��wFΟ׷ T�R$6��b��;x����������\���\Z��2+~�����5o���g������ԩ�]�s�^�{Zo@K��]_W����=���U��W��Ė-[<x:�A�4��B�1�<x��_��_��/���U����}{|�&�y�k�@,\�5��al)�]9h�0P���/�u�I�P��kB�:!��Y����.���U�˄�;�0����;� ��0�T�:��#;hȍ�{|bb|����_|��G����!��`�¿ �*��en�]��8qr%b�/^����5PC���O��NcT(�@1֊�B��q�0�%�X�=�L�E�z %�Y���8 �u�ߧ����Ȩ��z=�W�|MZ��D�0�#ĵxRX$�E��y���$M�4EV5 ��������g/R>[�g޼�n������Ƹ�<$Ff^(�~��ظj��_�/�>�����]d�bR2�4�RT�,?��!w\�n|t�S����v14l����Q?�t �}��m֔8W�1H�s�ew���;T.�p��c3!#Ƙ� (Q�����fbm�&ǬeIȚ����O�R�D�q~`�)>��,ߧ�~A�+��&�Ќ��=�p�d( y�|���n����Ǿ����͝;'��E��0���`f[�Fj#�g��<p)c���	l�1���kA�sM���I��)�ub��Y����RMxM�8����3��C�g�S����L@R�Ƽ�o�2֍���n�s2i�ѣ"�:Y���;�D^�2^�]ҽ.���3�d�6�C{��י1��1��ю�x����Z f���s����++ԃ��{N�i�?�;��_�b��6<�獧��\���^Z��2*`��Q�n��ݏy`u�o����	?%B��C�%���Z�`����	ra0L*K�,���C���|�L����իA���[�n�h߾C�����]��3�v�ᑮ��6ovtQ��,�ݭv�йݥ��b̦�� `L�L�Ŧ\؅���2��$9r����_o�(�ޘ:�]�9sf_ܾ��C_��6l��åK����.�$-l�lݳg�{�uBV�\Y[�`���]�E�������"5���o6g�0�_�!��4�$9Ϻ�Ս7,�l�TE0`@à�=�!��q�A�zR�����8�Q ��!�X��!��u���@Fu܋����%��縞�ޔ�IhÊ�yHiH�]��t/�WT�W�D�:�"��|IT,h왕�7�Ÿ���c, ���`�캫췸�Qn�M�`@�}�v�3Rb}��e����$�G���M�� �.���3�o>*#n�t�����ڥ�QT��} =����\�q�T5T�##@��l�Yf\�����\#�ﵵ�ǝp2y��,_�7�p-U@ݾd�G�"��f�c�H���1�隍Ƀ<�n߾�����{���h�R6��Mp�o�L��49q����i��d#,��0q9;�&{�\�ݐ�oI�$i&�֍�T��w��<���cE<r��w�2�Rݜ`��KM�x/	&��8�uh�FwBi/�cd�Pt�7Y듉W�����s\Ep��o��s *>YGs�2�ߘ��Ђ�<�串���2���w�5������,}�2y�f��8np�M~>����6w�ܓ�]w�3���{�wʵJ�����LJCe���߿a׮]w���++ ���vXCat$�b��/<%5pjpٓ4E�:b��y������;�|�e��K�u��a�ظq�ݴ�������ӗ>��?�����"o��q��J_��Q',�0�@�I?7����{�<#��c삎�3��$�����Cv�%W>G��ٳ{jί���誫�~s����~�Z�t�8��Xl�W���U�رc�����������jJ+V��Ο�@���TJCGt
1F�eH��AC@f̃DU7˃B1�#04�P�8����nd����I���JE�G�	˂�@y`0&�Y�`a� 8�����N���&ip���O?�6H��"F��
ʍ�}���.u.n�DP��n\0�+SP7T�1q�T��ȳ�r���"PQ�/������iw����;�|f�`w������Ɍ���Dp	��1y�#{C�v���(������!a�ಃ���vMdL`Ģ�@Z���2ѩJck޲�����i=��,Y7��@X y��L��zX%�����3N7N�Mԓ�' ��>8"��|���q��7���ɡC�܉'�1�I���+5@��g�~˦���?/�F5�n~�s>�az><���y�.+v�e�<��<�[��毗�.�f K���d�oz�.nXd��O��7B"����Xp�(��\=g��?���8��>s��Yo��i.~�����s�ʰy���_㆐e�X��шn���!���}�P\3���5�Μ9������x�����Vi�ߒ�W�O����/�я~�9�ni����qT��+�KѥC�Zب,��W���뮻��`�y2N��y��L꿳G�9x���v���}���}�7�~��Gs���헱9��^L�8�B��@|�[��PH�ط ;���C^+(|�pY�x��Y(�o�$�٫���-��ϛ7o���>w�-���?��d��,x����O}�_� +�ڼ{��?~�a$�]�l�DG^��Χ�)��1ܥ�(A�Pe���E4�f����~h�}�8Ep�lY-�~��ʕ 0c9� ��=p�hFP�-�+�0����ah(����닒�`���PU���B��]�����P�b��Ts�)�)�WH��P��`�:����wc�1b�Zg��h��X�*Q�A�-$\mf�F�%�`A�ا :T��8z��\��8wHQ
�`h����
���� ��9~�ƕJ��BLR��J���tu�{ȱL��ԩ�c��~�^7���D#1��d�P� d2��D����{Y�6���K���/&��rY����Eznz@�T;A�[�x��3���2�=0k4�s�um\UJ@�1aX�0na,��Ë����^҄ع>�Fs���1a�2 �a�޲7Ӂٯv���� �]a9 *Z�V�'-i�s��t��@"��c�*_,y���X��X����W��s�8��7�,�U�As����s�kܴ�
U9��=W�З��ʦ����뮻�ťK�������o��ʧ����eR�a��OX��o��'NT�dU�T**���6W���hG��^�ˌ���G>��o�����d���2��Y���Ϟ��y�޹�޳n��=7�8ub����7xc�]�L�0f��J���&�_��,]����x/9M�*��&&y�]Y�h�ι�=��o��o�v�m{n�馳p�����
�U�`�<w�\���<����74,_�\_q����]��12�V�=�"��#ST=t����DQ�$��`��H�}�t)���������No�N%���`<����"�?�i:�[�&�A!,���EL�90�U�]����t��g<�:{!h���zM��Q���v�[@em5�I���&F��mA�Ǌ�i1�7��(z�,'�RX��$ϔקK�F(��1�v�k^&�j�*�?�:΁Q�X,�O���Z�_�?i�����/�C�, ��dp_u� �!�w#����x�z�q#�z�=�l����I�@�����E<(��}�Ր�c��S:������.�x���g�pã�=�|���qW]�N���������El�4��0�Pb_�>�G�nf��>űBc=�����0��z�|j��`bǩ�1�.���A�4��� t���}t�d�(�K2F�Ń���1�y�x�.;��K�8�?3�I|L�X��m�g�,_�U��93�a�$��Ɩ<�X0���N�]2
��5�x2�"�F�})�h���\��6n��֚5k�/?/}�V���VZ��S^�pֻ�{�/~�����o��ܹsE` ����M���Dj~�Fm�������g>��Ͼ���.
V�T�׾�v�6�t���#G�ؿ��e0U������d��9�(���E?�w��{ީS��ɸ�ױ�pۀ�t�O�Sވ*�c������:��Y����_�v���5���ړk׮=�'�����7�����o��Us:t͞={�9v��c0H�,Y",6�9���.���� "��\3�%���	XV)m��:U��8]M�	��.g�1m����F4@�NF��y�`�/Z�ȃ�v1�a�3_s �@Y�P��ǹ `p;����$�}?��~��I`��8 [B@�3��SJ��!�zZ�A�i���E�����F)NT��b�5�.=\ڎ��7�4�Q�▧�4 4f�[�hd��,��T�$1V
��~hw߆�'pD�1��C��@P�D�x��V�b])F�g���3�\�=Z�'y�|=h�Y���.�SC���V-pj�Wf���W����H3�o\�"���  *�p0�����X=�����p�={���ԍ��Ƥ�!�-�ϴ`�_����ǲ9 6̀�X�ce��8v��Z�"?$ޠ(j�aP�&)��6\���16�;߅\Ϭ��B�yxn�M*Д@x^�~�z�,8��b�o����|o�7�J���z��ۍ3�f\�x���3̓3c'^/�f����St��/�d�rqV�]��h}	� �U�|��s�Ε��Tݰa��6m��c +��k�V�-+-p��/s�����|���'�u��%�0Ei�rOr�R����|����l����N�&w�hM���]�h����m|���M F�,:z�?�0�
H\�?�344�������o���_cCg笞e�VT�l�\-�+����;��=u�䉕+W�{������U�F��U������,��_����ʃ�y�O������ۿ��˗/�����1��Cn�)7� g�4W�$ǌ1�d����B���1O�4��X7�>��#�`�2��(ZW&���w� '^!5H��U7��F-��i�B	�ޖ��b�p��KeB$	^�d�0	Ǐ�����=ݳ][�#�ZW�J�
聻�[ww��A<�	��F�f��-`+�	���ۗ;����F^m����)^�.�*	pD�O(�8\��ot�k��J�!b�]� ����}`P;��I��> Ȃ�&D�IP�X�/$d���Tmi�W��$�_\�R�Xƨ��_,�qҢ@6Y��Ҧ�����5.Ēb��KËsx��h#�S�T�g��'�]wݙ�w��n�u[���~����C�j�&�k.�$�F�N,3�V��E.�qZMP��2�a�����{�Bi�SAƟ�T*�ᜳ�nq�-S#���1�qA#h����vS�<����̗e^,��r�Y�}�]�gJ�"��Y�3]R]��+ٮ��`*�s���m����a��l�Wd]r�� ��q}�?�~Ȁ�<�ō8���ARq?�Y�b��7o�������UZ��PZ��S\�h_��/|�����j�mIZ/H��T-e>�\�v*&a�E}O���Gy�����W��~���)�^���³��n���S�ο��<~�
�����Y�ߍz#h��}�����O��\"΍�/:z������>������W�Z���[Ԏ8�BR�^���hG$D4�@V	�J�E���������B��(.[��E`��&�ٲ1
��!��.[�n���*���[N�.���ꮳs�(�y�\�U�?V�q�;<pT�9i4{CՃ�ޤ]]�K�u0j��'Y]�x  ��@�'<OU�q���@}��s�� +��3q#
�*�X�{�0F���b�þ�箁��4��$�'��$��L+s�(�B����Edf�|���*�p��J�� �x"�2
��̴�3�F�������V��f}��hΫ�׬�����Tk!V��wv���'��p����(����+�{���ɩq&�NT�#��Q�1R� �F
bB�S����Bѷa���|���q��-�� S�h� �?2�g6__�Ύ��#��s'���a9��_���}\���������������7�䏩9��������s��B:�Tc�ɮ42���pL�o�S�1S�wd0��Ė7���w`��8<��>T�\,�\Q���~�a|� OB�@�x����n��3�`>�;O�cQ������τ5+W\�� spHD\�K_��;����F]��c��_7����ڂN�]3��9�2�x�(���a Z`lgܚ=���>4�)�4OɃXs����e{m윽ntG
g��q�$�t��s8ߙ��ncByM���p�N7�$�^
��.\��k���e�N�����A�*��i)-p�)-:i����^{m���@�7.K!	�ԽJ��HN+-D%,*��o����G��[���=�k����N�C�9�2p�W��s>U;`�#o�.���㣏>���^���]Z�r�����&�,��拖WZH����"w�S�`1���V9��40����#�C�12(u)Ԥ�L���OA/�hmm���? ��]��bh��E%D�<�مVc�|}�cp 
+LED��C6��y ��zRi�ۘ��'"�B�>%~QG{0& �<�.�j(G	Ϣ�����X
a7�F��˸L&�l����C�.b���Fc��Lx~�Gh+�7��ӧOq�Χh����3�:��W���0A�R����qn!�h�)���BLE�o�AT�t�RqC���;>Qq�=]�\)�$�թ�svO�Ļ�(��L�������g�/�8����G�U�Y�$�$X���)i"$�TU��%���0/��b ^5�^S��dhlH�csxx(��p�\�³��G��q����Jn��F��כ�:}*�`�X�>t3�*g ���H�7\4M3�������1f��m4��{�u-~��θ��?���5�u�q�����8���?j2��d-#�ψ��o=&7�z����G#���B��l*]2fɂ�ْ`���7�e�g��}^�l_�E�h��ܹ3��Dq�<����u���RI ��S2]�b
�DWA)�e��q/���2�L���1�򫟳1�oݺ���}ǿ��[��U~�K\}
K#�Yu9r䶧�z�_��=~rk_zW�q���+���L|���FU�������[o���k�~�_s��P�>��:�S
����޽}��7߼���C|��^}��),��aDw��� "&�s4h$�9����GI'S��	]��.��`�74g�\��=
�F�*1|5�H��bI�?�����@.}V��F4�!�ܜ9s�'��P?,����#���~>�-���@�mƟ5�T�]v�aSu�Pê�]q�MC*�NN'�vŝ�{nw�	�F������ݦ�a6����^�O��`�vS�'ST��=<�o��D������ �T�/@��Xk��,��,ZT�Tw@�N�+�WI)��n9�UH�bo�G�ߘ��Lt1rb�}G8��	�+����$\�:%H�U��#?�U|݇FĵQ6&a�	㔆[d����۶}6��W����q����t'O�L>��*O1XL6m�lg2n�$�(�~�؞���ʁ��kX&W�n3���#Ò��y���A�"㖧�P�� ��1F�5�q}3 ��H�lR��4>����󛘟d��O���������7c��-�lVF1_��� ���k�K�߹O�Q`���eF ���Zu�d�d�d�mn�%���	B!#n2Q$�����\f�6��
���͛7��z���y�.�c�J��֖��t�������g?�w��ַ�:u�T)�g�>Ä
��ߨ���7ހ�[��b�|��G_���zժU
-���X9y�u�?zÞ�{�����`S�X�Bc,@ D���]>��U�F*Ɏ�B��`D`ø�ImJ�5)`��6��v |ԈM����G��R�F|�� y��Қ����C�1Q / K8���3��׏'YX�7l�!y�����#~ς���ȅ���Ӑ,��\�%���P��'̱2r�U�8�v�7 ȠL���V���|0 c�=��2ڎ	�𬡙�wI>˹�yƕ�1-�R�Qc.2�D���P� '!f
@��	���q��Y?�-w�����P]B�}��	]� ��j	���� J�i�Z��=]!c��X-�!���aܪ�gB&��Db��O�$J�����4�B����zlxD�z��GM�������.ng�զ�-[�K���uw�q�����Ξ=�8 ��0V(�B����븜!�u��\�H31*�}��2���� �јƐL3�-��k0�Ϙ[��At��x�kf����rP�D^&#n`(��8�	B-�2��1h6��e�L�����\Ǖ&��Uo���}' A�(n")�E5m��;ڲ{4�p��;b�;����̄�������t�(u7E�%���H��?���[��r���<_ֹ�
%Q�F��x�{U��̛�7���;�;E9g�2���8�L\A��z��069eP��c�.c����*�/��,���z��92���8V�z�-M���V�>�++�l��$ކ�5�\��ƍ����������wYJp�{V�V��5G�}�?���@AO_d�`�j�����*N���2��Ʒ��n�����k&*�R
��(�"ݷ���w�}��={�^(�͛7��
% ���f�X�^�����3
s��eCcy<��R A�y2���h���w�)�M#wΜy�ơ
~*�>�v)ɨ�3��/QJ��ƛ��H O0�7)�\�XKB��\-Y�$�#^�T�[�l���/��µ`�,��8
מL, 	w�GG����H��`��8<�5�[�,z�M��\����̱�w�����xF�2fx���AcD	�,%@�qCߪ�/��801t�DZ����hN2�[���| � ��#-�u�\����S�9{F@تU��z���6�n�3&:���sM8(���$�����L�%���	?S#U�U���}��]d��B`�h���/FĽ1TM�Q�S"���FGGD)�^oHޮ�$����֬Y�v�����Kn�+��*��'���c|6�nKC����U?W���^�������%뺊�J㪺�~u-JL�D�~+e|8F)&��lX�~��J����[Q�"��!�m,�A�d���M(�K��a��2�+��i�:�����I׶T�'կ}����y��	0�Ւ����܌ե;0��$	N�|�b��p�������lڴ�'a�z=T9��R��������<y��ۿ�~��h�ǗI�������V�>080X�$��W������wܲ'��K&������_���?��;��E���U�6Cr�L���t��/�V��k�Jr����|2�í����|pP��Is�`�|u~-���ӆ�6�[���ڠ�ށ��kY���r���B2U���|��/d|����n�ʥ�R9r$�wI\�x�� �effZ�#<湺�-Y�؇��������� ���ј@ႀ�U�VfSS�"��M����nP[l5�>�+ f��yt�X�`�p�h��z���|%�Ƿ�퍻茡�.�x�4���r���7�����2s,�4i��n2����t�c�څ{f�8�#ԍ'�,��E�g����	�70�ϦF)�"�)�W�� 琥C�躒Qi��8�r�h'XU <�)vi��ͻ&ׂ�B�lH��$�	u���]�pA2�7 �i0�-$�u��o��PO8�	W�P��{�+_q;��֬]��%w��a��Y�����%�;��u�r��p.ǎ�4��[d5���낋�kǏz����?�{�z���kY+^�-7):��9�P���M�m�Z��_`YP���S�2-�ZY^�0�?�\{�
(r�j�u91
{���ʹw��9`��Z=�5�ڣi�I�s^��>+�%K�#�N7�R����kȁԯ�&��S�|x�ǜ�~�̙�ƍ?ڲe�+,x=�Ε�,e�R��ߣ�%���w���w?��P��n1}��8d�e��[ayԝ��ҥ�'��W?���;�Z�|y��}%��p0�6����x���v����������W�Z%F$�e5�F�\I��j7S�{҉��[)�a���vE�` D "��B&FZW��%�8�`*ѝ+�\�=pċ,�H� bjP�w`�.��0����7�XO|����ذa�H��:u�MMN�����!D�g0�	T𒟚�+�~�K�L=�q�+$���z�:u̤=`�h��ʝ��hT)k%�I������i�0٦SC����(�R���Ս1N�� )0>�h��ꥄ�*��U���>�<(����G�/���l���S����'�S��U�B1����PWFOEE�wdb;I`cf�U懆G�8�������Jf ?�j����鴃a��P�7-w��I�\W@���_����p���7�֭[D���?�� �}$�2�-2-�l��˒����O���߿\��yLʊ7u�s���>
Sd]���6gr��e����Z	M;�3�H1�11����$ȶ) �� ���K�*2j���V@#���7�[a���#��T��c,/S��MN�Ā�~qZ	dY�c,�i�;�/��u���&�&��*ض��9f���a�6+N�>�X�z��6��	�]Y�R�TJp�{R�"X	F���������[O�81cE%Y1a\Ze@�Fub���¿�7�rۛ<p��H�[){~����fU ��������}�֖-[��K�
��4���{��-L^~�Z�33��ت��N�� P�{��jN�R�|�c�y��H֋�� Cx!�|��FK�+P?�@P։q;I����b@O�l�$� ��Q�Q$3���Z�rE8o�$
Ʊ觑为$IiG�9�䥎:��0���p��Q�?��7<�hc�5
oD�#�[xR|�D�HF���gLc��C_�Y�#�
�#d����{��17B½
3��sf˙��o��j�;y�YQ�7��2�e��F�)+%���=~��ԅ���T��o�H|J@�z�A6�ʊ �+t����jG�\��S	0
m75 ic֍D��dA�bΜ�"f1	iy���A�B_�$�lV�h6d����������Ȯ�v�l ��8q\�E�*�W�31VjTp���>�Z�?������*��Ou.�amx�<E�^��3{^19nT �3����@�l���	��~���8$�32]�J���}�#�a@C�2�LQq/�cv��ۺ�����B?��;�c���*�g���gEF�O) �|�E֯�~['l4܊���l�]9 ���^A�"�o篻�ז-[�t�3WJ�%WJp�{P@��o�G}t���k�z�aJX�`�� t��މ�
^���%e����z�O������ox!�te��J��`��@Ńo���=o�����6ްa��a��![�KJw� M�/1���$��;�IYC���V}M�uG����+�}4@ �ꋠ�Ri�3g���ꇇG�u�^A��,�>�2�')��U�[��0����/��*��M`N�� � ��\�k�:uB��!�=o�|�>X���vS�&l�ϛ7��ns���0�G�!�>,9z:���6�rɈ�T�Հ�9�㦃h�X���[Y�{����r�%��y�!Fߠ� �4�'� ��A�M� ���&���t���T� ���u�� s�Vx�q]�)�^�+�&�E=�>���!iXG���\�?��h��p���Td6m|�[b��w���955�l/���V�jH��մ$�j̅�Wk�ƳA�Bmu��@\Q�L}F�Ao��6w�}���۷K�� �}�>���	�q�����kk��:>��JX��:��̗"�QV �M��]�#�-�076_\��02���2��7���NV�.�ED"*%N�T��S�9�k� �k��I����e9�5�a�6�����a�߸u&���5���Z����	�ak��':~�Z���.��i�f� �b-��L����lg��,<���ee��2�o
Xxu��9x�C�C�	�G��a�ɖ,YҺ����߿�׫��r�,e)�\�~�9�X������g�Y���a��s:*�A�+��0��R�k�ڜ9�{���v���`蝭�ꀿQ	/��0+O�>��o��柼�����^o�Y��J\%�.x��)���>b� zadhD>�10&a<W��I:��7��tȲJC#*�����j�����=�jn��1֙
�H�;1q�@#�* �`#e���'jn̩�
 �2�^�'N��?uK��Aɒ
��Q�-2��Q�[�;Y/F�g��`��7{�Mڟ��7��ڭds
ajh���4��H�}��ɡ�������kA�}���"�^=���&G�P�U����M�Eͩ%��y��ql%O�c`��(�]LN�f̙�D5I��_�o�~8^lb� T�Jc��L�I.�]��I� �!�V��s��x�p6ڭ���F��p'DΫ�KSnF]�|����+�}睷;(�q��n(�����?�󼺰ze�ю�lP�M�9�y�h�昪�O�x��Na벌����+��0�9�;�q�Nt�|>� ��X�/��ƻ��Thk�#���+��^��4���ӲA���(�6g�-c�s�϶e��P��7�Xmv�R_����~���:9�;��������m�.ec�;�?�6'U@ۿ^�>��X�+�Vx����%)EΞ=��Ɔ^^�z��a��E�B\���)%��=(gΜY�ꫯ�������~o`T�0?HT'�b(����Ȩ��ɢ���ڹ����/���6m:S.x�Y	/�j02��:uꉷ�z�� �dW��(JksF�������ٹL����wY��-�}1ƅ1,h�ku���.@:�F�Ӎ��PRP��v�U��2�ls� 0�\�-v4_b� ��V���m¹]E�Y?1_��L�����D�^��)	�\Kd��UI�u�ʅ�@׈�p
�{( T�/�QE�j�5����TRj��t������|~�o�$�2�W;��-�1�o��L%��CWCn�|tKLl~�8��!L�L�zF7Ke��*`�o,�ʁ���X+a�L��J�Ԙ���h���i�qd<�+�����%C��r�Hn�H�l�ႛ�� �&�����@�����z�-�;��'n���� �O�:�>$���z�Y�$#��oN?|�}���.�V1�E�eX�Y湄��t]�sJ*F�ή�m��.��.�T����6ސl��"��9�`v�:���P%�g�		Y?�W��H ��m�������9׿�D,*�ж��d�O�{��Y�l���HU05�Ɵ�͂+n�w݉�y�k��'�J���. :>>�M�Z�-έ[���
k�����+�
qY�ҷ���wX� ����{�'�|�ˇ���1�4A�,|X��|8X�c&��ͷ���C<��ڵ���.�L�%��Px	��η�~{�/��6���֭׸U��D#��QTeKb*��~���D�U\Sc9�zi�TƝg�4qw��qG5����(6Q@m(a����d�W���f��;�W���ܹ�R��E*׈_��"�%��!P�@�pM��FY1#�!�k�5U�f&Epɒ�bl_�� p;k�����8_ܹ:H+АX�p�"���j��u��!�.�kx�l���}�Jk�܎7
�H Px��a2�4������W��s��"� ��@��_$T�k�iQEpT���^'J�?G�?&�=�M�.�Y���VL,@�ndtD6c�va�����(mq�#�&shݲ�.�gS�0�{���N��`��
��n@�\�n֔�&�Z���Kr�2t�# ۾�Z��c�����͛?q ����46 b������uB��|��@��E�����c���3�3��U����&ۗ:��9�UxK�'.����.e^��N#l�9ǺJ�S� �ދJ��H`�1�= łA�i�_�1�Y�Y���g�sR�m�
 ٌM����[�e��
�́G�O����8]A��Pwѥ�'>ʹ#7�f���
�9�xf�<��R&<�����^�x16i �S�~��W?�	��������JgU��\����wX&&&?~������ߋ/�H�<���;Y+D��S����u�*b�n�q���|�[����\w�{V��L���F%���#����ݻwoCPۼys�~��`'��ÞĐ����qz~F�A�d	̋U∪��MD� �!{n�T0��HĴ���XWО��`��J\te��X�z��\��y3�f7&!�+qB���b��*�y��i2a�Y�hq�ƴ�@j�w�(��PJ>+a��-�c@Y#
�������#PIFZ1�S�r.j�Y��1�ͺ%���.4�1h��K��1i��$8�6�0��C����V�#Q��Y�e˖9&�U�H� ��� dp�Ę�>�3@ъ+��b�p>�e���YP��,��d��'L��:9?��Νz�FX�(=_1�쇮�G���76�0j�ʞa��?�5����
c[�CQ�+k7��lC�c��U����{衝nq 铓S�^y��)���;*6!��Y����`�3W���o�; �����;X���9�Aօ��^�Ջ,���'��d1h���A�*�EƆ`�m,�UJL�րW��YWݸq�D�Mo�B�s��֍�����{#��s�W�#����a�JvȀ����L�sqc�*�2�j��"��m�S)�#��s��΀F� ���J��!����6�8c��=$R������9�c:�5+��ن�7n���K��?��%�*KY>����wP:Q�l������}�ه~��o��ǃ�&�k1~#�=X��7��lPeS��a3w��5�w�u�w���,�wɕ��.��xml��W�y睻_~����h�m߾��~�����6m�i��ˑI[-�d���rn��?]3<��i�7�� ��5�Q�����ni4�	�Ȫ0�+����EM.\����rm��y�$	F}L<#u�0�Ui0�<�+���f^/���N(���-�y�b�^�W7�L�
1���\2���v�	<���;����T�{���RW���"�����R�}�� ����qMN�����x��:����$�A�
����V\@�B�1Ī���HW;�-U�K*�^%�i�Ұ�.Vv��u�]�Ȱ�������"Kֲ(��/�K�#�Y�57�L�P.���4q�-`������ӭ[��M��a��mE�P��g�qt"�Q�|p,���1)��|�w��q,^��|H����s��0Y���,�֣@X��͹�"`;�;F�ЮoxY&��9pd��,]�-C�AP�6`�������>x�I�P���͏�L�1d�g�}d�KL��:7n��>���{�k�e���|t��t�����hb=�� �`�L�Z�j�����W�X������R��|b)�����}��}�?������yX2���&:������k@�p��ԃ;w��o��ϻ���eS0*��|��7�Xw�ԩ,�*q��` �6$�����cI78���A5/WO��,��$�-�$�]P�ӎ*^�ʨ� �禠�5�.)SEP�NQ|�@�ŋK[����Ɯ; �����U5ü����s����
����!�
`��E��Ѓ5*ӎ�4���#a6XO�� n���%���>r�4V쎷pi���H��!��PO�A��n�Q�^�q��+%�#��y�>˵n�:i�L�D�:;vL �q�
X?�����
?�����y��U�"�� w�)�N�Q7��c��H��H���Ec"���L�.2��qGN���
�B�OR�ھ�x��)�c�k_�=��cn����'��V)P�D_�Մ+i@urt�	`)�
�2:��jC���J���2W8?kG&��ɦ�1�R�U�mu����Cc�Ȏp��g�ޤ�-����x������}ƺ�/s��&���xL�O�����b��)˔�D��^fl{����+����Ϝ[Lj��+�z�Q-��l�M������9�RnH����c���5��dɒ�믿���+W�����2�,e��W�s�"��`�_�W�WW���{��E�:��jj�H��!,�L��К��6԰���{�z�����kW����k�0&���LNN>���~�瞓��͛7��[��1*jp��'Cŝ{}��m�g����T�(/x&�$s�U����ÏƎӤ�1/��]������Bl�S���
��1M��R� >��k׭�FGFD������[
m���F��s!� �$�0IB�Q�8��� ��u�&/H?a~�LsHQ|©r�5k՚�����q	��X�ݒ��5�����ʊ�"ڄ���� @�>E���=P�
��+V$m�J�Cr}0H8ǆ�%�u�I�0���།7� ۡC�xMK�6 ��9�������hԂeԹ*�ӰW@%����Ec����9U6�`�3���y����62'��w�k;</�pI� �$�΢R#�����s�N�m�6�i����a�'	3\O�膇���3�&�M ��¤�h��O^F�p�72�tU1�̜M}DpB�O ��8�v�!{ȍ9d�T��'��u�G��@���y������s����_�#����c���z�nw���x0�U��t}���"*�s.	5�J&��E���*~_��8��[��B�
�3~�(k�@/��q��s��a[a�S�v����6�0<߇\�X��,������/sN�;w�/��ş���͵�A74<*�#�!h�ϙ;1n�>+A��>��p�v����=��W_���/�X)��e�������~�����3�ǎ����`�Ɏ���!�NFj�иp1" �V�#R�d��6�qB�����ŋndx�	eW1C>�/�`U��jK��lfZ ����"��B+)�Y�ʑP�cp:�Уy����O4��Wu=I���h7��Z��#�#�
�
����]X�F
��qNC�n�"�˱��ɚ�.��y+�\UkQ����n~����ͱ�[��%0�\��7�FN��q�fN���͆��������y����P?�%����g I(��¹ÈIr}R��%1m����+��a�N\������a��#��3X7�ȜQ�]��:���	u���2��Wƍ�̓�c��j�@N*��o�}�����!��U���� ����v=\�@C�y '�{vf�g�U�m�fB������f�MON����{���܎�F����������Ȱ�$V���c[���Mɭ����_���j��b.��A`#�N<��f

\�ȴ�kU���g�4�*��ɥ�/0t���"Sd��\`����`�*2~�|V釟sS�X�l�x�l����IL�2��z��#�G��"�d�82��Y��?�߹������r�IʜkKW�4�q�v��eg�#m�u�M�z��a����]���eֹ(�VX��NaN:th0���n��_�_���o�s�X�W(%���J'�Y����������Q�䲡�A_���蚃EL�~L@�d'S��}��{��v�M7=�T��,�z�K%���>v���Ｓ{�k����|0nw�ؑmݺ""�]��!H���R�F��}IV��%;�.�(�L8���Ν�Yv��DQ
�!�eX�BX��9�l�ҋR�O@A�p�Fyܱo
�9�	Iu����F
��A���)��W�5kV�}�.gI]�8�o����;�� 7.a�F`�xp �ԧD��^�1�r���X��nm��,��i�}cW��P��R�D0 HW=&�+�$�`�C�v|J|�:7{E�=1X�P\�g��@���X�{��s�c6\��
�D��!�4��n|��.�r߈�0J��ZY�J���� ���7�	�1��Wը�)| ��Zݳ�$v4����C��ק'���l�j�x
󷅟�5��
�MO�"��?6"���7ݣ�>�n��z�ɹ���ڠeǬA�Q�H7%it+JЗ�0�l�4]Lv��X�ۂak`�WDg���$	���~o�[��(ۥ�w]V(��� �7�z�>�qK�+2W���U?-&Ν�v�>���i�Ⱥ��X�@�c�,kt��IߥzM���1�F)�u�}�$�f�����]��h7
|7�U���dSmx�|�ԩS`�&6l��ԪU��&��o��/����,�R)���W¢�v߾}��������`�-6X԰�MCIc2Zp����}�1Fb���~۶mOw�R������Ƃ�������w^|��1�[6o�j�vl��Q�H����' 7]K^�I��/=O������Mb�q���MY�v;��&N	\[���V2��;� ��Tm�9���9،f���\]zp>b��\��׭C���H�+u��ߡ�Z�#1b� �P/��ł��x��+�=�7��!��UM۟\u�ޝ1Jz�ÊQZ+c(�o��t�h,����K�4GA��v��L������rJ�˗/�qs�<a�O�6
���ϼ�n1�6�� �`�v�%Q]����_��k,� %��1P�.d�v:)��)[&J�(��2�3z9��+�u��(�!A���ONN��G5�Ձ0IM\�bb��L�b( M�:4}���1�@܍7~�=��������ȑ#~�޽�q��6�g�r���Ev�~V1�r�1(����>+���W`杯�>����ٴ1H����Nk��@��ː�8��}Ḓ�e9pX�1視�8���.#�<�K�-��g��x�^-�0}l]{���}��$F.�q��_2��5)��Z/7��Ƅ���X+���? m��v���b�"�{4��e�R�LZ�1��L����\ V{6o��wa]ŕ���R�_����s*�`���������-?���n����` ���N-�y�V�o3O��i����iTY��VkӦ�Ǿ�կ���O����*�"n�#��s�k��6/�XF�n��l��
F�����[a|j��V��� a��kq� \��U��0n�\g����2^�+Q�@�Id�Tq/u3��@����E��Ipy�4;=.;s�\/�/q�B{�=�4��/W1$g�����ЈF9q� l���2)-����@l � ��=S��LW(�H����tot�Hf�TzX��Jޓ�� �1V<��
cP�
nȽ �x�}1�]�� �A6�����3�`l@U �2��<�1��2�DІ���5��3��4q�j���c�(x�x;v�>�uq�
�ɠQ�nG�c�>A���N���Q8�*��)�����6��� lF�dL# �8#�g�VS�(��w\w���?�Sw�������������H��52����f��e˒�s��5-4�{之ŀ�j�j��&�M����'p&���ڑ����C?3������{��˰f̥���e-�b7=��M����W�g��b;m�-�� �p?� rO�����-'o�-�C�f���+�k�,[��:����}�熛2\C���I��Ԃ́�4~��jժw�m���K���?^�����+%��-],�v��}ۓO��_���?ʩq]�.����_�"��BW��f�Y366?�ַ���;�x?_�%k���П���.M]��w������+�;V��DE��S�3~��s�En�25*��c(n�Y�%��:%�B��@\	l�8�-O��$���k�,MH��k��l�6��ap3Y  9F=]�'�sR���g�z�@��`�� �{U�� k5@��2�fQ��kN,arL�@��/�X�A��i���*�g�� ��1��2 !8��`F��G�N�����v�{�a��GQi|t��B;�?��;��p)�J�/�� 8�)���;G�1�d�0b_ �a��(�E�,��n��n��*��c1�'��-���w�4�mQ�}S��eίV+�q���qފ+e�E�!�m��8�F��[�fU������_T(���݇}$b *���gFU��c���cdؑb�Wν�^���֚�[�<�ި��|̗�vE����N��ҦB��2̣}^�,�r��[�)�̘��?�7���c��>$]�C���\����X�n���S:�����Q����n����?���/<w�sf�;�]'�9!&�:ɟ�Ǫ<����'TI�<'c7%Vg�7?A�/gFA�8=3��6�";~��x�&�Iw�&����HyՔ�Y��k�b��2�z�
�f�Z`�G��q���٘�H������z�7z��/���w�0a�� �,�z	I���M0Ԥ1�ݑ��Z����O�q�v�j�� n�f�����~p�럻�����H�q&7����~�{�>���X��a+N�%@I1}Y����b�l輜R�?�������]������Ҫ���,J'�xؒ�!��FjfF�ѽ��5�@����C&��:�^y�`��j�D� /�^8�~�e-�/��EkKN�kYF���t����TS��d�u�����ngJ��T���fB?C;L��ʇ�3tmJ�cN&��T/z����0܇�&MN���r�h�py�9�����Qg&�
�	s��3��R�:di�@'Z����,�w�*�-�V|r�|�_��ł
�����&�*��p�l�	WzN:_98nv,2|/`\Od� R�<sЩq1}{����NT4��`�n%J`�����$s&Y��a?�vԊ!Y�N�*a��&�o�M�:��v���`��G��l��`H���w�Xx��B����V����31߹���.��j�Ј�>@�����)�s裥����.��-{<�=r���e鸣���.��]�l��#8�$��Xt{�B�����D�d �=\��M�h(�?3��?r�\�Qt����^���%~�7!��a��������[�';>�<��C'�<%�_nhVXa��p�B����K��7��9�_�)�k��D�p?^���=��Դ��onuœ��3צ�-2�$��x����D�O��6����C��.*�n"#��e~*�!�fr�JIm�'2i�n]�b[�dR�,�@z�o5*(ܙ��m_�N*���7�X��8<��C�����C��k��$ М��s���fr�@-���,�q%)�6[��&�C�3�5�M��`&rĤ�ܭr!�Z��22	#E�Ƌ��e�zt�="�,��^�\��ԓ��J�ri+n�5�'+*�8�]�p-�V_�)f�U���X��4>c�]GP�6����tu��n�U���v�W��y��[i�$6� $B���Eج1b~�<����H���w�4Ӟ�ach��b����0�drBm2������G�s��N�G$F#��#|�n�L��f������{^7{}��-�[�s7y�9D�Z��������qO�_2܆7��^p�;_!q���q?����Pѵ�6��ej>��Lk=�?u�;�Sb�;��s��6�9~��A=�Ѵ!�se��4$��ȫ��`���I���n�V2����$4���aXNQ��I$�[��a�_w��*��P�oƗ�{��^��LO�?�d�?]��!���gQ17Gsg��cw=߼��:V�#�&�.7K�afm'�_M�nl~_�D�m�x�8�cvJR��I{�\���{F��6�����N[�\{��Biy�M���<d�#�%�1�Vr>h/b~Ⱛ��<S�g[J�J�E��PYAhWY�/ w*k�2?6�Ё~��~�M�ӞN��A��n��R�Ɍx9�;ݷ�G�zB�ɺ�f|�3�һBJ ��b1�gYC~f-b�����ن���p� \*$\�I�c�@��p"<@:��x�C E~�%Z��|V�UH}&:�nm��c��ɤ>�ى]�w�������� #��sb��[����B�,�5b�6P���LP�3i0UD��~w	��!�)k���>����Yx�jB������S�Eي�~���5M�m���1�I{do�k?�M.
V�5������Q2N��d�꺸�'4Z�s����Kzt�"c��l���,o�e�K��M#��.�T��q���<[e���:��gM�u�0B��Jw5������س@8*��}J��ފ�Ƹ�"@�2MA0[k֬&'��=�&x�.�P&���5�\�������_��O"#=��ųg��m�����L�?�ۓ�I=0H����S}��p�2����Տ�d��9��^}?�:xM?i:�~B2u���Q����K�W�y\�����揅��n�11񠙴Þ������$V��������q޶�z?�H<3��+�0��۱<5M�|B6ꐚ�jo���͏Ⱥ��CC�w�􉰧Ӷ�&�!"�P)Wm�&NZdv� u��xx+gdD�e�#a -F��[G�U�iK>Gh�U$y�\�)�<��/���d�.�����ޫ�,����D��
�{9�}�j|�~�4r2;"=yAB[=LS;4ORUS��3YQ�f�-%,�TÜKh톫�M戧�����X>�E���KwV�uHѸlz�e#�Y�{p��W#A�O*�ѡ8i���q�����_=9��R��J�.����������+�d����@L��`������`���N$��
�0˴��$t|Ǡ;D����DA��u ��7H��儝!G!�2[T8e"*�/ɷg�KulB��,��[�z�Z.9.��É�5w��`TL��qe���B�#"��e"�QB/�t�d�����d��w;�m�����=�1g�>��D�����?�ɟ>��y���K�|bS�r�p4 �_���|��-����3��5׿��js�ў{/��}�G�����5y�N�B�Pw��T�duϷ[��-=����*t��'�����h`��j@M���7z-*��� {�����z�G���[N�,��u:-}c�󳄆�`���Ħě+#��!��iق��xO+'���aF��<g�Q)�Eu���<�i����l��@��\A6���j��?�v�R5e{&pxt3�.���'��cj�����XƊ��9�l$m��U��lf��I��O@d#�p4{��ک�2m�z�r��d���̉��	#n��������0�}<��x��	�O+1%Ő�z�R�kp��&H���3rWkrݒwu�X��+_�I��×+&_�oߎ.�@;S�g���l�lH?*�j�O�+��.���I�/x�*ơHm�����<1�`�S[��%=
2S���N���j�!j������� ܎Y˄Sd�c���kw/-���u��®E�$�-

�,ImGY��]��#]��C2%!���ీ[�R����>	��'ro�h{`�u����`2'�.������
�2dGy�=�`-H�l��:<wd܏j�;y|B��	!�ٺxxˏ�i˺���̾�u�+gW*���d"��7y����^���Bl!QD�i�_z��k���I(��,6^��jq�r�֧���Fw�����*�k�M�ۘ�fb%�����!!����bK�t�ñ�6xF\=�w� H�t�GHk^��E�f�8H��%x��+rrBG����,�1����������R����l�V�@*��4GE����g�
@?�y�|ַ�\�v��{��4[~���)>Bh@��af���y�2�:�v�/����}5z:�v��ز;�SP�.u��Q	�B�nH9C��򌛝VT����,�����0��V-^<���`�e����J�>�{5p�p/ͳ/O�ρۿ�nc�7�3�`�������?ّ�u�!	M"�N�m��{���W�*h����]
}��y ����v3g*�/H'^�	�#Fʈ��^!a�(x�R���zJҁ��w�4��E��k�\⿶��5�Q5�įYGA���I����	��͊oˉ��\�#>��3ԘM����(ہS���s���C��3w5oO�o(���$ŭ$XFL#�\��{	㏹#��߷G��l9�w���&��F �d��D���
��2l���>�j͉5̝FJ!���<0%KC�T.���7���n�Fo�|�C!u>�C�i��O�)%&˂�ڪ�	�, E#����`m��D�0�	�`���[ᛅ	wL�*f��ߣ��\D�;]�Q�C��H�Ɨ�OY���7�H˞r���j+��=��՜^����l�r����7Ѕ׏Zw�����;-_��g�_��.�IA���e�݉$������ah�Y�ls��mG�ɣCv���	� ��	�`>��N�����P����>�2Խt:�����@���ČԮ��C�N۩��$X�IG����}���CN<+���2A/�8J�^ٶ=���S�Ǭ�y��ak��Q��.j�#�����B0<���#V]�4�^�����w��|���I������0elo�.�i�w���t�bu<��`���y_��gb�D��y��&�弹p�L��D#����{Rhq�@���_��w�o�A�;;���/��V�9�A�]��F���Lv�_�c�m�T��0W|,FЬw��B�A��z^��,z�����E���I�@����U��C#�#)�l�e��,R�1���~3��p4[%C�nFCÏ��ԏi�1�|�v����G����25*8�ݑ�R��S9�}�[N�����$���kI?�Uh��P��5�G'���w4r��\lY5k���� & qn%�4�d��їcG�q9��bA-I!&�������1O�	bާ�:x�m �0�\zǉ����m�&q��O)Ű�"b{��Щ�N\o�2�A���X}��"�{JN[ ��7�%*��9�����Pm?�c\-�-J0�b�C)�hxsY.��T b8K}��Sν�Z':����U3�v�{C
?���gX���s>�2ʵ��e���L=L�U���������q[ޞ���zd��F��沃�T&�۪�U�k� UԒ���Q��>�l��J��*r���C��^�����@���OdP)�Ԛc���F�m�`�A�s��.~�T��C�ج����ͷ Z�L�u��`�����P/��M���2�n�I�e)�jk_9��
1������-)�{�Ueo��2��jP����Y.z�_�m�PgH����g�}ՋD�&���?�{�EOL-Np�U�^����'�eP�]�O��d�9��w�N�@=ZQfk���?@��ִ�<�����n</m@��T0����{uE�����1G	���O��<ng0gT��gm[�^ԯ�����l���z�ߥsZ�W"�0>cFL�v��>�,S�va����D����-��{������:1�؃l���	@���*�#�:�s!k&g�~sQC@�����T��}��Dw����$=���\��E@<�������:�/DJ��
?C�K�G�	�t3a�r�}c�����)_z�ׁ:�����g�C͞��p��9���$ܝi���$��ެ'mS@���l/HБ��N?B<b�}~Nc����(�o�ݐh)�.���1[�Z�AX��������?�{�j>P����w3�I���sAij*I�j�q�Բ�u�~��F$�(��_nN��;f�E $��1���Zj������g4$8�CV��0d]|�mʠ�My[����l�l#�I#M�0?Q-�j,Go1�����I�Cm�Ƌ���_���Q�����1��?��=�n����4CB�rL}�5uB{7pRaY\Y%>�x7�:�4;$<Ֆe&�#�a����ɼ�-���DT1[�]��D�n򿴇��2%�t�j���l�0
:SS��
)p���%���NU%���`4Z���!����j�	r�jM���~2N\�-��ۻe�&~d^�X���[:h��d��FNec��/�p2�z�\��4�pT�rZiB=��k��7|N�ZaZУ��κy1ġ�^��R�u�8D�PK�~#&�f{Sml�$�b��"z��uQ�k�``ة@.aNE4�z̿�88��Л�Ma
L�!����kP�\|�oa65`���͜�yJ��\͝��g��ۈHC�{�z���^����b���� �B�.�T�A�b�@d�"�::M��a���j��\I�xW׫0=�g�X�M�_��I��2������H��\��  	�C&D�t�j]Z�Op����_Pk�����ν��	��(2���Xw��P�!U�P+Q7,;2�u����!�my_��3�	�v�+�^Q
�$V�V�Y(������� ����&5 ��k�
L�W�R�!�@����I��υ���e������%���狂X�5Z��a�ɵu���]�Ap�',����dD��93�Cjp��/��)��[�E��n�\�!m��X�5cb�/�i#/-W{��Z/c!� ��n��۩$���K8�)��L����#�k��������#�,˒�ݡ\dˈ�^�QGI�Ca4��/�I9NY1]���`C�.���˜��_TRN
+�V�U�Ip9���J��'���O4�qNO���Uϕ�鈯���
z��z������q�e�郜~#�=Ȇ����3[�A~�Zx<@.?j�t�b*��_�يG��6~�Г0����4��O/6�珰�CK���M[��'ŨϞ�C%V�W�¢��s�6�9�֛ 1�Љ�\�y��]�݃)m˿-�^+�<�e7#���`@�T�W�kؑ���`�u�C�ye.�yB�j�|�͛^
� !t�.���)K~d�W����-����Z�b������s �������H����}g��g�է�W(��2&9'V`5�8(��a3����ֲ�e+�J����p���C���Ő�#��9���v#t;�*b�A�\���'G�2ѫ�̆���G�o5���8uO����k�!~�\B+���r�.���!e��u�8�R�A�m���&iڑ�(�a��E�<�
`2JS�wJ'O��[�X9wV&�s5����]ٟ��n1-y�����O�����9Z\G�(�@�2����0�Y<vFl�ay>D=�q8Kom��q !	n����O��x����~��
�����i�p����/�82��T�����-�w�A5�[�7��^�+<�����|�}݌{~��Ym�7Ը��;�=���5*�#E�Z�-['�8n,�Q����=�F{&eb�{&z*h�JugV-/��My���[���j1��Ɋ���`f罓W�{ �k�
`b�\���8j
��0M&\���-:��R���칏_��{�_sش�@�
��zsAMv~PGx>��o&�l�j	ߕnm��A���?�߉���qɐr ��b�l�������Q#Y���(�]mDw~�JH뒷�6/�+�d��=nf��ɴ�'�h�z �9��>]~����a��n��N����i����]a���$^w=A��|*z<�̖����R;���c�N���\��6	�	������ف�QQpD$`12���Q�1	M�fqH����H�X	&�)�v��ca�8��"���Q#�t�=ߜ�K��г�����{���Oz�v��h�߮ۊ�l��	���6���<I�9�Ň.M6Ԅ,��5<��E3Dxy
|-�>T ��0����~��&�W�VA��	��L�n�8Tȩ�g��{~ë��9��d��e�
~��Up`(��֠?��p@y<�{%�(D�N�o���w*��GVтP�I�Q�f%��q�ʶO�	��֐�5�]�oX&r�4��[�ƫuM�u��OúT^"ާ�C7^mi���'�E}p����n�4�R[�BE��w~бl�l���AGn�|bsl��s�z��"�����?Eeܨ:����C���C7K[c��*�Ncyf{���)yx���HZ��i��/89q�q���J@ҁ$����"t��ԝ"�d<��x�F���x9΋��qh5Bt���)�"(�A�}(�m�𝸈�5�w�!U�I	�G�Q�w��[���?,��K�օ�!l�������':.��ؘ<h̴��q������͏)���(}�Kt_O���Z��?4��)nT#�2S�|k�VOG�K�:7/ۘYM���ƭ��-ɳ�y�����[b�}>f�i�Ƕ|�S���Y�zTG�m�%by�/��_>��DQ�7:�)�7�����!�G ݢ���yyk�/2a��J������J磬oET��
�3h��cP�ߘ9�X�1Т�r�:�E�2�nS)�=ثa}[��솆o��3��cc����0
�z�:�"D�X���_Ǥ�6P�Q�q(���&��ۮ� ��4���c�}��b��3���!�������L\�ӹ�^��e/��(��6{~`
��&�Tn5m�-l=�W�2�v��o	��9�r	Qg�
f��Lr7����W�=u�y��{�	��h��A?r�ݧL?�I�}����4�0Z�<�	���ʪW�F�Ӎ���M�;}�~����îA�+��	o/����T�@P��J:��D��ٿ���6�	���kC�q���
��&����	�oZ=ORQ0�Ɋ$��8ߙ�q�ʤǼ��Z�a��",�-�8&�\���ӷ�[չ ��E{A��֬��Lrg�-^��[�~��V8A7�A3�jN��r���fx��kXXX�B
������E�+V"<ܸ���B4�,���{�.}�5�
�j �������䑮�Cz�"���wL�ۢ �7&bЪ�\�dS�ӷam�ܓ��;йdT��u+�3� �0�r�����eĲ��f-u/v�{���M�>�ª3ok��<���HUt�D�k5��e!J�O�9K�N3�T�;���0�5�vG�cs����Ih�!���_~�l�C�}Ou�=ܚ0hz����j�絎���'���R���l������*���9B������Z�z~Q��njRc�`���֒ �?׋�\��:�>?,5�;F��,�Jm���*[\�i��=��QN������ RLyl��4v]c<������gc��+��ʧ��{z�����h0��}�~#?2���c����>-)����B�1!��?H���9�D���@�f�^�j�`��!�@o��a����l�e~��a�\����T�h@.�3U5I�D6�۷���AG����S Єj��=ߛ3�l�iP/~���$=�sL�����S�]�lr
� E��jz�y�����?%��ZO�ǝr�E�\�d"9�C�X�G�ߑr�r�����	�*j���JN$�����olS�a��E}���9'�&Ď~|�#��b6Z��n�cF��C���z�����Uwa�ۛ��e�r=QH���j��W�����4��]�@����MA��_�Dy�<�W*l�u$�c����`�e��2 �q��^���W�o�N�Ozw{���Ph�e���fo��څk�6�0.��}B�zR&p��3v�
�9��ԯ}?ڦ��?��� 
� ��+WV��G��,�ɍ��a!\�}G>����͉�f���]�S��
�������/���_?u}K�x7q���v Z��5��<$�������g<1a֭��R������"�j�?ɚV�`.�]!�������S�\��`pa^����:�g�c�_��U_���o� ��Cޱ ~�ߛd�ĉ&h�f�}�:+�*M
:Ο+����Φ���h��_�����pD�P�毾��5v�r����鱠��J��ߵ�y�%S`�^V�Sq����W�z�z&�#��N��Kp��R�{��^�-�OP��w�HK����, :ݭ�`mjrrr��#t���f�!ɠ�7V�cgr����c돧VlPGhqUu���tU�p^/�\�^�3�$Y���}Kq�5��#��_��D��t����>G�CF��m�Z�1��wyI��#����[�y�M&YC�*�9���sAg�;J�FIm�.2���w���.5�+"!��佻���(��n�V}�=*�b�/+X@�0t��Ȏ��RY���Т{�!,�p�,b#S_�yN(�~A"����U�2��Ob�����_(	;�8��ٍ�6���XA
3�:1����*n��s��iO8M`gA��#��C�?:��� �x�~������^^w��1S��_~���b���Y3�r���oqOP�]㽝8Kl8�:!>�?����~�����.9�VK��Z�Ml"	��t�j�m���;���{�/j�]���Ё��G{�2߷��}
�T���[��3R
Z�CB���L�bb�xʞ��R����$��R�v,��Dp�1�Yla�����z���L����0�̵BԂ��S	�O���}��������W^�p��Ps�p�Qvb[-\-��"�VWo�uZ�G�Q�P��?�0�S	����Qc	tכ|�Xr�bU������r?X�@!l$,!N�9�)��]{�>��C��1ߚ36K�u�=���E̻����5��>���c!^�4�ur�4m'�����+�ǡ`S��O������%��0q��ʑ&{���S7�#���~��cM�i�	FH��^&&H?Ө�n�̸�为�۪P�9|_�榋h�ݢ��侔�D�ݠ������Lv{v~��EV�4,in������,(t���`}~��v�Kɏ�Qk]�F-�lAp�c���RL=��	R�{�9ưԲs��P��S�M�_Gi�M��M���t����܈�:�t;���im�[�i���w.b�U�����]�R}���]z�/�6�/X�].Xf}4��e�af$-�"�����z�*71�!��^2�wW��li:��|;�Re|%Mp2�C�wiu1���&�z�_�����l.%{.uUEN����"�^�{*���Y$���cG�7��fP�~� u��ca�+���ul�:ht�������^]�(�[2j�-���OePF�A���)�1O�/�Ku�_���&��VM�8kȑV>�����iXS���` U�ПF����n��ͮl:���R��w�s0��)���b�o3>e4)�O�N�Y�b�{-�}�\�>�+:"�}���VK�����k�%����g��ü���$��E�ݨ�/6��u�t˲e@�ɼ��r�a5�=�Ė�&NNP�}�KТZ�5;��:�������n�?1}��{Le~���!׋dܴ34�H�qc���B�3�1!Cb2����ڥg��\-5��^�}�tLgq'}�кgk�f��F�\��s�����>A��1�D
�K�������i�ʀ�8SB�O_�f��O�1֩v6�����/P������鲽(͏�������2��<e~�����5�f����dzw �I�����Sm�^+���;��v��x�|�z�(Zr�x+����E��������p�蜺���哑�EJf���Q]p���F9���r#�?'��Y���B6q �ʄ\l+j���p� �69��^����8�xө��T%�T
"��Hz砥L|Ѩi��k�,x���a�P�D�T<D4�p�#ғ�u�|��mM|�yT݄�a�i��#&�v�T���l�����\td���'��`���G�~�_#�����3���Y�0y����	�-����Xp�p���v}�Ws��&�0vk^v�:�5����CK"}d���w)�����Ҳ�3H�U�g�������� �)+V��t�U5�l+�H�P�	1R*�Ex�2���C��<��G��'R�>x�8*�XD8/U�A�q�޹9�Rp�~����/4�T�to�Ϻ`�IM9	��p\#�-���P�J}�ϯ\[#��o.�Ǔ[B�]���J2�-8yX������rV�e:�*�$�=�[��)����5��ݼX��Qls��;���-'?�V��I���"!m�V�ک�g^)�)Ⱥ0ͫ�� ����u��@1�}�&������[��67U����`S��q���f���H�$���'���R�ik@�����yϑ�������6cc�F���X���O6�����UW���C.��ǉ��HǄ ������F2�D"+�&S��q��0hP���bfP��
�п7�{��[�#sN��G��� ���2���^�k-�-�N�8�C�v���zx�?.�S�$~@˶k�1i�ҔG�j?��?�$��/�q��a~77)2� A?'�X��XwE��m�+��J�'����ԗZ��plr�#��*DȷV��hw/��y��E�B�o�
{�ma6��B~9�<ò ��BJNTC�	x��%���ok3�]<�N{:f1��Z���m�ٍ��r�]���Ҭ�8�}=� ͱ��-D:;,�Cޮ�?	�yƴȞ�x���vZpK�;�BY�j^!۽l'Z�Z@-�F�<+|��qD�1���_��m��Cd�zq��_�������G	Ë�𤆇�[k��^��A�P��y��c��zK�*�,׸#3��{N��6qga_��͌��ϴ2�!ի2�A���M����2
Gke�3�TnޘtE�(G�o��o���w;�WP���<bE�1��[|��΅���=L~��:t{w�*�_�{~��*!?0U�͊�,ox�݂�{Yb��mfi�@�U�c��1�� b�~�d�N�����0�� �|u3��E�.u1�<�e�[y3P�+��z����̬��7��r�S�j%�n�d������p����T��9o����A����d�1�y�K��f<Oi+x�kjC,})`ۧ��5�ݩ��@��w��X�3����`t�Q�uIf���)���B�o!M�D��1s��w�|���׮��eP� #K<;'��Aa&Rf��M娱*��paM�PC=�=#��u�gt�+Vj	
�P/�yE��ֶR1� ��0�.���ƕfm��C�V���� �hw����0�� ���B*�=M��D�uxE:b��"(x��_h�#(���b�}���o�C�+�"v.�Y��'�5�^|�8e��j?�f^��h��V��]9�@&+�n��㡾�6�wn�G݃���D�¼��g�q̙T�d�b��|�T�fYV& �I�kZ�������'@i�o�"�XO�����?����L��uߑ(=�G����v�dVB=��076E���$����5]�I)=jUa�Fzp���b���ON"?�'r�����^鞩�=ܭ,��ic	y�$��ȃ*u/5b��#��(���Y�I�F����}�����P�o����R�9��A�V	dFA�4m�:���Մ�J��%fI{�l��˂2Mĳ�~��h	�^*�����g�ð��hx-�^�2�؊u��{���V:W{w<�#�;��1+kl�ڼ��(�^��	A�\g���Lu�w�"�q�R�NZ���u\�?ޟ�N�m:b H�^�l���h+��=;zezī��4�?۳˸�ˊ]��\p��+L7D�uGe��}�n-�;�X�r���;s�kr�̾�.a忨ILx�U��]��r�zFې����K&�Hs�*�sÖ$���M��U�9ч��ڄI}1V=\�oo�r)ne�8B��z��)H4�!8��!��k�\�]��$���(��Ց��BQW۹�ȲD�u����_A�3_�+��vې`(�9�z�t��nՏk/���7^]E��<kS���ܙ�p2��.���=���ߥ
��NCT�c����iD���߆l�_d�':����Bܺ�t�6F�&�EG�80����w�B���D�}�����H��)�z0T�= ���RLl��h�i"$�g� ���}ᩅ -Q�1��<�	qtK��G�J�U��EDZW	эiɁ��P2��Z	b�>H�� j��5�נ�~3��>�V�NE_�"l�>�9H1c�|�h�嚹J�pì����`�ʊǪ���U��*&X�3���Lը�Vw���M�[�}�84r���Ȅ�	��,�z#3ԎEZ�0�	�1LdYП���X�P��0����r4��X%4 ���O:�\̊�p���Y�J�M2e���uD���G�ϾnL��/�,���尺�G��n-���*2�W,��Lr%�� ��R��k�Q�y�ع�'��G����vڄ���*����wj�U!���QW����?��54�,���o'��O�-V#m���I�����ڞ�%g��(a���8��],�N>����t�S�Np�}~�?��Iz=Lh��11{�{��#��x�(����Z�)[[[NC��N��H��h1?����[ o����AR�5�p����~j)�R�����}q0V@Ea!�5���o��h=X�n2Z��xEH����*�I��ps/G݉-b��;��,;��0?�ə%���Oz�c.A�u��?>�p�o0�Qb]_*��są��u�Y���~4[�<L���"3��O���k�x��/�~B^Ǚ
�rp�F��e�U�~`�����%?��n/�Ш�'D��0����48PK1�,Q�':z4`�� �h�Y����Ny�7D�$�#�9�q�,(�g���b�dJW��$�sEY�)3M!B����Ӻ=�T�����΋J��/Ow66���a���<?8��~c��K�I|"���3�y�6"�Gm�N����H-i��'����!� w�[a��[C�<���l�r ^P��ףjVm�ߍ4�[踘�a٧������ׯ~�Sxd���Sk~d�K^�E\��1b_"^_�sd�/2��0�L�1T�Ө�o�����@�z���~S9���� vrwƏ<v��S`�N3�u32Ǹ�]4l�1��<秓?�^6Õ��M��7��Y��u�K�~�yy|��1�.�b���atF�4�rg8-�z�U�����pBC����cM�����s���9L�����L�����0>�d�B��}v�sP.���Yٓ��嘂+R��P0/GrD�6,��3jL<:_BB*4��rE�Oɹ:�?��̙dcv�s^�uK�,�`B����l�1��r�3mO5Y:���#��o0��u;�㿃��aJ]�6Em��e\��Ĝ@wbN�1��b8!�c��-�֌X?m�1��~9��w9�4M�Q�@D�m�\Χ�F��˴]��;����Ke��}�9y_��6br��3��$n6<w��jl2�Kh�c+U�}mj�8/�����ֿ�ey2i�4��1�)U��9�6�G�0d<If#�8��<�6���a\c�؜�v���k�p� kb�NE��`��f㏭��$!=�x���DO��͋/��o�:jj����KP��J��Y'
�=t�(󷔰��D������h���s9��U^���E��ow���r/�o��H91CH�=L�%�i��eR(ͬ��^��ƽ;��[�\�E=�%�-��^�u(b݄^��k�ح#�|a���gz3��Fω�
�{�I�G��B�ǼIl�{��v��
S�D�X�c���I��$$[�ow;���J/�T�R�!X�!�_���g-�b��ޗ��	��t�)��7A�����D�֪{�ٺ������,b�ǟ��#ʎ7��FxֻA�Ș7`�Ғ����Eђo�֚1�.��������:�	��9$�����ߩ�L�b׭���'�ML�6���v�!~��u
F���-��lb 8�L��u��A��E��_�)�0���/,�����}p�{A�[5m~N۹�y���?���h�s��]MH��Դo��޵U��,y���l�YLY��%Y퉳�n�^��&��D��i���B�
b��(���$�Wz���俻�ޤ$��˂"Nާ�]1��cF'��� �(�j1g_��l'Uf�-���!�L:��0�ޚh<`G�/O�T�њc�`\��F��J�;�����(�S�����%N>�]zwC������F� k��I��X���QJ���4?�j��D�L<Ċ��p��- ���I�E�Kt-|1̇�������oS��3S8�I����(��ޫF�w�T���|߅&6��<Ԑ�����9e �z�Pq�s촮e�p�z�R	zp:p l�G����ѵ�C��O=wD���~`g�XI���ʾ2�Ļ�+����!�����ݧ�]O)�p4/�4�4bS�_���dY��Q:5&rXy��P�3�nPi�="��\%-���?0��|�J%'�W�%yTX����v�kp��;R\!�V� ͞��OO3�`*����>W]��nkP|��к� ��O��f!����U�v�ѻ2���^7�
���y;Y�e���o��nr*��P `��
���J_ܫF(��Q]��A�?(���᫙�?f�Msd̢W��-0���}��f*t��*Q�����Q���������̇��Y����sy��ݩ�W���܊6
�D�'r�K�A�"��o�ɿ��D�^��n@��Ӭ*_r�6X�OXر0��Gc��7,�b�ڥK~��O~�U`u�ٳg���K/m}��k�˶�p�[8֪7fG/�4�����U�fDO1�� ��MR�nSҧt��K�]�9ܵ�=�O�sq�"Ȁ��L���٬�'UT��/��0���R�8�s�������`S���w�uȅh�0(IN�X�>��K�Db^b����D�h/�`L���%�Ç.�b��|BpE�_;J�ϝ7*�MΧ��s���4jN�1�q�+�2}��G6�}���L��ʎ� ��������>Gp0����%E���O�g�" �\�(a�0��Fa��H��/i��8�c%!�E�b�`�^�)کI��b��pOp7$���1��C p���G$1Z���H�s��b�_LH*;�ѵ(����dC5ۘf�
f${1ܳ�a>��g�ɩI�{@\��D����G33Ӯ�����W�7������?��:,����i���Y�d�u.�r�ɱƮ��'����hb f�"��H\Ra��~����7� G8a?�v8�:d[W%]���HJ H� ��y�y���ꮮ!�r�<��[{������%(L��F�+�L{8{�ok}K8+�W�#�ΰX�K� �����_@�؉�M��&64���W"b++��8}'���KY�\�f��&��<�bSy�<W!��`p�,+�ų�y��-��|��/t��~����+宩���S�Ee�B�/t��9|��D�Mҵc��3̗gGuLe�Ƿax�`�*�S���r�چ�� �Z,�D6�����ѳ���1�x��Xal\�xQbKO�8��G��o��[|�Nn��eX~-�\��K��K��|�\��n����/G?�ɏd��.�}7��I��U����uw���ح�Fv�p㷕��Z���$��*�%��������{�_ޱs��C�]cc�c>���:�&6�j���g�|�ͯ0�*��̘cǏ���(5����T�����O'	�SE��j�'��X�n0j�k��J��C6t��~��dx�e�T�������`�8���	��R�0�p�,0�����<"&.i0đSii�9s�q+S�<��X=�ϋ���I[⚚�
���F�.�ߏ�ݑ�1&���{����q�C�β�3�3k�Żۄ��.�"4"}��;�b���4 :hX�?�]�����Z`�p�|��I18t���r.�ʒ��P|�L@�eF �s��ɸ����xF�$�,-/ycY�b�✓|�o�S�`'2ज़���m�͜�+(�v������-`��q��� $.�I���
� \�$��!]�\a ��ݰ1}@ ��$����}������O�*���ss����J��W*S'N62l�� �xBf$<f��dЖJt�m� ^��:H�c��E�#Ж�AmT�b�H��P`��}C��l�u̇�����ӗD�!0�wI߭�H}�c�ԥ����*�)�.J��,W�@�`*�8(TS�>����Q���g�0\�v1S�<2����g�|�W�RGd�%�~�n?��:aT�FS���Ǉ�\��ȫ�J%w#r�-,,,�Z���cǾ�s˛|���X˰�ڔ!��'������k'N���,,ܢ?��n-�n�Nꐷ�H�D���q^B؋56.A"�-F�(�U����t;�t���U5#��h�R��C���G}����`���G�'>���������]�v?�i��G���M��V_�m�\/e�4���ϊU�E 8c��#1���d���V5��w��gQd�?�pBՑ
Y7�Dܷ�M(vE�F�Ir-��������dݥ���%�٬+���0��4�o�kM��(p���rY��+�b�I>\)cp���X��(�? �;�jЩ��W��Xdc��⌔OttŻ*�.:(xv(	�G<;�C|����{���h0sh#0� � S8���*M�y�p�z��ZP�����sq[1��4���j�l' �p��C��"ڛ�+ʞ���M�qTV)2�z�3l����]۹�Lc�$�ʺ��{m�h�����>I��p&���4|<h��A< 5��vp��Ks�.���Cw���B��SOɦ��Y�r劜�y)G^O�I8 �贊�Y���@M1Mw[�U6)uL�"�c-;.C�[��\z�6�w�un�ʴ��	/Rq��K�]}��@LE�X�Pp�/e�g믬��g�A ă�d�!�X
���U��*��1����	�v ���a�e�^'՞W�u�M�p�[�ϳ�������C��'ܤR���
����?Ơ����{�^<~���=33�����װ˰���!���
6�Z�%a�!7M���c~e&; ��Wn�4q;xb0zE1ͮ����7�`4:4�L��.]`#ݭ��:{��7�߹s�{|��={�����\k����.\�p��a��ɓ�䬰a�LG?��9-�&�U��]�uM���b��!4!�ƹ��0ڱ�i�l�VitO�jٮ�,�vW1Q%�i&r\�����Ɔs���F��!ˎ~�V+|��0 P}���K������z
`��8Ǳ(�bt ��nWT*�����
j4�|V��kцn@�v����V)ѹ�x�J�Qe����#e^� ���YH��N��Q�O�,'|! ǡ��l�"�����Q�ur��R'��ߖ~N�Pd�q<�ڱc���8�,X�b�s��\|Vl��d�3n҈(�����X2�l7��~���ͫo7�7�lRb%�$���ny�E��Q�:�V��c�k���Y�җ^���~Z�)�_��sg�H�����l��cI2i�4GDw���ɲB�V!�NpA���( �q���l8���s��I����:�\�LN.wǔ)V8`�d�#�e����P�D����߷l݂gL�!f@��9�^�F R�����Ҿ�k6�������H��S�� �lR����߾�!��>c0ֹ�*��x[���K�]� Qp��"�+E������e��^�ï�հ˯_��_����~�V���_/�~��#D��8�xY(�>���pQ�B	7	X�k�;U`��u@���-��C p0�Tl��}�6X,:�zü��[w�˥����ŃG��_f�D�7��r����������o}kF2�'&&�V�mj�5a�"���g��v��_]|��D��(��}�&�a��4��QfIwSeW��[T�:V@ ���5�V1�2`�&&6�G9Q�S�uA�L�Z\.U|L�U&,��G� �����=�,� Ȅ�@���7��t��HX T(ۢ�΍���Pœ^��+���
�f���vX3��>	���W�//e:%Ƅ~����`�<+���o�'���$��8p���	NH�#�� ���j�*K�{����: ��g��O]3�9ѧ�9�����z���P���V�ʡ�����0d�dΐ�iS��G���CA�=�c��$�QI�	�E�wz]��7����c��}�D�q��"Z�iS�ӄ�%�1���W�J��_������1�)V����̈́R����;SD�OaA7[��w#\�� �IQ��[d�Rʓ���+�}���YDK*������9�:%���K���.� �<Ϊk�W̦�p�Ǝ)3YV��ӧ���C���3�� H��>����µ�C��߇�S����yb[���Ǉ��\��:bv|�'�7o0��sl��:�G�3��a��f������, �Gm7��y;��T�<��]�v}���K||��eX��׮�կX���v���o/_>o,;�w��%	"����~�X#l��",�3�q$n�\Ï�!n[���={�{���F��t!��K����x]��ܘ�E?��/v_�:�Ԟ�{.=���?>{��<!w�%;\���liee�<�f|;,���Ď����Ps�Ƴ�6������[�km^�����<|�o�����m�U�C�"y�-�;Tɍp;U��!j��:���D�@�#l�����҇�rNI~�.�K���f�a]��\��o�R�",��.%]��I<���`e#(bp����}q���Cn3ax)gc4�v.[`�Z�	1u+�e�3�C�]�Ɇw��فx��Ms���t���w`��G�X_�0�aT+�c�l��`�Ľ����`�Dv{+���:n���
�a,6��K�-)�>4���n2>S�X*��>�%�R��&|Vf?��26xg ��9 +G� ��W���F+�3<b�T��I�_'�w�_utDD@ ��wuie��o�(�r����䎎X�K@�^�el��?_A�������O�a_��h"�3�+@�M��49D�\�r� j�ؐ�lk[�������:�y��pI?wT�+�Mo5h��*b0�Q�Ռ����T�֩�s�Z�N�N�Fx����^�ʗi�=Ү`V���ťY�+"��h�A���1a̋"r�c�ܰI�1V�q虍��K�Ѐ	�XS�_�sa���X�ĺ!����ׁ��f�B�<y����HF?�@ *��<CW4�YC������Ź ,��`r]F���
���^
�:��_%��ZZ�����v!��>Up��j���S���T(�ꅐa�R��"*�q6���k��p*�tm��m��4��B���L<��?�[����ϣ��ς��/��9�ʕ+x����ww���
��H���i:,��b��_��:��Y][)��Ƌ]p#=���;v� \��1� &'�7:�l'oc'd�{�B�]b5�P��R׳p�"�7ĭ�7o.�<p���c˵���˕�O>�]�A����󑛳�����~6Ɠ}{�.�9����ȖE��_����6-..��?���?y�%�ͭ���	��Hk�A$c�]ۏR�Q1���L������,�U�%�'yjG���02I�FL!f��4��1V�[W���0��&��N۪�(��EM���`	@����Q��"�8�"�q����b����h��J�j&7M���e\̎��9�7�j���o�>ڱs�A�݅��Xa�B J Y:V�Fi���@�_��"9�*e+���s^�#p�qc˻��ë1��O.�+Psb\�F�����jeԝ	�_�E�J�+�R6W�E�X. '�+���رC�"�#d�5��0T0����� ��c���&�Y��� M.�¹�օL?�7�0' " ? j0��D56[�%ڑ�רci �@$�� 6j`�o�a�)��J�[�F"D�M �!o��q��3����k��c�ז������So�.ܑ�f��2�g�[&��g���}�s�?�E:���S�8I�L�G���(�GN�6Y�D�f���YvEu����x P���s�Q�2|3.f�q?P�L3+j���c������J%��!��_��:��Ի�ʬ+�
�
XA�A�X�^������Yڦ������������gx=r��ZW�پ�G���g�\_�s8��X]�C7̠-L���7j����>�F)�*�V Tn�ƋX��Uwt�瘛��ޥK�"�!�:u��g��9�#�W��eX��׶�կVx��a���t��/ɯdD	��:Q�]M���˕L����v�Iw��$yn�T8Frb��pIl�(D�Ԭܢ��0��}0r�i�kݼy˼��ϰ�]߳gr`}HV����`�9����m/���7�x����_�ǆ�Ι��t����O��G�͵�Qy���ʯܨIRbhv|i��W����ۛ������2�Ab���x�{/���z��O>S��{-���k+�&��L\0e*S�R�FO��5^���WdUGGM������0@�D+*]�*������mݺU����^ %0�+��l�Bh@��%r�x(Q��V˪A5������-[i�Νf��D��D�ʿ�p��9���ׯ��:�& -$�����#�/��\y��q@`��m���� ���̮��Ր�|)������Z��Lq*��A(��;���u���c <Ѓ]^=c�G�����\9X�x�m	? -6��}W��v��~���m��W5JKЎ�gxőN��i���pC����.`�gP�D���ȑ�����&���!H���Hl�6�A�h*P�[�J�0z�h��9����]f
���Jm�Z�B����l0�b@��u�<;���9�~���O䲺���e�_�zU��(Ί��ƌSL�W7nE����M�^��a��u��Ƈ	��JZ�؂����:9�l��s���ڝꆆ�)H��MU�Y�L^�\>uu�Mm���bǌx6'|'�o����oD`Ez����=ս-p�[�����㳮z��:�hll L}��tΪT���� �ɻ6fv���
f\�@��z�_0����gx�����S�/tG�Y�
�� ��89�K��=�-�\?~�����{���*S�a�a��.Cp����'���f�g�'�r�z�UOrO�� aL~ �,stn���,��tU�A�	Vh̍��*��N�=$ �jbꪂ�x���>������������ݷz�=����V�ܹs���ޗ_{��u��g.�;//-��M�47;_�x�.?�@�3�N];xp����ܯ�"�����XX���ß�����5n����?jU����w��r���K�T_��⛍�t8y�6�w�7�[+�r�)�SQܧz�I�^����e6�I������LT��V41��dcY��R��6M���	6�k�y�j�Q
I��P�̀�#�\B���(�ඖØ���3K���Ģ���g�3�E^�V��QW���M��W�B̠� Q�j0�U NM��C^����`��z�b��J�o�ٺ�]u��s9<�n���S�I��̯�$�X'�uv1Mƹ
j`a�Pw0{��PY'��Z��
}�
���)�� ��`�A���Q�~B�%�2��G=�=D0ԥ�2�F�#��ñ�w��ߣ����g��,x�ZC�g]��!���X�����<z�6�!`4�ōM�}�S�nSd /Qqg똄��	(�+��?�y�^��6��_����W��K�Cv��͛F]ﲌ���]��� z�Up������,dJ���cR7�9c��2f��
�9
7L����@� ���M��-R%�B��\L �kn�^�:����z��B��6'��	7Te/����0^�=���I�g!ç̗~�,�������õL����LgJZ=���X!PE�+��Qw�jOmk�g�Oa����8wI3m��8�뿫�S�)0���36Ѯ^��9r�Ȼ�<���X���iX�eX~��\�������h�_���oJ�������6b��m�O�[H�nt�ԻN�"
%c����"鍢�%�f�Z8M\���9 ��.n�R�4��W��v���W^}vl�<����__�|��={��|��s��陟��'�}�W�{�w�ܺ�'�\<2��4[��Gg�Es��4;7����c���h��}����.����*����kϽ����{�rW��{�KtσǢ��B�o�D�?A�htu!^}�U�fw����C�?ah�.�ҿ/�VM�:Җ%��5_b����i��VAܯrX��?>v!J#ql|��V$���y��ĹgE���a+����%0��$~fu��r�F�����"��r�2ŉ<�A_�X�]�?�Z!ѿ]и��;w
�0�c''7����^�N�\$�p�g07o��cN�6W�s�H��CÈ>�A����F4pO3�{��q��a��/v�I󊉰�N���mf�)� 1���@
�����m'�Ʃ	
���-�C��+�������כ��c�p����> ��NcD�I@bj|?2R�v�ʂ;���6�ai��D%���=p�����$ ��ba[%�W�$,l qO�`(��0��	\_��m2"���`����B1����j�������*5�Y�����~�b6����l�?:��0~d������H�O~�,A���b�(`1��U`�!���,���YG@LD�F��Ơ�gh��c�0FT�ӱZ'{�q)*���&��4`f���1wh���0���v0i9�PY0վṹ�ۢ2h� _�:Q�5us���s�ald�1�r�����I2�!0S��V�ȵ����Ǡ߄
���?}V�>{7f]�݆�O`����d�ؕ�\�|��{��+����x��s��X˰���!��
.�۶m��C�N|��G��~�镕Z�=�5��06�s#Н�XD��A�O�㩻�9Q� ɄK%��Je��Hu,E��dB�d��+�V��c�0z�o>��4�?{�La���s�ĉw�0Y����#V�^z�GO��?}��������hb|S�Ղ���Co��v������+2q��{�G�Ƶ;1XXUy��v�ʥ����<���o�?~��ⱓPa�&j���i�.��׿N[��W��t���ͦ�[���t��F�r�v?�mݾ�\-��v�0V�"�^����]�l4L)�S���P��_�'�X�AV6&%��N$�[QԻ�&6��}�8��vt�J��[�!�._���J%'���f�+��q��z��F��4X$F*��}��Ao?���P�=�scuR��xB��R�.츞�'�ĝ�v�r'����Χ����[cGG��� N�	��j��Kx0Bxf0Xp�S�-o ���*�)�:��C��x�p]��A�`���*q���%�+�*<�ŋ��?��4[���R�2B��q�Ho޼���Pm�޳Z��P�o�:���E��wײ_EoL[;�}6���|k�q��tUcS6�π��[����}���,i��Z�:�8B�$k��3�N�r����ǽǎ���3�<BVb�Оx&��p�{����b(���w�A�|�A��![�� !4������o���:��f�����[&�Vݹd�˗��Cdu9�>��T;��X����m��J�|Y��!p�2����,�ul[t�<��{�}%�B3����߲ u�z��gc�tp�^�������;;Vu��w�����9�@�s�1o`�A�֭[�j333sǏ��E������I��eX~S�\���'��իW�}�3��v�ޤ\���.\�8�	ј>D���˼���&���rI˶��`1�#�
����)�`'X}���:W%a(���_�B�stA��DH ;�&߫3~���g7o޼��i6_?u��/xr��},(��T��O_?��K���W_}��ի����30Ȣ|�W� ��=+�$pe�q��|��v���6=3�Ў�;�MMM-a�� �	����O�^������݇�|��ݏ=��ч}��/D�fs�4�kl�N�vNo�?�E�پ��n��x��fvw��?��9��Jk�%���)*͌���cJ���ea��W��.���p7�s����vD�O[2��S�o����>K%dz�"E�/q9��1� �m �b�s���h�` ����W��A|!/`�Z-��bd:݆wUC����˅eT��zb�������A	� ��6+j1�EЁ)1~.¸"�x` �3��w�|ū;���\Wޑ�RJ<5�`Hh�Lw�X݀����:�~xG����0��VO�$n
uW�t -q�c���5݉���`0+1\����㔡�����{�u�-��l�k�(�& Q��d��$E�
��܃b#RWG�I�;�،�I� ��� _�Ĳ�I�<���j�)����@�7`��t��L�b� �qji7[q��q��
�RA p$�n�5�*��C>���3�>� ~����K�
������ �G.�r��Ӂa� e0t��^�j�sl�~�����(����1�#��\�)8¸ޅ�����;��M�2�s�3+�	�|��z�ǻ��(˫�������e�h < ��?9�P㧴���A]�
|a�Z�	�9
��kl[��ʦ�s�m�K��Y���K�s������NlU6�Od���yq���G�Q#���m"�~gee��}y�رc�k׮˟_�a�߬2W���^���wGG'�b���W^;y�ҥ�++��y�
���0�&ٞ�Jǉ���HQ�8�cwF�L��͠�qV��ϲ��+)(��ɚDT-T#�ss׏��^��ڵk���8x��"��l�.�P�}���w�9�_�����8�B�����&�TD�H��0�X"��"c�u�x�⥙�����f�q�q]�sⷓq�xkNv����[�_~�G����W~Z��'�*?��g���DK��$�:�h�\�W7o���1�ON�WWkt�[ߧ{
����
]�?�F{��z�A�{z+5�D��I��64^��������S��9�B��#�*4��mC� ��f����h�v_��@F@�5��<6�;�L�^X(��U�[�<"`�T*��E�8�Y%0T��ׂq�E�����s���� ��������+¬�x^Y�"�j||B�ۺuk�w���jYR���gŘ�|a(�(�S�'�)�����W�b/������pS�L
�`t�7U�X� ���B,7��p�Q �rWaGب�#��
`��u2��d8�3/܉ʰLA�LG���`���4�Q끾�;��r(�ĸo/�[�Ȩ=8��v�,x��9���[ ��j7ɷf��؇FO���w�k�@��?E� ِ]����L��V܂kuSg �����?n���s��>��;�>S�D�]�ð�;���eY���n�V}R�W+Z!��
�\�:�V�7L�S����	�٨�g�}�����&�$������:�����e�0�c����˞���`[��w��`9�o�f��*{��;����]��+S����I�a#2,�g�}�A�ϧ��� E�;��;0c~sL�ok�ʠ���3xG�{x�@K?�|�r�s�<�w�߽{�x��Ȇ*1�2,���[���Q�.��C�Y�~�z��c�W^ye����l�,���D���
vئX��w�
\�bG����N�X#�C��6�(�F��f�X��WT6;�T	r����o�~�镕��l�߾���c���s�'�{��C�/]�Z�N�ADQ��"���Qjx�f�-lv������Lq��]�l �Q��޹�V��\�0ǆm��a����kС�j���_����?����=Z<q�����^���-S4q���Q��3S�����G��_���Je�|�Ϳ���x�Jlj?x��V����I��w7u+e��a�L#�Jv�m� ȟ��^1��'�I��Q6��"V#�J wŽ�I%�k�F)_�ǭ^KT�,���zd�	�>Ʒ�$�.~�����A�c޸�.r��e*m@sQ�l����8a#����5�?�����R 5$/��  �؜߿(W�1p���1{�Zb7F�N�2/j섮P��tn~��%cP���Dr<*�������+�� �� Mn��K�`�U^ݩ J��
�n��͛7E��ۥ�# (��g�9�V[��D�w:�
|ȫ[�V[�;�A����9�"~U�q���䴳IEI�c[F�&\��M"l\�
�dY�HƟ�"3�����Î�g���m���5ZY�I�v��6�]�� O#U��7�������b%�����s�tV�Z�A��D �\n�؄�����_�߱EΕP�H:���±�o��d�=낍��˘�F5>���'�G'�� ��T +i\��:��c���]�t�¥𹘔I
��\���:zO��k������K쮧�����Nڞn�
�����?6����8�����} z��u�&+)  W�o�h��Cf���{��k�$���ñV~�S��p�8E�0���`��9�u��ɏ����'<�3V�2,��e���%g�V��ɟn���U�T�������^�o�Q��O��iPzbe�dRvƑ��R�ֽ0'Ƴ��$�*���j�b@#"����nd0q���b��d�\;$��~��{�<�/--�ؐ5�K�љ3g�5"�0{nq`{��v�a��]�~��՛$-����{�w�Ju���K�����[�m�cG�o߹mfOou�o�m���;���g�3ѵՅ�ZP�N1W� e�hOt��t{�C��^���$Go�Wi��mf�\�-W����e|�֦��L��=4>=C�F��+M6X�Y0{���
l$��C�.(���],�[�7�ʈ\/�t�{�(�%��H�D6`A���H
��	�i6�bP!�n��6�> ^�LF�5 l\���8m���$�9��8k`�޽2�BР��v�3�;�
ҟ L��.R�k��u�	�|���8��u�Z�.��*��A�u���ǸJ��. H(����P
`6�k
��ٸ)\�1o�:�{1���NiQ���k׮]�o��"�6r�A������Ʒ)�јH�����_ܒc��)R����裨yW)��$�y��lw�Z�&��i�����1f�^��xc%�i� ɱ��j2���� \�գV�)��n�ݯK���������E������[�裏>BN+q��Ar�@�?��L	�ǆ"��S���� XA�/����y�όx
�z���� ���d]�t~Ņ���d*�ї5`0���ߤe�}���Ϥl���-(����X}��*;���M� ���c�y"�<��T�1>yxx���I��)}���'��9N��=cj�e��p,��>�<uKV;l��94��当�`sԭ[�z���s������ҿ,/�˰��X���_Pܮ�m�P�;U�����&��+.//	�a]D�q�I�ŢuҤ�n7�"Z��~g��
��D>_��$p��?��P�&�Ţu�|��6bWF��Ǻ����`�����wq��:X���l�N��}���'[h�V�?>s����\�2[�������]����E��osq�<�_1�w�?�/�r�#^�*�-�-~�N��^/�-&h�Օ�r|͘C;h��Cѩʗ�шf���8����<W3I���ҠM`v}�a�ڱ�K�{Ԧ�W���1��va�/*�]*�|\)UL�E��F,���)i0^O�e bO���5�����J`����d�A�`Dv�� A��i4VI�|p�?�v;��k�u%LpC��*�5*6�����7&(h�����*JL�y����i)�-�Ov�CI��I�W)e/��&�bB�?��sF�>��O�7�k���qZ _�K������	{��n���I>�������*{�q.�2�/v�!V12:N[�Tb��k��u�x���Q�L��P��<{6�k���o�GS�{��?c�Ց���<�D�������ɖ˷�x���K���@��ZmY�g_Z6�|��/�׿��t��i��ϻ�#�9���9���Lf~L���MH��s�8��t<�c*����A
4��L`p��]�g�CB�,4`�R��X��8O��fF�:��Q�3�W
|h�i<S��
A#\㌂.����k)`��6[��_Y6%a}(.}߄u�v��>����eA��� ��?Sڶz�l[d���Mw�����L�n��z�!�#�!�_�o߾}�ȑ#�ٹs���)�╇eX��7��էP�$���ם����d9c'Ԝ��BT��T���:���*<ქ�� ��s�?m�5�a�a7�fyٹ�t�J`�����3Xa�EbY�n�]�L��+�5
jj؟�U*�{y�³G�ue oT
["�
Kі-3��#�F�|0��{���Zu߾�[ӣ7�ou._�-�ޘ����2:w�b<���9�֞�9bLk�B[�zm�L;6ȉJ����W��@<LEy�_��gViӶM425M'��E*1Py�O��/\�=�mʝ���7�Ԉ;���Ǩ�};���8^�j��6XO-z"@^�k������;X({V� �uQ��"U������W��Dx��!�3��0��7�?���D X�J��%�՘�= �� ƼJ𣝑(����� b�t��X��Z�2/��M�&��!n�j� �$�\ϖuR���q��z��y��	ϣ�z8@���
��M�U��c�Źъ2^��&@	��W�I�� En+����$�E^*<���߳g������ݾ}[�?��[��K��eVH�ԑN <�rc�D�S�-�����'��Œl\����� >�o�8�m��nu�}��y*_vPY5���Z]�V�A�++ ܄�b7��xu�fz�$=��St��Qi�sg�"�?�u?��`J�� Lx�+؈1�_�e�cXBA���770�����J� ����;����U�g#0��ϣ���>��!�b��X��x`��#[e���f~R F�2]�c�8��:!�;��&!��F��������E�@_h	c����
T��H=?>S�����S�tc&P����&N�B�`5������G�� J�d��$iܰ˰�:�!��
��k��o/�Z�LVBU�����b*FJݕܮ����V�[&��A��_���.�� GP�7X���b}�����	���</$b	��A��x�����LX�Kl�lDġ�F�e���{�ĉ�X��+W�"��O���Tytd"��.���Q�A�L�N��1��{����}y�=�m?y���$x�咖Ș��	�:�(�7-�ݸ��Ya#�vu��Ǫ4�c3��ߥN.O���7):s�v���y���4�Fk�v?t*�n�j�.��iƅR�T$�k�ʅ2�c�c#��`�m䪂R`��;>V�f�m��P`VFL�d@3�uw/0��^M��hץ�e�ә��Q��8*��I`B�o ��1�Ӎ�B�xW,J���O8A_�.��cQW`��B]<9#AcH40]ws�A"�L	U�����M����Ԩ�A�:V5
��3�|�Rǽ�7�&�+nq�n9�b��&�6N��� K�%�=� ����]|v��u���nj\T�>���&	���OiS��`y��;j���|���m��
����H];Հ�iʔ�g�c��=�Zu$-��UB�W�)F����q��bz.����s�ԁw���<=�������haᖸ:�9�fYC=��@�(��ϝ�~L�i������>����8C�3���:V5��{�<���������)��ϝ���G��� »?pmS�Y79��"P�L1ea���^��-Ŵ�m��)%��Ӷ���@E�*[���C`�,�F�i��;��q��V��w�ʇF�X
��6-��P���s�������2J��k7I����y?�9p�{u�}������sЭ!��a��/Cp�)�~��x������;��z��V�fE��Ci/�k~�:�������.���C'o�W��@�ȱ^��ܼ<�ry�LȒ�8���.������(��&��\>gDT��������t�����[�H�z�F�&�\�յ�?�a�D\��^s�����+����o�[/�BW[��l�fS!O��=J�I��:5V���u�D��:I� wX��1�<u�I\�]4�۶Щ��<UL�>������g��kS��˴�\`7����N�������fC4g��GPW�w�����-6H�H	Uǧ61 (��jA(�ce��|_\��c�fP,bG�0��~�v��GFXe^TU�)���qP�qD�={vӮ]�;%;�k�~����� c,�3]Ɗc��sɃe8t�Z��;�+_� ���]��Ewi��]UcU�OY�9T���{\m
����������/_�@	灅30�6�x���gs�� l����8�@�8N�G�`ȣ͝Јߍn�8���i���C�wѻ�ƒH4�B%��cU��\d���E_b�d7]77����?\�E��e�6䄉�@]�:��ڿ�M�AU����)�90�f�����_z�����iы/�x�F� h����ӟ5���(�l�Frh����k��z!h���6RС�Lp�lR\�'�t���ҿ��Хl]�[}����?�\�&��ʀ�`�-���O���-��(��]ނ5�o���kz����^znȌS L�g	J����� |@��a�غ�k���0����wY�o�:�b56L{�B�*�G#�!%p��.]���y�������$��,�eX~�\}
�}��:77�ڙ���y���;7Ɋ�x$�E�	[]1�Gn�,܉���go�;W5q3J�Y%A����V����S����+ۀ{�;o���Kr�\��� ������u�Vj���7(07XN��~��Ŧ�l��vǜg�T�v)�i��=t|q����us�?��k�t��4}��&����b9�Zp�j��߈���)����\a���-��.�����أT���T�#��Lh���q�����t��'����5���kw��`(|�O��1rJ��U�C�Ӓ$���G�,Xa�?�C�$\��< v�khS9`��g⑑Q���$Ny�J�(�
�i`I��w����*��6H`POM��� 80]N���Ё"Vy����0(�[�M���%x`}��b��-�SHF�s[S Cy�0F�̨���%`��MĈ�mO��S���P/��^���[ V`� ��X����q�*��/习��h?<#�� ۃ9�����)(+�b�}�z���6)��`��^�������̰s1�n�+������x���mP�
v����	�ưc�위�z�/ک�jŭv�tX�,����V���}�Y��/�8p�Ν='qV��4!;��2�Ȳ����B����.�n��X����-my���ƒ����i3�BJ�\�+�Wx5��-)�n����X��FD�m̻�{n~Q�y	��Fu����s׽�z��n� -����;( k���z�Q$'���3�Ž?��M�' ���2�a;f��$�\X�=��X)�6%c݌rm�y!�~�://�5�<|���y�<ӥa�a��(Cp�)�[��O���tڟa��Ɗ�e�qJd��;����������Ww��-Lc:\��&mD�v�;�PD�xaaWU4����9q�`��K���q����� ��(���v�ټYγ��������R��n�/,�~�צW��.��Ç����ݸ^�o^�h�_{�޿5Gw�n��O=E[&���Ƞ�U7�?��������2S�V��5{�A�-�t��g��k�^�?�m�����>��ʵ]�k�V�o���#[Vr;�+H1��C�]�J;�p�2��00��؄Аڅ��Ȯ>�GGG4uڝxiy�Xy�]�:+}�yf3MMo#ܺ�u�:�10���ާ,�c��Ѿ [�U�Ѧ��]p��Eɿ�"����|�+����1�xw(?��P�ٍmMh�,�75���Y��� �| P��B�����>�#���@�oS����� �*#�sn��(�	�\�����pmE�ŹE�Q�,���2P ^x.��${fP�� � ����n��S1�It��3/�����T�u��s�ScU�i�`�Z햸B�^]�A ��`��]�o,s��
��1��W^����Ks��裏>�R'`a��G��RZQ2��q�FYkS�pe]r�;����ΰV&J�.���ͺ�9�E��7޳�A]U!Pz�H�?9�I�U��Q�r�\K1�!f���:/g�_ȶ�MD��f^���)Ō�`L����b؟)�w���E�]���Ϗ�sY���᳇
�DEC=O��O�ِ�
�k��68S��`��rNj�����ļ��������}����gϞ �⯛4,�2,�5e�>�r� uggG�ܽ�̹�g�n�h��Άn���r�ł˩�g�[Iuq��@�,�$�=���W*��bT��1�Ū����	�A�'^�3�#r�rJ|.~4�Fvݒn9K�5>FY+�(+�$?�=NL�ͻ���ھK
�9���rbď!��c�R�AM4��⵱ǗY�^��[���bϘ����z��?{����8mѓ�>Cwm�I�6����!*W��d�A��̵�R��[fS��J�fh�w�m��	������#֢�Z��?�-��j<u��i��x���Ta�T�Խ~���J-�+$.�&h�0&���z�:Ԧj�������߅�����$}���H�N�rK�)�tM�ݥ�/Q��Y�����lȏ�;!�],�Xha���UF�%�%; 5j�����ݧf�cZ�.�L��I9gn/.���"!�g�A�H�l�墕������(����a�0#���c���t���'�{�['�.����jy(�N��1�2�!��̊0Z�O3u-���惂%����� < ]8mf��I\`�7�@��i�[o�A�;�m"7����X�7w�"�m�|i�� �"�ɉIUȾ$��3�UԪ�nN$I�o,d�#I��"^~a�z��H�Y�C������c~n�@j��A��p�[��Da�eW�#.��k�gC�׌ۭ�H�7�Mȭ�������Ϝ�Z�Fo��6\i�:!���Je~Jϊ�\Cu��yV�B���&��/;���,#�� �:`N����8��q_5���Jn��]��D���y�UMp��H}5-����(�[�B|��J.�ɼx~�<yP��u�z�� L9|ς:����}i �D�3�0�f�4Mx�B�p=V����;m�@%,8����#)�e��Hl�y�Y.g�~;?X7�`s'��H���r:�\Qڹ Q���yF�Xǟ�#U >:~ \ǜj[*K��#T0��D[� ϝot��(��<�s`��Yl�9r�։'���7i�8,��[W���S(n����go���^�p�����
�0� T���ȫ���l�Xr�xW@Y�X\�Đ�lUK��]iT��J�&G�0����ڋQa��n�W��{�ĥj���4���43��c;q�8��@�F��ŀ��^����b�9.101�7o2�v�z�v�2R5��-�:;�)>�~y�����-,ƿ�M�W��f���yƍ�J�Z�&���-��_���:?��T��I;�>@O|�Ezu���o��l0����O_3�W�΅E���x˖]�����q{M�Ż��V6j+04���-\*Bt���	c%�U���*?���j�Q%ܺ	���q b
H><�lc�4	c�`�
RĞ�A;��х�l|l�$����}��] ���\���Qb�-�ȳ�a��m�O(�~H��~W[uOØ��?����e��Z�X' JeNQo\��
�47$�����N��ST�^�g�X/H����vˬ���TwJލ��i������x5X�y���~U�����^@ n�����X߿���جG3)�ML,̯e��TR��x��&�V��r�A���!���_�e�M�� )�������j5��wO>��y��رc4w}N�� @Ѷᆌ�R����P|!�i�r)`��mH��]

p~00q��{�5n�%�m�L������w�@(٘���O�_r ��5/I�{>V1�H��g�{�`���gδa 8R1n
2���ݍ����Hv�$7A?;��"�e�ގ����4nIrl�R��I��*��z7��#/&��Zm�؉O(C��Yw?�����
�Ur]]]|�g/�ǭ�r.�|�<�����C�ݻw��u�]�0��{�n~��eX~��\}J�������������߿6;��)���{�yr�[�.r�>���*o`���!':��%����ps��FE�E(X����bи.]\���o��#ueY1����®�XY���/5H�nb�	��4v�W{f�tim�&�M�M)g�1p������/��;�t�إO?J{6�ж-�&�ݤ�IN��K$l�OFh�ш��|�Z\h��k��x�#'̣۪�7ѕo}����f�-6>_}�.-4h��ݏ��l�%ᅊ5U*t���w)����(��*��z&�ϗ��Ɍ����,����p� ��2L�Kb\צl$C@2&�@*���J�Ƈ*�P�� �[��e������>��V��� �b�f"����D�T2�O)6��v��Va 5$t7��I����V�;�>G�L�!g�xuB؈� ����N3��X�B�����si��������C�~�H���U7Cax�Q�t��: �2���{����:KK���oB��M1�dk|N��iM���.T��b646��9��	��)��l����upc��čz�,���F�!�_��3�zSd�Eu��e��:�ՠ|м��"���ܹsR?M��eB׹pl��vc�~��$ dJ+���M��R8_���1�1���D�6��Ξ�pXB\��Ś�������Y#`q��y���V��pøw �o$F�K�(����3�2:)�'�,���-��� �Fh��]��mr.��O�6	�!*���-/�ca� �J���p~э
}ҿú���uhC���)xe�BU_͑��I��;F�`n�.�����-�:��8z��K�v��>��9d��a�ߺ2W�b��g?{�����&&'��Οۻ���y��|u7.�W:	�؍���J�j<�����/L�:���;|8_\Zx}�V%�? {�n�r���S#Q=�W�A�A�V8���N�ɓ'�e߻d��)��rӝ�.4��}S�b��f���56[�ofv�����-�x��3���(�{��u�<}�x��ݦ<R���*%u�+1Ȉ!���ɉ-�Э�s+�A��ov�G��'��o���]��?P2{=�� ���8^�s�{��<I��i�aC��$�0��Z��i+|/�hj��+��ڤ�N[6Ы�:Vo4��hBB�@Q��Wq�1���֎��(	��@͉@������n;��B���_�v�����jɊ���kW&.��l,����s���%4�����r�R);�q_R�q��:Áz��q�F|��M��0�!"`�cPouD�d|`�� �T����q;e�ˇ�� yT�^����YɁ�@|���憰�D�N��³(á���d���rY�(5�{��eP�O�_�(��Vm�4+��&�z��\G??0؂*9�b��}�+:]�4[����S��Q�\��n�����׾�5���O˳}��G�#�*i$nW���c�r�kip�:�@��(I�k�阮~�j�16�3cӋK( ̀�R%N�q�&��k�qn\\��rk�;!��T]SI��ޡK�Y��m�A�P�j����� �(�j������R@�2I����{���@A4��+���#������}E�]#գ­�q0�lTL�wXw� 1.� ��s�����g�M�3�0b���Y��1�8�1�F�-[���r�
6��>|��?�w�g|�˰�oe��O����I����[�}��B��g.��t�G?~y﫯�ʆc	y%��%���+`,���#J�]���&�{�I��Ǝ?�T�)�](t����]�v7P�o��΃p����{�����1x��PN<tm	�'��c��7��)GH��Y�P����ʴv� �*e���<�|ئO��Յ���B�\|:�=�����T<u� ���`�΀�L<26eF
U��t��,u�mn��M�藾L����ޟ��)��Ec��I�?C�V֚���CTݶ��Bk�-u�j��f 1�M~^x�u� ���$`	09�`�а�H	�&�H%�h�jLI�������J�щX+�.�H�ʥ
�� �ꈀ�������C�ۈk&D�#U73�s�uF�:7@5�B�J1gLz�45���U�y����1�R�&N�|P�X��8��T�:�[*��5@�B`�8P��	���ŽD�˹�i̛*���#�����a�n�`�pM�=��0�p}�;��M.�����7?gp�jj���)�TǤ�q�m�v�)�ߍ�8v��i����٫ F¼�IL�2��c͏=������������<��s�1�<;ȫ�����7^B`����y���Ú����NŰd@[��p�s�D7�6d��z
�4NG��p�ʫ���I��e��6����X"U�" E��QУ <
��I]��>!�{��,R >�ﴖྞE�6�s��˥���I��`E��������T:��3�GGPW���/5�ܿ�p�h�m�6Ս3�t�r^FA�2�P��
�ܳ{�^�mb��{�>F*�r����Gw�}�x��Oo���2,��e�>��&�wk��I5�9rO�T.�����`W �K��ۡw�ă�eq���CY��&�	^�~5m`Б��C�j��
���i�_�,//	x�����w��̩]Pu�7�kZ ���t�,)�b���-6��y�V�P{�tL3e�y�J[�8��𲹔�N��L�����fz�N�1�D��MӆTu�o�dV�h�J��"�oݤU6��츋6o��<�x����k����/ߦ������9s�U���O<AS��1`��-4i�K�n��m6�[�+�E)nlt�0¡z��dæ��blj��I"���D����G�"BK�ۻb��V�l��&���1��CcR�*�Pf Z*��w$�G�^y9��L,��@h�� �,[�.���W��87��@՜T�T�%�H��pı30ڝҡ .�I3d�@�^e�q�իW�&����

#fK�u#ܳg��������4�k�1�E�v���ڿ?������n�*�û��Y�����7\�2�	!"39���B#��-���
0��̕�(+g�{��tMR�<����<Fd��+��5u�[�:�`�U��Ƈ�3_����'��x�3g�M���DU������J�%���~���� ��Fl�^ς��q�
P�����I3n�((Q�W� Ub�q��S�as�O ��'.e���q�k�ϣ�ܸ�\�R��������5d��I)62l/ʀ���\�=TY�;1�z]wO����z�R�@J7!�Na��ez��]?d�u�(X��y
����"�Ӹ8��p��{�wS��:ƪ�����g �B=Du��ޑ#G����������!��a��.Cp��P0qrY��m)��:u�ԗ�\����t�2bc�X�s/*D��t����'�*���2r���0��;&x����v�Q�u��j��+5յHw�� N�-hr���X|��}�СC4� ߻\D>I��VZ2���z|�XT1�1}�k5Ȭ��$�Ǌq�AMor�L?|��r�T0c&�y��>���ln�w�v��&wn�V�6�;lX���ڦ�fL㛫M�Qrk��kk�8{�j+m��w������2��?��o�evp�����=6�{��u�A�c��[\���S��'g\A�R�غ�U��z����"��V�P��׭�h�:J�����J=���-�,Hc�q��~�Q�T�\�`_�/�������\��s�&��w�}aΐ�z lah�c��;>NFU����*��%i�J%ʾh��nv��\r]  ��J\���� 'v��xp0L�b��x7p�S]�τk�qR��ǻ�<_x?�l� ���y��Jc�p�� "���=�A��l D��@�&S�c�]%Yuo�`Xc�t�މZ[��j�~�I��:]���d�,��@r��[��Ed�������ؾ]�+~�w~G\)ϟ?o`�i`���rWs��+�Nm��P$�T/�5�|x�(F�h���z�W�<}�w&&%��}�F����D��	�'>��I�Ф�W�*Z7�?���Y������y��FJ�N�6�{��z �,jȰ���B�ȷ?e��=��%L�#��A�C6̏?����*�q�s؎�O���Z��2�S��n�B+0�Y�3������us�����z���y����X˰���!��W*�X��n'ol۶��=�����a���ߕ�$jH>`WwAe�P���}U�J� 6��n��w�g�3�1;�Z�-��16��\�F=��Is�=�� ~�(�r�-V�������R��m�nԣ�̟��"�a���0�,��-jON�ĽG)�`�[��ȏ�L��5��B?^�ѩg��}��{�Ƌ�F{ܦ2������F�iʓ��SHL���R�����+�h��A��Գq��� @[u.]��/c��C�Gj���CT��s	��bZ���T��+Q�,�ŽV۬rU�HMo�#�ƀ��2-W��X�6[n7D�*�l�5�U�}˖-�Joc��Hn�������4	���}鼖�lĭvˁ(�������W#6��HArhx)��b+:N1�  f��+Ta�8�e�Ԩ�
��s�UЩ�	(�w��B���C�]|w��}�2�0$kF�au��5p_�_ϱ`1�����;	�8A����;��
y�n|Ow��+��B���$�nI���n�([��l�LV~�Sk5�p�.ɫ�X,F�U[��:l���	*P0��q��c���=C������w�-l ��q/�����	$����e`�fc�<�s�9�['^���8v��S�}q�ke\�4!#���+P��N
dC ��	�֜��M������eo���T�����Z����\u՝Uٟ�^�������{��1Rm�i���\���n��J��������xD�wεد)�^.Ú�� H�^
�L�Ҙ�����	:?a��q� U���
����w���/_�ܸ뮻:�N�z��?��u��X�eX~��\�+���j�k�Oпφ��Mx�Mj�UT���c\l���q� �q"V�պ�(���.`j���w0�`���t�UE���Y �s������W��b�d�/^�0� ���{fu{�A��<�Bw{&����(�b����f����|�G�W���h<sl���>��r[|�US�ܦ�7��5WW ����(u�$
M�̏�n��<��M�X`�4Iq��ߺbnS/�s�9���h�R�O��?5�2�3 ��x���:T��@G�x���z(����������ys���iS�fFG�R(і�M�o��\B�f]�je��/�P���$2ҥb!�����X��x+pA�8��6���A�[vN;|�<���`g��+E$��Q"VF�	�jnh��p�]ǌ�V�1���o����	��&���B�Mr�� I\���H��_��ٜMk(έ0���T
y�Ν▅8+ ��³1��gwn��u�Mc$�s
�����
�T�@ѱ_)�F�Szr>>�� (� ���p/r,�@q����~�T�wm+��*&ji�����hv���("�mX#O^���h7[||�A�s�׾�5�������Y�� ��GH�C��V$I��)Ф�����M��;�u/��{���t�=e~h��z�2V�\u�M8��\�R.������{���S��
I<����O7� �9��r����\�?�Αzݼȴ���#�3m��(�H\���z�?M�!ϵ�3*���H�K�cڤ�X#2�л(*@���m��Y����hC�=u��s�Z_��JI���E�W�����TES}��ǱV���9TUP}��[��O��@Q'>�<�K�<��_MMM}�ϻ��ѥa�a�O��տr���իW��nwz��8���@V����D圔�2��5��d��]�<�R�|�n�$x�.c��w�^!*v�݉St��o>���Ӿ}�D[�Ԉ���G�O_�6�,��>|mD��R���\�VM�����h5�4��$�ܶ����giit%�?�޽_|�=�������G��{�8Z���uW�ԩ���X'^D;y^����R��u3{�Pe��z��9��_��g���f�ԍ���|Ӽ][��Z����c���Aj�m�.�h��=Tʍ��wceUܮ�f�i�����u����>�˦�OШ������	S��iu��XQ���� �GX���`��pA?!�%a@�p�8�<�ce��F*�ùĹ�'�V�#��(�p5e|�3~�����`B�Q %
����,+���Λ���k�g�UҜ1N�B��(��� ,4 ~ x�,���bh�ر�U�x�O��Bl�[�2_�2RU��o�y%�MQ�?j�/�nt�L�	��p�K�k���pn��
yo�3l���@p�Zb��1'���E6
GGG�]��R���
���$I�u˄�:hZ�6}�����_4��{L���>��q0#�����;�ސy��Ξ�|S�S�L�U�*��'�S�1ِy؋���2_����wF�"7��wo��T�������c����8�,���{D�  @$����H��DRRմz�f����o�~���y�Ɪ����UY��W �&�g��K��=�v=-"����*�WaR���n���c��sM��q߇�uX~�a��k��K�-��Iܡs�A�_鐿�/������N�V�b#0$N��'o�3�eS>����OgTB�m��>�>p�_�c`���%�r�B�\�P�Q��6�"�~�3}"c��śDL
�JؐabU�w�©S�~377������B�a�6eH��ۗ^�����\�{�(�wtPT��ݥͥ\!x��`A`��%V��-\Zl.���,���ۇ�1pG&WXbP��;x� !��ȑ�a	0�ld�,��@K}���*b�g
p�UQ�����Q�0a)(*���5���{�G�$���
��;tHg���w�����Oi������jv7��������O��]K�c�쫚��6�a�A'�T��2j^��.E]ڷ� M;N~�N�WT��9�66��ZH����y^8��C�;�4�o����>v]��KW�.i�M����R�\۠����(�Tk��}�f��^�;W��6�)߇�ꁈرTv�6��E�I^k�fs����Ŧ��d���������q1}�Z�Hb��8�K��cIb�L����>�V���Q���B}V)�(�r%��haa��	��Z�ٳ��DA�]�� ����PY׽\�RI�}�^޿��޷���y��lS����%J"�m�>)�]�;�<�����Є��q�B`ș�g�d��n�\[=�X8�K�H  ��IDAT�0}m��X�6&�c�!A�;���XO�>E/<�<=��#�����X�$�M"�Ѷ���K����v��e�⺋m�/#_��F�ڊ�"!�k��1�3�UL�M�3��$z�K�K�2`����7�XXJ���v�M��q�s�#w�t���rc���c#k��ɵ����Zp�X�P��%����roRg�ڠrM|�fE�+�#�˱h���>L�:�쎷k�R�XE�4����v����g.�.�y!�O��r�J�m�t�}����Çʿ�������?�2$W�����ſ��[g�n>�����=���-pK�(Ȋ�·���)��ȧ�
m*��ʉ�K��%e.F6v'H&���;��v�z�'�(X7[Mu��uSw���m���b �v=�MYu�T�*�_�� e�31�1 dr����{�����cj�}�
��Β�(2a�e5�E���hJ��W7?�FW�W)�x�C����l�yFOE]�d��;*��@*�#�Y��.�=���C��ݴ��'(�{\�e*�n�H���.�gL:��z��'i��Q����,�����0�bX�Da���WS�!F�7�Z�M�Χ��1jE!�/.dꌕ�SX^��1� ��i����lq�3�k�r�Cx� � C�i�B6��3�޿ƈ����D8�N�rYT�ӌ?��t�.�
1��̼�Ɖp<����osTi�S7H�|��~)�eKgby�+\ �'�3�3���%`���k���Ц=�A�n�Z��1u�:��p�B�
� ���� nX-��v�m-�M�Q�VqK�����$��.�����2$lxt3A
��H>���bb�g���0+~���뛋���h먼S\R4h�:et	4�e�Ѷ��#������v� ���s���i����wJ���:$V��䐚>wHmcH���EV�E,�b9�`=7���>#�;�k��Oj\�%*���ϰʄ7�9߽_YK�๮e��r���_�]�ov�|�����֩[�ܷťI����~!��q���C�9$�`��2�J�ꥶ����y<�v#�<v�H�C������wb�ϞK~�@�����~�}&V����gi(�>,��ϲ��?Ry���_{��lll�+~����W��v�����
%q�H�����t���X������Y��\��1,��s\'t����p�B�S�N�vsᦩ�H�c�� �w�V�E���源��;����T��1�[K{D2s�"V�\L 
JŅ�Z�6�֚�8�P��?H'T��_�ȇh�\�>�Gg��'��n=v��k*M��U�*UxI�B�T8yEj�[R(������=��@}��4��ߪ��%j$��������cU�BW�=�U3Rf!���2jm-&pE�D�
���Ni|d�
P����I؇7
t I���b.����w�l|�<�sjc@굪�։l�S#��	 2�*�8���l����`��L	(!����X-�J�9ѓq��e{{\�r��<V8V�B�Br[�d�n������_�Q��-//녅�|d��7�),|8��Y( _8I�7����U�D��ǵ��7Wє�t���a�\ej�[ �+�`#�kI��q��JI���6�G���e@XÕ)���XX���V cn�����^���.���wޡ�ׯ��A���� Ue�ec�}�8bG�������n��$��lC s]5��9 M��W�xA>w)�(ɽc,��p�"w�Ͼ�m.0��;DO�������*�\!�B���K0��#��u���N���p|]K��!�n{�<5�h�C�sB��R7J�Zf������gbE�߫��Ӿ�w�ױ��M��%�҇r��L��!�'I��+�3�gxIY�T#��w�{��W�wɉ'�j���?�g�c>vsH��eX�y�!��G*x9�K��f�5��W�/�}����.�?���Z��>����o#��K�\�ωC���9���;.���9�ٕ62ُ=�m�����T3mIS�\2P]��㓞�(��Ƕ��UTFv�1C�DFq}Q�Q�&�n=��ʄ��%����-�"Z*�jqW�ia�@���9}��a��*gh��W~~A�~K�C�(�٣wR}���KE�Llֻ�m�Wu��G#�o��E��]����؏~L����ӟ������h� ��U��~U�F��~���NS���v0����o������c�*i~��תV��#��v�������0��Ir%�H�����j��r�b�X�T@qYN�!V�{N��b���/��0��-q"������k�8\��XzD����$2r�VdEb�� �Lrb��<|��wA�\!�
� ��\��x�9)2�����b���%s��v�۝MT��􇍃��\���3]��Ye��V[.L�eA3�d9'W�M�u���5"��,#�����J&��}
B*��Dw�m���Nw��~��?�g�{�F�F蓏?���רT)1�,)�xr�^_�W�e�ߵR	`�w�J� 8�ܲ����6/���2kl����X����@��{�&��K�.��.�mZ�3�S&(b��A��+���!:@��b7�~i����\xHH���Bڄ��@����9���2� ��G6s�J�XMI۴�F_O�ZQ���Z��^)�U\�����6�חs��9�m	���H�������?P�-�q�\G'v�x� �
+�Û?z��gw�u�K��������ʀ�2,�lː\�#/���޽�����廿����}��?;s�L���>J��d�3 �X���kQ�j5௏��h� B\�du]�h��28p+�u�q���1���6������9Y�킔'�'qcpC����R
�{i�|/�\y,0�bz������������CJ���
���1��f��#����t�3_�-]���}������}w�C#�I��>mvD�*�*U�Z�,PT�t9�T��Լ��7�Ё'h��Aj5J��_�{��Wiҫ���]i���L����i�)M�I���eE1��r�����Ŝ��t�\Thf|B�C� }uuͨ�e�%�Q 
!�ւ��+/5ʄA!"p\tp�+�-��p��UƱ8��ȝ�ͣ�0������c�A\s'��j"�҂�E?��Y��`��[�X�@��9�ļ7C�'H6��W������Y�_a�2�ZL�4u�mZqm�}�V�A���C�}��L�8�d-w�B��C���&	�%&�E��f�L�u���Z7�	��с�ઋ�oln��#���g�Տ?��I�|��y���WT,�L[��G�A�^>쿹��׀vx�l�߲���]���	�&�}�F��_����X�no�3�1qȀi�K�1��-�����N���Q
쳰諜@�����<��#n���wɇ�;w���l��X����2Y\K�۷�k��>����O��ȯ���ӿ��:��.y��vɣ[�8����G�9�w�;/�\is|Q�d�̟�	�x���TK;?��}�^?~������a�a����/݄_�+�������m��5�\(��X_��W�.��O���%|��Ŕ��4߽�.]y�� Iq#��L%A����F8�� �0�ߴ$��;%������*Ґ�����3�+�t��j3��z�+�1�2u�l&Z��D��hMS� ��<J&*&O�Z'��Vi}|���s�n+(��i�������o���ou���ѣ�Q�2E��(��mJۚƓ�.�*��J�]���?]�I�^��6B��ҷ|�!nVL��￡���4�*Խ�A�|�֪eH����[hfn��ְ�k5==1��B�V[����n�.�u�_�F�u��������U�ӓ�Ѩ1�������l�!r����y�,Reчg�7�)[�ɂ]�#;�pQ%6uKs +R@�U��V��X�@�lr^C@"D��O ��>��1��HE��X�����B�w�P�� L(  ��'ل��\�'Ι���c�:�H�<W�Ή�p�o��Q�D[�Z,Ϛ��B���
rP+JnQ��6A�i�s����6�C�Ѩ��j��e������v�kb>/1�'�����y��4�Ï>����SjϾ[�ˋ��>`bU��H#��p����kX�'���qZ��wV��א+��c��_2Ro�Ȓqut7b�qQs�V�Are����&��;�s"�X|���c����Lܕ�'$D������g�Qb��O�ꒃ�~v�b�����s-}>H���Y���w�J�k7���r����ut�+OB�zE��Jֲ+�d̤m?�	�emq瀌�}��k�\�6����&+��x���}a6.��<��,@��2hb��]WdB,,,ܜ���~�ĉ�����
�2$V�2,�2$W��Z��&F'޽C�Jѳ�I����~-�X�8�(�H��@����E map��<	1Ȑ$v� ��LA�/�"ު�=��}z��;��$��?��j5���qu��k%����
)���{!�:M�%��\U�ŒB��4�P��|�S+J�N!/Q2ƊAg��ت:%?���z�5�6���G48�a�[��`���I�|18.���ڴ��r�-���<�����_�5�>�!����Rҡ/h��N�MS�=td��ަ����8�[��@��	/�E�:̈́���cU�����ztlJ��U��W���4�[o6I��tv�E�}�u�}^�h�tw�H�����I*'LH��M�赸��UR����3G�k�B���)B�L�Ig�T��ʈ�>�_ �^��:����+���E�h���7�d7�9�k�d�"f�#�k  �q�>H�$�u��R�Iq��?/d�1�2�E] [���lI� $	����]�c��!��X��hm}E�������޽��rG�ay5�-��PPI��_=c�Br�^/�_Lj��}�VW��q��7��
����N��X L]f�$����:=C����
�&1t&�(��X����*�#jE]��"E?��v
�X@�B�����R�٦J���r�j6i�	;��u���}\��?�w���t����K~�
T-U���׽,>s�[���~��f\Qj#��M�xÜ�8��r�{����*�6.*')(8�+��{��zn�qA��L���� �#9��GJ>�L�f������)�gʨ,}c����il�Nc�<���jl۶��'N��sb;�o�����ٝ������ .�e�Q�΀%0e|x�+����I��1<M��9�n�I8q�!h��:�@�����)�)�������^Yo�E�o�RY�p����?:f�@��C2�)��}z���bu��ޜ���.W����RQi���N�}I��m�!�y�ĸA�����R����,����{��_��������Xy@o�77���hECl||��
��l�A^��뽲�O��
\oӧ����\�����-/o�,\n{�tjJW�8�kҪ�m�<��D��/��o�ѽ^Ej�@�q�`�ݠ!�u)��*�H!dJ��$�"���͊08V�ƻo��I4-���1=l�jܠ�<$ Q�W9�LB�B�8�^}p[������9�	�"hg��f ��F6��c��Ԯr�fs��OAy�
���՜��0��˙}�M�ΰ3�_�V�)��,#d�={�rw�H����0i���,'_�B��q�L��쏭���iz~T��_�>�=mP��׮��=V��N��>Fw̒��f�녍s���o��	� ����@u�g�f��� 0Y㦯�Z�����aN��M!���>mT-&f;��� z�hqͼ���GPifm�`d(�G"f�.��<�ޥ�J%;//<���\Ӱ�'Z�Q��|2�������Dm�^�u�����;���/��7�7���aj�q��
'�� =��:�j��$L�B�I���N�ϵ<UM�e�ם�x�B{8@2����������1ӆ�/~ƚĵF���O��ivD�Z�|G-��ԃw��l��qS�/��`���$~=av�f�d�L�/H���D��Ϻ�W��i��7�"�l���/@�9m a��wJ)�P+C�J�h��v8uz���ٲl�keN�n�e�n1}�r����r>i������j�k���[�R�;ثrro��z��벻�T�E������~�jˎ�--Ӱ/��v�ζi���aAq[�����m�\��o��������88AmJ���z���`?}��%	]��R3pw���?MyR�Bo�R6��8e��d�����r;*��dk��������I���B�I%�z�a|����xH� ��ܦ45�5��z���;<���q���Z�2�J�33b�˸�e��e�S満x����&[Vt���z�x���h�Q�}�rKm�g[m�%��s2����K���fE}7.UꓓTȽ�\x@���G�3��`y`fQ�α7 ��`�s��H8��f�!����rG�f�Ě�`��
��H1���DI)FN��%�T�z������ZN" ���Z���T��RS�x<Z�w������Y�������F �i2�J�#xx|o���S���&g�6v��.�����������eĸr��n(=�$��ql(��$�� ���-u..��uE�8i����|{ ����DHN��_m�[%�wQ�E{gLM���wC�Qyz��뢃�ztƸ��^B�x�dWsh-Ss��C���i&��g
��������,q�٧�Z��%�K��C�3G;%�c@e������lf���;�l֪͔(5�Ѳ:��!W�I��J���pq8�i��� ��(L�O�)�#��F��ű��QV���EJ��{Vry��a6�1�$�@��a?qKD2*�r�D}����!d�!��-s*{,n��ho|��t���Ow���L���|ہB=��|�^�����430ǵW��L��׊�GR�FJ�j��(
�mIχ!�H^��`J�D��+r��6�ԁi�93�����GJ�D1mN���D�foF^��t�?��r�G�Q-|�Gz�ݬ�aT�{�u�ӻs�]�a�r��	{׹��}L�_�o2�:>���J@�ʑ�?��o�<j��^�ѓ}3NK�].����w���~{�~Z���>��ܦء��z�UG��x��ɮb�b׵{�4Л�J<��/�˼�H|��r�,���<�a��o�ĩ@[�)�a���hi���ez�����A�ʺ0��b��#�[�;y[��ܜf������夺i���)�n�I�2;���BPꕸ?���H��hZU�i�;Y��=}Q�7C��c�!�eO*,VUAӯ�t<b�V�o`�L��O��sɲL�4�(eX��v�	�=��1�H������^�Z+�߇^��*[2�/�MF�j�Ş�����~�����cX�ďx�w��<�DKj��뤐�7�����ڢ;�Y��h����� ��Xf��8���K�_��ˇ��g�H�~u�9�I�j�/䳖�{�JYVi9����o��Hj0��r}â��׬j�"Z���.�6a���h��ЇR#B��`y����s]]��b�Cp�:��@ȣ<M�ZZ�ã�C�b$��2���T�}R���|�ۅ������i��>f`|3>��A|�^}T��0a%���N����O���BQ{+n�7� �n��~�41 r�!�tdZ����X�+H9�lE!�Bʅ'F�fܥt:�;oC�o�8�%d	c ~2ͼ] ��o��J8t2�$ �Ó(�\:���qc�_���{ߧQ�P1y�l���ҩ����@4@Nr�I%������A�C1$�u���T���t��v��ht3���k�h9F�"���s�(�83�aq/ݣ9��9�V[
#_§��E;5�b�géN�0LŠC�UG!w�%Kr>g�kó#�]ߩ@��A�b�(��zS-J8c�%�cH��㭬��W<>�4&\12�.f�aUڜ.F�����pO)<��,�9j�pQ��g�����nR4c{��.��q������ڌ�tx�Wx�.��$$��-~X4��X�������S��p�� KZ�%W��P*� �`���˾�v|	���B���^C�i8E����}��s��P}裀T���OR��Ilh)�~]!RVS�_�#ٯ�Rx�$>�T�k�3[G�4�%���H3-��;����$��ix����7r)D�#
z:dhK��4�Aˁ�E�tb�Ŕ�Q�LZ�S�;���l�����TYQLK��N
�&��o�_z�DXQ�H�Ūan�Y��)��}�F���M�e�jN���m�?"��8�f��p���``o�e"j��f�h�pe��d7�+���CM�z��>�MU�3%/������gJ���kG�m����d"���]���Pk�cu &�U�����ރ�!�y��qQ�?AۃEc����3�\O=t��l�m=yP|kdO[RӘx��)v���*ǿsC�/�D��6��*�A���v��q"��H�HPXI��T�a}��;�y�O�$K��y���.�"��'2Xj&2� 0�� ���݇A��'��v�2[n8�I�E��'N�;� �_�
�ڐ������Gx��[R���jm-X���v�|N���~����sZ�zrJ$)A����ePԦ�4��Y�tuI ��2EYX���T�MoQP]iR����.�W�Ylt�pvY��/�����h�N�0;��{J1?,W��!�dYE>��7[]�:�����۟ƨ�Ӊ4�C?|ebS]2�NϽ�b�OPи?�ˎ���,�1z�FF�-��@�N�C�ȥu�G���m��!i	���4)��J^��"���lr�t(����;bl��27���Z�_N��UM�bH2�d�f���7њ�~ˏ~�͢M ��h�[���;W)_��7 �#y���?�4=��R{���GzS��s���m϶���f�A�_�ꢂ����0��@�RGoCGVFs I%W�Ϡ�3B�l$�7��lv��t�9l��P���+�w
�gA@�c�-���aGkk�\��锠WD4��8<�G����[��.4C���haԲ��n��)r�ruE�*"	�\���!�M�	я2-�H(QԂ�LgJ�~1t�}62�n�lzn�0Y�hk�6�:��r��b�m�3Z��˱:���a��́V��Ҧ��;�l��1�J�:%����� sp� ���L�;��^)�I���H5��u�an�r��d*rA�jQ�C�Ƞ4J�s>�5a�����@�22<_l׶S,�q�� �t��݇\*^&j`ŭD '�/�Y�B�FQ#ui�7�@�w�8���3\Т;�4�C�����?�'J��=�7���V~u(�^V��'ЮP!�ڄ <4NP�]����$�Kb)n��f���1-kuW'�h���&?Ǯ�녽�E-X`�i���#�e|"��)�Z��$��t�ñ
�hы�X&��d*�r��0vN�*�]�8�e(�E�[ꞌ�挎�@��:����R��M�{bd�zy��ײ#c���ۼEC�;U��ei���2� l��˞@}�V���J����˟_�n�H��#�؛3=�&���\J������޻,�c�i�]v}h�к��&�f��M<����]�C��N����w��\G�.�i�]�
�G�	K��S�ZW�j]QC�m���{���S�s�4����Z[����%��G�x�l)��y=s���:��1h���/����m�ܡ���.au���9xxxwAQ�S���)$ú�Y����]�����k�6�W�*��؛���"��#��)P ;iRh�0�����mSu~����S�r�1��bL�d������n�v����L�=�ܹ���f��G\�f�j�	P��B�ǖb�*=�5��J<���]VS��O��̉$Z"t�߈#_�6
�+�F������]v���Mޠ)��o�Dp*���=��ˊ�Ѩ���\�&SO^�ףkPsc/����{5Z�R+��p���~?O�=t9�hl���:��ۧ��B������-�}� K<��{�WJ�Lk�@�J�Gr�����\*n۟��{1-	6ܩ��[_K�)C��m��Vev��.����OT����l%�A`��r$�Y���94#@���C�-(ϯ\+��a�`=bh����SS+�����t���|$��Ug9�Q`$�C[h�	Ӯ�}_�0�߃rc�^����A���8���Wa�,QD�-+�����U43+���Log��IO���bTg�8?�>Lo^����_.�\�tF��EA��?*��y�Ln��E�;'��9-ri=ڌ�Z��F�3%��O�9|2��0�2Y�����Z��!�����˨��@���%ݿ����/�8�	F����`��/I~�$��3�jg�c
bٱ�l9zG��%`z�]�T@i���;�1�Ο��>��1J2��k��޵�&l^LĽ5N��z����Q�Wv�ì)�ٮ_I;��]��gSa�ڏ����v�K��ݥ}3w����W|Sy]E���#�_�C�Vq�����s~3��W�,l�$}~�ydtv�H}m����ͪ�a!kY8�#@v����)ڛb�	�W�?����D�Eo�!�\�W(����LI������~r��Ѭ��}��������<f�Me����<�� �h��[�	a:s���<)�ϓ��1�~'����!�96�7�aR�<�C��fE�qj�������g�1��ˁ�<�zC�k�ߏ��[�+D��t��(�6�*��V�HFGC8�<��i�`�B�AFe3i�����ai��N�5�x�_	uOyhiE	2N#�İ�pW�B���.� ͈5T�v|;�t�q�%�w��Uy��b��]P�.��0ϭ���Y�1�9qW�@��kҳ>��A�������unTJд�W�x<�L��w���o�e����;L8F-;pO1{!�vҸ���{%���A{~��\
w!��좺��Y�!)w_�HA9tB5�ٌw�^Ui^��L�:\���(A�8=4�i�b);:.I$/��>��U}�8:ٌ�ky�u_f4E��}���F�+/�$)-��������z�*@M�LcӀD��p*���|*tF:�F�}�-� ��
g��������o��C�G���jN~~��ӛrI������##4�|�1��n] �A�*����`'�����岍M�d;�RR���N��?��}v�A+��1l+�/ZK8Qx���,�������ć�m��¤3Bv[#b���l�e}����G*-����G�[eF�p^�,��o�
a��k�+m�2$�!��ȯ�����gz��$��u�����~��@��L�j�JSd��9���~ݍ|rcB�@UP�3�t�떇,e>.�$�08�q���;M��+S�r�ir������E�UFg���CL'�\_r��h�A�L�՘��n7���-��ym�m��6>+nc�+mڎW'��Xa���� �*����9qd�� �ϗo�����wW����[B�P���[3Y�Tz�-&3�u�7��<����OK�R�_~�V��D�82��]�w*�G���W�5�p�[�V�
c��
?x�FS.�$��+�g��Sǩ�X�6����k�JeZӁa���3{�-�UȘH]�܅`=�}6<�疲XC~��0� U�"5z·���
,�i�#9�ڪP�0iW�>�\�:��'���ې�}Z�\���R̽踭|G3�r��=��W�'3h�`��2A��*���|*��p,��G4�sr�k:)J���u���7��p�c�
Ύ��ޟ1�?�,�sI\�4�e{�p�R��׆_v�'y~�5���Z0
��T�)�C��C΅���!#m�k�̈́�C^,�qa�������i�:P�  
���nA��Ly��lG�?�>�- )�A���t1 �MfCe&�n�a�����H�P���k}�)4M��On�ɦnjt�7�7^���Q����_�&?�D3��}�'�������;���r�	�ٺ��  $��5�^ݘ]�A�:�����_!�������@A����w��j�y�,E���� o�i=���kN@�:���>�d��l�t��
1�eR�rҊv@�\��9np�:I2Ҽ��0� ;���OzL ��}'��+����NL�F4�q@��w]�L���'���U�� �˟���C�j�`�5旚��$��^e�(�l�ʸ*.�u�e�-mR9�(�H�=qm�w�z�q�kW�|���.�&v��NMY븀a?��'��NL׽��f�^AG�w������p�ϱ��w�����-��������C>c����ɮ�1�%ș�=]� {k�f�"�d'~ϋ�����>��3E���.o�:8�������"IK�&�bk؆�j�}v8�h7	V����_��h�mB$$F�����*?�ʆG�!����\x��¬����~�uW�j�PtHt���&�qw�!�wb=3��Ӌt��k=ڜA�B�E����ܒ�	��%�P�VZN��K��~՞�2rw��LW��P���˳��7���S�����T�"�{��3ob�Hqb����C�y�1�5hL%�6�Ӡ�I��f��fU�<�e��Q�5������<:D��3��p�\.�yy��n*��d���Tb��T��x�]z�)���u��c��=��P�J���^#�g�ͥ/�r�V[e�����S�
���ſF�!�_e���h�Ah��Y�:�ނl������\��L?�&��2ր��jV��\7��^��e/��k���Ӳw'���픢^�����چ�]hc3��eq\K5�O��� ��{<Yη��=��nV]���N��|�ќl��V�hY�D��ۉ�d�s��*��H�#w-l���r�1Z�ߴ~(�[~IӉ�� :��;ތ���e
�!0M��7�
G���^2D8��q�{c�mO�?b�y躬	L���� >�PnrX� ���t��y��@0u=ū�S�YsW�(�y�Z��7���.:��¶�f���{�S�rmS�52>���ă2�^��2r�R��l2 �Q1���"&��̩n���,cP��@�Ӎ�k7ْ�����x�����o�tR�׀���t��$M������G�7|��/���n���A�c{��jvd�xFI�u����I�(�uT�~q�ii�{�~wǳә:����N�'�߀\� �����&C2<=�&2���:G�ڈ��YŎ�u�8V'���`2����,F���x���܌U4��e�,-��#�9hJ�#�ʞ��Ԕ`t��7��ξ�I�zU�Y��f�m
��+m=�E�3h试�?
՞��.Z�U�3��e�iXݨC`� H*�w�4p�ڰ�V�~�ͧ�C'�5�]@/ڂ�-W��ҭ3��5&��*�w��½��-c��9p˓��2H�@��\|W@�C�W\�~��~�;�9F2�J�hX����-���3JiKY}�'�TP�㺨Xip�#ɨ��ސb����Uu�T�p*u�>�YdT���sRon�	�Y>�z�nu>'��X�͙�ӭU��BX4�BxS�.!��@E2M�
�*���[��բ�q2l�W�y�Q�rލT�gPG{?f7�T���9��>�0�-䰉
���'*�?p�ZJH?:�Ơ�RCv��j�1� ��v�C��4�Ǳ��@ VT/���h���,?����8����ε7bHD	�W�`j�5m�j��*O8��o1�E�N'iz��[wf�-11����8DjP�	��r/Q	w1Ǹ����['����#��#�B��M�}g�2x�r|�:���b5��Ǜ�%�����+��-�=v�f�	��*�<�yi/���� )�
#�G�[��O�����˷�{��)7���f3����|�qs�/O�U�}~���;$�]�#���,�!E�39�Ѓ=G+V�V��*/,�4���Uf���a������m���޾T����E��\_��zK?7���������]�Z��҂�Nr��?���|��|�-a>ږ&��F��3�A�^N�~W���d�:tl>`7��L�aF�Z��	��x��?��.K����~�ե�?UȤk��/��� �����_W�Ӈ��NPԴ�N0�����Q$��$'�=�yj���4G�.�T���N ��r*���IV��̺Qq4��L�p����)̢W��}G��9�l�Z�*�0yL)A��+��C�dĬ��(��d}Cت�H��i�G]߾�FJ9<ɫ�qF�8�7�bD�
���,�7��;�lt.~�q�z�%�jW�̀0�'�%����R�SB۽>ԓ��:m~�Ąm�20c�&".ō�h���Hk?:�M�>��F�wF�B;{NC\8��������dmfuwӴ�s�c��R5vͽ�L��dfl��ơw0b!$2:�E 	���nrۮj��hs���U�Iwg�6�Q��/s�:-D��,�,'�sqJQ�k(q� ��PD�~�׎�{|*,���2x x�N�g3QF���"=�U�y�Io�@q�����-��dm8� ����&����<���49K�";�m���7���b�ѤJMk3A��D����`uk��a|��Ӂ�T6Y���4z?qq�<y��.:q��c�����l�s��*�����kJ��,Ko�r>Yvu��ú������V��2)�k ����!Fj�Y��i�:�g�*-r;aQx�5��,z����w� ��{��4=Ouy���&QZ���S�7�Ң������ѷ&��dyǼ���M'n�n��ޱ��"2
gV���i����MX6.��(
��'�Z"*|�^	U��M�_��<��ۯѓƾ�Y��ߙ̛��I�m�f��:�2��nY:�V[�F�<{98n�>.܄˥��d2&�㮙�ƫ��wφ���C�$��� S�[�N  Nu�'��/R�}@����O������j�Ԯ��{��\�*Zh�����b̛_����ʓ�D�
��q��� �oF:�U>�.kek�n�O���g��d��-�E���-����5�����^�]Uq���GiDBQ�L�(�t��yUq҆N(��f��v��l|G�)��a�Tr�gix�y�g�,�K����nk�F8�p�]U�dc��~.o��sy<rj������~�~�~�(�^���E�
���XqOT������/~ B�Vj���=.Du�s�s��R[K��3}�d���K-�9�_�����8,I�n�z��������ԩ!^8�H���7�~�v5����f"h�r@hJ�&�Azg��?s���3C��U�Dtd�pP�y$��7ctd�"�{"\m;@��6�Π�c�'x�1�g����ݮv�
��1s�
`���}��?&�����T=x�����x��/�j�2�w3�zu�E�t�d��{c�q���܀��o�
�����G�(���-�A��/�s���u�J4���8y����>�G����r	��$B�L��i1���������=ք�X���p!l��i3� Z������Hń�-�ş+�8,J�U]���-H&�<!�����ueJ'�3xLB�%>�>��E�|n|s��Ǹ���9��DՕ�����sAy�E��in�Y�s;4���m�m�+�}X|���Z�0�/#Xˤ�o�S�6�޺=��ɷQTp�"�i ��o�X8ң*�rI�M3v}�ދT�#� ��g!H���D����_��y�v��5D���d����b7�������J,������ƃҵ���/��0��8!��0�����`�y��9��[�=��P�,��>�H�j�0��^k)!D �N,E�9s���24Q�g��K���n�eՐ�j��|�v��cA��,>�5�56]T�LP���z~��O~j��Mj��q�JI	5=4#��IG��v0���]I�p'�:ܘ��u���p���	פS�cM��/k^�����6nKiP�i���tw���|Y=�~����s������hx��P+��V�����g���&SMZ>��7�+=s���8����y�F�7vV���-�&@��ۻh0�bfu^gxO=�AaIpq~VCq�d��"���������J�LC��<���ɹ�Ƚ{ai�1��a���C���>0؄�C���lZoS�3,�Ì� g5����=Al�J >_/w��C�+1p�J� ;J��a �ا��n���$2�|�S��r�윏�����K�l]��R�MA&�(ˋ�n�%n���v�,�Lu���&��_�&�72V6��=
�D�ME����l9O��a�k���p���a�.*�8��:J��4��Q:��fw���t�y���~z�O�6�zR�T����zv7�b���M�C-֦��LTn�=?���D��� c���x�a*BGc�[Rϖ�!,�I>Wqo׼���0�-�z��y���Ԕ�����T�^�]���yk,�;r����W��F4��`�����*�gI%���%L���1��ˮ)��A���ZV��s}[������[����[0����+Ig|���_�������kO�����_7c%�N��������^�P�ݽ&�P��8_�V�_��N�+� [��&�f��xd�C���g6�1�P��l�X�h�����)�����=ᶨBrƒz��~q�n1�n���r�$��F�첈ڭ��I������D��*���b!ں�[���O���oi��-}���d�[ꓕ$&�L���S�?t��hӪ�lX]���*�MI�+]DK�04˩�CGl�]E,+Sc�v�$�����7�?���0_�Y*�;������K9��&%��J
^g�.�i,���*Z\��i�|���j�6���tW�b�?r��+ n��T������=��X�� 2��бBL=�((QMK��� ��?8�9�^�����qPNTPF�d� s ��g"�T/@4,��Z,Q��S�,�+��(�Ǉ�ky��+�L�ǋ;���7�v����Z�ۍ�C�C(���y�K�X�Dϙ�)C�pdX��-��W��Og��G��uOR��H���]E�͛�� ^NV�E�z������-C� ��u1x	�{�ou��o��zQ���Rs�eQ�Z�ێ��z������n�k�8����a��\��J;G���`#���ޖ�f�:BH��e4��|.�0C��������^�j�Cv�]��Hra@Bɤ�``̍�F�OKC�{vҿ���A��
�߲�C����a�)�,a>�4}�(���`�b7����7�I�=�n����)��E�t2����s�@�g7��Q�o�{mû�@��?s��^�t����)B������͙ĩA�L�P�?u���:�O�)�LL����(�4$���I3�@�<!�S����c�?;�k����\�-{.�>�1�,A�Q��P���b�36
���&2r8K�kyI
6#s)5�.��4�
!�2��I�j�ZH���RM�\`L:��vT���l�u6ʥP9}�H�b��숆C��$��^�xO��w�ib�K�	;��ݐ�+�#� ֋.���*���n-6CSc��8���<�^��XUj$f��׺�y��^��	��`l�윕��J�K��.l��$Y1F@���ia�.v*���}	�U�'��"ew%\rӆ��F���q{�՗�
}RS����x���rx�n��<l�yM��>�X�$�eEM�=��=#ѣ����okC<��9sz)�}�44�}zf��a��Qm���6x�xR�G+!���:XMha��%?��6�!�)a��L�/$�&DM�Æ�n�r�bH����%5�����ӅVVVؑ��-q��;a��@�D��N�JF�6��7"^ThƜ	����*�����A�v-6�i�C^����5�}�r�j��浪�?�-s�D�� r�U+v�;�!�@_��"�sD	�l#^Ĳ'�F�-�Y=+ۚd]��p��"m;��w�ư�ʈ<}�Z[z���yu�����Z��Ʒ ��e���H��Tm¤�.�������F�����Fq����*��V���?�I�}�ypa�0�ev�OG�26����$�U��G������
���������6�i�+"�mO��]�����i�K�I�2��Z�R{�����ku���?�v�0`z�,�d�i��V^}��,1����;j�/X^�,���NJG�~8R�r7uU�ߒAw&FYo�5��6�ѡ����R�`�x=w�>j�S�t�@���b1�:j_�/6�?}l�?��c��;�pb���CB� D����J'}���6]�<�RC�M+Bwae�!@[�M�B��UI��G4����yp�J�Ȓ��M�Z!bV�����S4�յ>�
��wP��E���W���^�ᒓ!z�������V/��t'�"��"�������%�ѕT���T*�P'⢑Otm@۲Ӆ%&�$��	�>��.���ϩf�rN�dj�Ȓtl�Uu�K^���)��W�V��[�6%T�-�9	���^4f�c-�W{@�`*�R�tJ��|�\a88��k#���HQ�i�`����y8$�:��-o�_'�R&��2�Q�N�@e����v�sY�:���ܳ�W�Ǔ��A����+MB��f�Oxf���tZ���Ͼ�G��rbF�Zp⬊�gb�6�g���B�6U	�*A���W���$��3G�o�8�����r4����XNF��9�ڤWDx{����Z�����F�6�.�Y�ް��wH�@+�`�$��MuF%E��z_O�CCO���!A��o4�4����ѡ���-?Hö�U�0�j��:�y�-1�-�3�U�I�"�QT�C�EOwa���)&v8�}�^l�W��6�0��̑u���Z��Y��R��f�kaF�*=H5̈́	��f�S�,J�)3�{l����������ȉ�_�������8�������
�n�׮.�2���$���EU נ.OB��@E�����|�>��������!٨=_>㕧��� ��-�����T2�]$���Tf��}�0{\h;0�rIx�;v?�P+�Bw��<�:�>�	�H�{F!$	]��g�l�������dNx�2�BI�����!�68�#oc"����|C
���_���(Y=�6�A#���o�@d����*f��6�e�pܪ��t�@z�#�����D,�x4�����Ɍ�$��]�2G���ƻ0��\�mN����.*��Xi�7��`,W�hRپ.��v�k
�8� T)]O�i�X�����U��?�8>�r��1x�����Rb�ö�mG+5�'�*q^񺘣�	J�����һ�{Қ�������l�@Ml�a*�ס��z).�`qB�ZǕ"�\s�A�P��JH�����E�GK�*�#Ś����3Nw�E!ˊ�X�`Z��K5�P�,Gg'��/�߰q�_�f8�˴&�n�T��5׬�%xz�U���[��+\۔JT��Z�r<3&[^��{�;p�ٛ|]�.��U���/�^r�_�5-��u(��^|�SS�r�Lݟc#63�r�`����U�b�A�@��t_��F����+��7H��f��<��OI����o��������T:n~�����i#�*c"<���$!���.Z�J�˘�%�-6�X� ���j0Yΰ������*H�0b�@z���Yh�����0��3�zU��تM��~�,i�\~!<�`P�ӒG����Pu��"����J�z��a��	i��������cN��FK��܍�ޜe�5��²7ɱC�#��lf(�ŕ����N0���~���t�D��dM��[QtZ]�Q!�c0`4��ʇ��=�n��3�2�*��(��u<�u-A��}���0�ᨕ5�wtp^v}J�3���H>�W�r�$����p�-�gݫ+|�_��!�h�ū7V(�`�����Ie7��L��d���n�PĿ������l���^��=�7�8f(�>���Ժ�+i��51'��^p��kGsU�O��`���Pw��s_�7;t����IKK��Z ��x��9x�Ց����Y���������]v�-�{ZZ~T�^~��8m}�;�~~XO8�������I5����qd��ϕ�����}tt�p�}���orΗ�v��B�&Y�-g�)_9��$=�f���T�B�z����͸��A��������z�|����ؖ?�fVS_!W#8��[܂�K��~E�&J�*��v�u�:�AQj�[�*Lxa�4�s >��T�g��{�������Հ�Q[󰨿w\���uV��`[IX[?�	�ʋ-!��Y�\[�W����*�k�=�v-M���_�eN�7�2;���j�*�S`W�F_1�F-�:�Ojk6�z���_zE�ᅑm�M��ۆ>���r�֧���Q��̾m�o�?��ҥ)iOE�,E�� ����UOM������{R�*��U��Q��4*�����B�`s�TE�O
�A�n��B��$�̆ �#/+�������Zx�Lش�vtV�����e�L�F}�-�F�aѴa���2[S�R1���B�,��sجw��4�1���j�v�)�Í�k���)Z���v۞� A�C�P���J���9�T��@Ȭ�lı��VվN̎Hﭢ��.�=y��|��$O�oAg���8�T�7���A�䜉��1Q�,G���?�v���Ra�[-d��}m��H3�������G����e��d�F�����.���3B����%	�܍C�%0����C�~#�5���3���O�u<�ܯw�|DN �.'�R2��R�f��;6�����Б	�4��ٱ}α�MwY��C4�ƥü��e.���ٞ�m�!_m?������x׶~�N¶��}~tw z'�e�O��Yv�6"��!
�6NW���y*D�G���,�����ݮ4�}�yE5x/�?��s���
h�I���u�?'W&���4���wIC؜!� �~7~(��2�	��W�$ŌO��D�;=��x��1zv,qC�b�+���d���9G)��/���L�ؒ�XV!�l7z���N^q�:k��5��+���`��U�XW�Ÿh���u�&�h�&��Ȣ�/7b-��N�x��=�?=b�D�Ƅ���A�û)(hԺTTL􅀟�jBYA�m<Y���#5	*���{���\u6��!FN,U�ˮ	�?���'ɒ���Kl[U+J�T�����4�/�|���	c՞w����Nf��3?��~�ko�������xO7�/4ڀq�x��a�rҿ�jXb�
H8��v��l'UF�
�2�|���i�ō���e�p�4��:˛�E:FDR�_KCI5T��F%�u���j1e�#��v��0i� ��V��]4A����s�g��? ~@��_6u�0�����+�abÐl��y�������J���V�c�H�׃[�qy���YcU�\1n�33ӆ���20���~�\w�,�U""������x�Ty�2qTl,�x�p��	@0�d�L��a`�4��<R��u2'V ������qc����o��p��@������/���w�]�'0��3���Y(\���֙WL�^���D�F\��bA���Eǽ�ɓ����U��ĸ�k�p��2���P6?�%J���K���[w�ﶎ��H�~��}������k-}j+t��sP�϶�8����X�젽���J�K�➄���ε`��<O�qb贵��Ϳ���h��s+�C�\I�`\��n�N�@���n���v�6o�=z􋙙���9��a�a��,Cr��I�����޷����I���[��z�ɧf�9Rð*IZ� ���BX(����)}���\عv�k��x:�!�#�����ueyQ�S��g���sT-����Z�p��<�Q���9�{v�͛�U3n21Y'��"�21(�PIa���S�;\��fG�|�n��q�Bl�-��b���ƺ�|�>���>Xd �TTU��X�ϟ���
�0-2Qi��S�X��L�uE�#Gh�{ߦ�����T��_P�އt��֟3y}�D3����(P�rWǅ��,�tT�6�E-��.����힞P���r��^���_�D��6պ)u?������ֺ�:��:�y��T�0���V[%^L�
9�@Hv�
�b��9��30 ��PD�S2!a�V��T��3�=�A��s[+�ZY^�c/,�0�eyi.� �y�p���3�!��[�h�
�f�ܽ{�j"�K�)ԃ~���Xaa��V+Z1�Lz�U2���8�}A=P���� ª&�I7F�s��K���Jb=l�P�_��BA b�*���$	������	���d�cN��!���ɓ��Dߏ<�9���}U�I�A��%��9��\��5@��ꏑ�Aw,�*�g�p�.�l�_����&�I����;�r�uE������{P�D���<�#����D��M�U��ۯo]�L;D Fޗ�$y��w?d�/1?.�껾�[!onq,fʵ��VC�r9D+�Xɘ
�p�j�˝̑>w�P?���|o ��]��<��+����[�8��!���5��ٜ}9�µD��+֔�I����(�������|lr���7����p�}����eX����2$W�X��������ܻ~��i�g��c++����`킴��,��B��O~�H "�ݴ�l�*������f�6�W=U*D:쮨k�Ղqۿ�5������7m������yrΛy��C��\@b���h��%��7^w���:����x�n�eY�@`#ɀ�U�@��(��V՝s�3������ά,	G�&.�n��t�~���z��'~�틟Ҋ�E�V�;�m��B;�Z\�ŵ5#��i���������j��(�@-���~`��p6�b�@�����3�fp�^�%?�Ya�I,b"���F&��Q�;5U�E���|�O���f��у���G�9�O/ ��j�������HT��=��ɔj����)tY���	�wz����b���ح���Law�};��)��d^}�ӧP�pY�F���7��ݭ��lm�{��s�J����(
Ǌ���H#@����$���	���#�rF@#�V0x�Kč���������p?���*Q���0�S���a�(�'1v�;Tn�&�yl=��Z�?������q�11���u�{c�a�+�� '�>�R����{L����L�3&IB�D�K� G�V�l�%ʖ��	e��.����ͻ�eW?HHʝ��&I}mT�4' 6�~TO&Xb���Wb�@���0�>u�����ᇿa���_~/^2.���N,&�Q`�8�w���z���^�ɧÿ]�+V5�y(� @?���
\��xX��ͻg-�'u����s��ZЮ��Ċ]�"6�KF�����C�qC̏݌1���u�萅!����@�.�.y��#�NC��r,�G>�gk���DS��X���1Q��խ�Mt�"�I��,�b�k�&VPi�Ș�2!�I������!\�7?Wl�b.�2�F��s�G���z������'O�s���������e\�e\��ʘ\�+��dL.�ڵk�T.O����ZM�1�(?T��t{�# �%V�����wn9��t^?��b��є�Y��(��f]��kqv=�}4����Dj�
�g�>�EM��]�#rA�zahR=�8�	秐P�ݟ�I0u�+/�#�L��?F��f�D����]�'�w��*-��lָ�%�	�"�4G$-��L6Kd(�N��;U� �2�3��\����S
��֙IU�x�]\�`﷞A����W��r��!=�C"�A�G.C��@��D��bX�j������4N��Ee�9�MK|EO����6���J	�fE�x�>�,���XNQ�!AD����`�;����=�|G��� Y� u��XI�@c���M"�ȇ�"jZ��p�R���1MLr�p�?va�������h,'��k���ck[y����.��5c�b�� UWg@��6�e�]C��2	�09pA��JLlX���9��3�k#~�I�#��\�
aw�C��X2���\X��g����r��� {���\׸�reG�V�>���Xq_�����}�o����mLL��|"�j��n���f��&���(�*|���kȊ���F��wʠ�8~ɕX���Xˊ\۽�)؇+��p@�X�B�=!pۧX
$�Hn)�m��Z��%�vI�����}o	E�)!m!@B��y��Q��H}��/���I����b�?$��K�n���Ș�S΍��bi���qZ�,�[ �9?gF}Ӧ��9"�{�܆�;.VM�c���Ɔǉ����sǎ��z��F�ʀ�2.��X���P�#Z*��g�l���˥b*�8��Y�������f�Z&����b庞���$������	�Q�_S��x��^���ͺ�J�;��;��v�ǅ��;�.]Dꍳx�Z��ͫj�]g0�gڹ8:�z�MUo���[���7���HǓ*M�����&�bnn�������͢ke�M,ǝ]�|ٸV�3��Œq���\^iG�� �bmĺ��fR�{d��"D�5t��'Ԯ��󻡷�oL�m���.���l������b�[���t�@|�%�9>����Hq��Z�W��8�S�J�8p��G��;?yB%/�a���Z��K��K�:���|��jy��|���5qtm�Ts�"1N胨� ��W�˫��j��tY���(ݣ��,b�F����kJ�dQ��c�_6�K��߅�$�xC�j��ar� ����"�N�:�w��2����SV��f��~f��Ȯ3��s�hp�P��~ �ؒ�J�5+f2A�ky"��a�*K��' [�#*�;:��$��~q=��u�t1�O�8�@���O��YH��m��X+ߺ�1�nL���z~aN�}��x���}��7��ī񼶄*�Y2��]M}��RC֟�H����;&$;�����]wA�2�Ņ�ʌ�v�sH*�㺫��
y	@����6��ߍ�b�$\�����'P�-=n�]`P!���0�T@�c�^�B��8n��k���ɪ�F��o�]�Z�B�h	���:�� Kz�Mr�o�p�=�Ϥ��H�/Ԑk�k����.�Nلp[8��w�x��O��(2����$��?or-X2&$X��@�&j��pӹ��'N�y�ȑ�i�x����q�q��.cr�_�XW�$��CD��Vk���~��Sq�٢�k�.	$!5XćH�����֌0�	�o��t��8v	>K�#��h�W^��		 [/m�dLe��X��Kh�7��ϞP�+:�x[}\-��ʊ�<}\M=���t!�hA�w�������AM�Ɠ:�L��j�Z� n&�`�A5�WSE���ݻ�-�M�/��l�,��u��cļ�����z)t�6�ud���2
�X�RK��=BI4"���ݭf&��/��ϟC�ëX�xKm���8��.v;�8�pR��dfB��
���zq]��U�������n�ѸZ޳�|�;�����˸���1f��^~S��c��o�����X&R��.x��U*I��e�5G�gܙ���u��Q��ږ�[}51���X� B���I��� �c�l�)I�j,S�)5=5͹����j ��̌�>1hc�� ��h\���[�x�Ō�3��y�D�O6�r&�_�#�Ty���Lds��'���]�e�Y����1�᤻|-�&�I,eBL$N������������y4�׼��Y���X˱�Y�lrl:�K�7��ˊ�ֿ��?����W�ϟ�k��f��I��q[���V��� �b�.`����K�nJ�B0�$
��w��pcً�0�Ƶ�;���2�:�1%`Z ��N�u5׌�d"%�.������b�B�8�g���G�~� hާ"����Cޏ�x��}��{8|GK{��KS(=.V%9Ƒ�I�v���W��EP�y�F�a2�����6��䚲���a�ݶ9��P,D\^�>�:H��k9��������L�y+�/�+��8����^S����۷�x���_ѻ��W#�8�q�q��1���S&�@ܺ�]|`�X\����.)�&��d�����1p�>7������Gۃ�u��>��1���!ram:M�'b�P����u��ULMdp����k�,>{���&��͍m�ymQZ?��בق���u��V��'��j"5�b��F��b�����$V��B� �.�p��� ��Z�p�h5Q�wKd�Lv�\#AD������G�*��!���\4�^$��V��$&�|�ޑL*�__A�����Q~�,��5��!�8s�@�H��<�'���*�UJmno�S)�3I=��8v�٭s�G���;��	Uy�,�^\��w�����l����z�ߍ��c:�/����|I�
"] �	�bZ	?�����q��溪���4U���#,n���م����o~��G���RƊB���E�s��w5]5��A����Yt�j�������
�ćX�-7x���g��_�n�M�n&<<m��vV>�e��ل��D�|.��q1	�Ș��晈I�m =' ��^_�7u�l��*�U�0��Ii,n��Nz����M�U�h�IN���kr�
��:}�-x�o�ԩS꣏>¯~�+s���E#����\7%E.��f���(vc���	�oN�����ZF�덊kȆ�k���^eUG�!���A��	!�"�.����@�;ѵ�aD�\���߈5�s����%�w)�	��'d$�|��_H�oc��1�G�DWH���\Te��ʹ���"��Hʜ�~��M,_�5�O��	�
�QD��Z��s�?�f莻g&V0��?�n�K.���KG�}yzz�I�O1V�q�?P���"��������q���֦iqM�&��6��KA���=�9p�U,�C;�����`z�h�0|�X���k?N�LY��79�X�:E�S%@�197�Ï=�����i"�k������ևX�O`��e�x��h��T���21�� �������G��,&S,���0�7�b�l%w���MK��	������o�o"�j]��-L%�%b����B��PYvњLB?�vN-`jzA��̩�Y�x��ޢ{O����^��*K�H4�d6I��`��&��KXX`K�R��f�i��'P۹�?�0Υ�X��[h_��{���wԧ���z~S<q
��:�T�نߡ��"�ѽT���D0hh��4�sq���Q���E�I���[�!�ctk\��9��j&9�0}�V(�T��n�-�5@�3yb!
v��n�B(9i�X1���wL��8�VU/T}�z����ʋќ��%��6'�U3�{�PE�gx�X9�淣���8k1Rb�����9nD�̿���(ұ�cI�!	�J5�
�{�܏��&�7��>��sfn�ݻW�D�C*�Aq��@lb��9�	�G����*������1����0����{K����"�; ]��]U8�4��R�s@�g�#7�0No�/\���.��CSZP��6�z��f��z4^*�ӛ�����B�\����d)��+0"mt�o�q�����c�R
tɕSǡ��`�r=�,���6�|'J��9!���"Ǆ�7�\����f���-�l	��+ oȴ�?�����N���tN�2.�2.�2&W_�B�R��=�@|{�ڵ�r�@�0-�c��i^&ࠁ</��KL��#n��*���!���8��	�������&������]}�ඩ
�$
D*�[Ul��ݿK�~�~���tC�T����(�P}�-\��D,����H�]��͞�\�!��`�)�1K�V�l�H�W�SĲ�vd��f��|j���=�*�S����fQ��J����G&�E:�D��u:�T��a�f�Gԫ�%���Ry����s�J-Ρ�Th�J���ٳ/��8f����}�cbjtS���^��_P~��?�vE�6�ص�K3�9�P��'��>�w�c�5���ϟ���Zj�I���O�n���5ܽ]�-w߫�v!�ʠ�"U+њ�9�Z�~���R��lĨ�Q"1�tܸ�0h�:_��E��ᘘ"�k3��*�Ĩ^��NA`�9�ڵk19���Z����`\Vd���y
�8�Zh�(���(�`\?��lQ�Q-�1�f��OD�]���I�$��"]��*F�O\ͼ(�m�+����q	��'�c%'�#�ޅMZj��N��W��vCF;jcY��޻��}�{�ԕJY=��ӆX:t��f6|� }�+8�����o�n�:5J��{`H-Q�5�E�A�%\*2���[���!��y�S��w$6��EW��)�YܘvA�Ȼ-l?�*$*|�Yb$�v�N��H�E���]�%��(�{}w|�x�̈k��(T��9B���w	���Ut�-�$��Ţ���c��C����o��sC����bi�X������ϒ�0"dB�\�}K*M��Ϲt�����ӧ�8|��Oh~}@�w0.�2.��,cr�.d��꿯��>T.�N��f��w��	k��r�0G"�k�2!?��t�+� _b¸��n5�$���t��2&�K��ō����h�G�A����5�۹�wޥ�L$�C�=/���Fן{Y5Pg��aߩ;T=�a��Z�������ѽvW5-�e��-w����ˀ��2[T�Z�!p�J�U" Je����
�Bۭ��	x/�rȤ�T��B��F)A}���z2�<+�׺��#�K�?��}w��l�[\�{�<�֕�ԥ�^�3}�_�����2���Ԋ�8�iva�*��d�*J?D���=S�z*�S���ǥڶ��Xص�K�������wi���;����j�N�{v�:�,�s�P>q�	�v��"����ιØ8�8��^�P�Ɂ9����M��Kqr^�g�����Mu��CB�t:���q=����&=,����@����Y�����g7Bq{�=��3���x�x�Y\��pW~r�m���<�y S���8 ��z�|`AZ&O���cw��s}�,����3�V��-��:��u�V�6�&�v'�ß}������~R�>�,8�Ξ={��N��3Y�:�x�kQ�?�h�%VB*F,X��$t��r�n����q��Y�ߤrP�+yw�=�{�X�Bk�CZ\����B��%��YK��f�k�����%�f���_�v6�nBj��+sO������ĺ�!.�����&c��	!�k���k9R����0��C��%�X�Ⓐ�����f(A1^[����eñ.�.��	���1�ʨ�򻃈U��o�9s�C�=A��t~�2.�2.�2&W_�B�E���DZ__�Ϲ`7��
-R�+̛�s�ny�5�7���yV\c �����`��,��p��` ��@<»���@^�81?T{� &�Ȩn�͚ތl+5����Ǳ��o�~���A���T���s#�6�O���#˸������u�2��)E�?n��n~TX^}zzJ���,l���j�}f���LB%�����bq�\!�~�W��M��kܷ�7��w�'�z:�U�D��mҧv���n����o#B6�'3귿�����gϿ��:M��-���CXX����D���dRػo�l�?��}��������ݵ��ss�O�A|�i�K�����S�vq/���E\z�,�"V<�űs�^�N'T4�Q[���ލV�v�zLȓD`�Ʉ�5ڡ����X�D��R&���j������P�"!b�a�`��
�`+�Q�sܒ�Hh �8+�cL�%�ce\�a����0?��ִK�7�,vd7�^7P`�>��p1H�ľf��&�l4�<M����-Q�%��Ȭ�C�h�!I��k`��0.������x���(�3�<���{��1���z("C.qä����|޻d�:#����K����,���9�����ENN�P��=ߵL�ZL�s����P��E,F�C���V�mRw��@ˉ�V��m����Z���N;B��J���``8��K0\K�vU+�I� dR>��o���G"��C۞���k���_��*)�l��0Ǥ#֯�����<Wa��7B�ԇ�J+�nb٢N懶'N|�o߾'h}�%3&V�2.��G)cr�,�`D	�-nnn�����׋��!����v���Ё2x=KV�C`��[,�u�qը��~���ͱ-����GM`��;��A��A'���q�D]�z���T��P�lJ �����)O}�4��W^�we�y��[��Q���Ga!�j��@<*�=���3s$�#�\q�
��Y�^�qA�7���� ����2���]��㱘J�>&Q"X�*�ճ��@{��c����B��J���o��D������$fn9�n��l%�5�ʅ�j���x�5,�ܻ�av~YibL,�����u:�T���^�¿z	"��s�9�G��Fti}�;*����?�W�]��#�\/c�w��l���$������X��E4���vMYF��$�ρ�x�Y���&��� A�;j����1�at~�[�V�D�5��r�Lf�b��4���W�UA�S��IR]&p������c-?\F<�LB^�̎�X���>+����5M���)ȷ��bq�im姍���Ș�Z�!J����`�����t��ͻcb���u�͈]�v���s����x��b���i3"�m-x�����X�G	�{�-�[�nG?�����q_Qk- �?"�!��\�ǡ۟X����� 򑶄 _,B@�Q��H;>�h��7=��;D�\둜?x�(��ɱ�}�%$�������ȭs�x;~n������Z�\r%�T#�ih��� Ro{/!��%V�x�בq��9"�B�>o����[�-sJ�錣�+p��=z_�:�6��'���o��:�e\�e\�HeL��`�m�J�ҷ	�~� ���bK��@@�۳��לP�)XX.@C�\l��n�[�	� �p�����f��N��n�.vq"y�&P�m+�~�e�P}D�d��)��u�k��΄��}&�>���~�WH|��r�����ҭa��i�RӘ���GKc�E�C�x3e��`]��3�e��D�E��[|c���&�(�'���^��"��I�Xe�u<U�*�IMD�� ������(�'ȶ=D*]��N�1ԛ�=;���yT��<����;D.|�+���_�j���P�_B/J���h�K��\AoLͩR��+�-��E�fE��/+&n�r��<���0��7��G���&i��e\��Z^�X�:�o9v\��T���s��'�A���v�h5� tzf'��`�F�X�&r9͉q�Տ�
�1-���H��LI�C^y���9K��Ջ�-���D�����RƉ<E%�ǆǈ�ϊy�L��+v=�q�q���&b��yQ����!�1���z#��}���jv=d7<#�:I�?l�l4����D;�V,ܧ��0�A��%|����c�=���9���Kx�78��޿����<�1��,���C uآ<Z�$�����V.����b<-`ݵ�|�5Ľ��;t]�k	�'����H�(q�O7�I�5b�"u#@�\����'�-C}�Zi���gR�p�u�ݰ�&��9.$Xε�>���|!��fqٓz��K�M���𜷖B%�r�K:G�{T�ct~:d�s�,�T�{*i��OA�v��Y��:�R6[�;i�>;�v���W���J�mc\�e\��X���Th���3�F�k����Jm���dy� rZi�}"��YՍ��U��e1�/Z �Bᅩ�.~!�� �K,y^�;���b�>�?D����}Z؉|�x)^K{�F�1u��q�G?K �US���6K�dY���:�,�F��!���	�VSї~�b����.��]w�?v��ԫm`���\�\e����z��J�4&2y��,��L�����]d3l�`���b�r�|����dH���t�������0���R�gܑD(�(�C"��n��c:e�v��%���tRy�wa��5� ����̋�����oe�]]�����ث
,X_m!�V�����g�7�py�:j�����_+&�Ln�wÂ~�<��S�ԇq�������k��Uqr���7����m��������9Q�Fc��:�2��@�����*��_����4���*����@�cIU�Vĥ���ؽg�I4��\�d\4g�f����R��z����ʤcR�V�Z��8]szz�x��JU��`�K�e*=��c&��荮�-�kt�͹��X���f��D��*�m�d���!�<2]Κ܋!β�1�n��t���AZ���4���%Si�~��H_w��X���Z�eb�R��.��v1��"��[�*B���}��o��|;v-����_D~r{��P^�&n��UH1���/�'��ۘ��2�q�[Ո�I��
b����7�@����������y��;��yH�½Gh=t��D-Q ���8�,�s;D ���)�{�I�@�7��z�3����ˊ�lu3�5[l}vlԎ,���i�XBYpܪ�1��ɵ��I#Ӡ�p}�D��Е�q�W(l"c>��8t���ߴ$W�k)��2%�p�>�17������hKU��H*7���-I_(��c72BwG.�Q�^�O\�J"�{��%Iǩ��Z[[���ϯ<x�o���6-��q�q���1���6ڻ[����[����&�N4j�/��[^�X�B�;��h32��.�w�}������Â(?=���HĂs�6Z�b�+q�1��tn���~_i���h�"rRi�ͫ�*�,҅�����Il��O#����k���6ZD�v-@r��Y�m��T��(n7�d6��T����h$�ˑS=bli#tX����tT<��*�M�6�Y��"J`�����L�$D�FANq�Rn_���D�u��d ṆE�e�i��w��"/�!�8�]�ށ������o�B��+�mU����m�p�4�]�u�S*�e�6�5]���U"E�[T{PHLK]{��=�"��}����x�mx�"R�[h���Dd�F�n��iLf1'�SZG�V�^���H]���d�Ƭ�����Չ�@�5:�^�F��R*����U*�Anz�T׫����Bt" ��{�		����&�˗/"�s��d�l9�n&)�=0�\���X�������3��lAS�h�*H�-��t[��%+C�7�Z��$��&�7D���	�=Cd`��r�e���[TTEm�]���' ޢq0ă'/��강6�T"I��G�R5�h�̈b%�[�rx衯�o}�˻��;���_�4��Ғ�'���Z2R��,�	�\k� C�J30^����8�t��xm�:P���Z�	y�	�?���z"bZH��[�h��8��1$C�ǜ/�3��x���Bo�Q��JlI����t�=.�B��o�b&!n̪3Na]6���FȣK�\78�O\!�Q+���u3���I����Z��}�q�t�F�%�Ⱦ����`��t����3��.)���W@��8K�L:�:)����)�����g��ziyy����]�q�q�S�1���Y��T*w���=�����x����3������C��qH	���-XНج��sK �J�;q�I��n�$�Xu�w? J�����`0��on���T1=?��wPˏL#��KO�B�w�A��U���Za�PKGe���Db�Jp�K���u���N�<�F��HrԬu�������U�*�"p��-¬F��ms#�����O�!`��*��&m�esm��^�Syu��!]��Tlh�h�L�����B�Q�Jo��6����/[�jߨ`��;T���
�zO��Q�[�$����Kj}c3^��RY_/M�U��=I���ޛ��Ͻ�Ū�Z�Z�ַ���	��8�,����bIjwqW�|���
�Dh���T��bR���	�N����#�����}di��Y-���-ݭ���P��]A���̮�,�����a---�P�V��׍�`��Ryv!d�'���6�.�V�݀VV*�p��ş��\�v�f�\e��u��f��!A���T��0.+ �D��>k4���l�g���uO2j~��Q)n��eE�L7ME�)j���ރ������[q�<'	�wT�5u��&t��㪲i6��>�C2��L����SF�Rp:�������u		,�""��q����>���
8�>&������%!x��K��!�)qU�xt��k(���%��q��M�;'�q�s��P_�����_y?���06��
�'�[�;~n_�ڞ?P��/w��~P�=m?��NW-P;����À��:�Z)��ƃk���g�xE��J� �!Sɮ��o&V���Jj�?��ו��w=�omm��i9r�'����L�kcb5.�2.�2&W_����*�n�=���~{��H2xeB�Z��Ǹ�'��)v1�!���@:V� ��Qp"��n��\G�Lsak��%39t�"�I:3��X	��v���~U�OS�L�!Un�������[���>����u����ձc_F���ziEum���j	�E��i��ڪ�4���x"��_&�E��|Gy��H�E���������T���Wx�6q;lRNC���)�D�#S��>}�#U��B~i��I"X]�c]L.�`���Ãlq!����_A���x����FI�����{�Sɂ� �RI�L��I5�+�¹���rq����*�c
���JJa���vϫb�ǵ�7��;�>�jp��E�Q�gW?��q��X^ZFIŰve�R&R��y}]k5{f"��Rxjڸ��Y��zu�f[�Ryd�9Uo6$I�0�v1Yb`$1V,䰰�`�K,9�d����<&拭<d�X���%;j{{[��,&[&.G��KQ \�3$���d�H�9ƿ����oc��%��,[$[�6#M&*�N��^����������U���M̓�XŌ<{�P�[n9������֗��^�bя����i�E7ϓ�{H~}���	 ��5e��k��JNLU�.��Q�S���b	*�$�ťl�����$��x�j'�nn����X�+��h��1���b=q�IQ1Յ'&�/m���iG��������1Q���+���9�l�=���{:��9!mtc�����<V2��$��]7�1�u�B;�C�z�`�r�KYb�O�����K��1 �f,��@�{׮]c��։'X�'''C��0.�2.��'*cr�',�b5�h7����zlmu���d��`���11�F���や���+x��*�e\�2���E ��Lk=�l��U��o	��S���Z�cv\=K~,�*CmJ�Z��jjt��X�QLM���w��|vBت��'�G����r��������^Ź���]��j�]��1��g�L*�n��/F����t*��~L%����Y�R� �"f�nooask��"�h�o���&�W�~W�P����X�Z]��.^��g�m�%�49���F���MaǗ��}��&N�>���P�����x��Ѫ6��_~����<�Qİ�J"�ő$n}e��l{k�U�צ�w�A](,���q`9�G��D�jϞ��JKMV	�|�VJ�r�<*w܆�Ew��K�Ԟ�PHm�H*���Ḍ9�Q�49f�~1�VQ"^��қ�M���A�N�О�Ȥ3����&&��N�� [vܘ�e�B���\�A�7��iks���s�5� �Y�R�<��K��	��y��5�?�c��4su$������X�4feD!f,JaI������ϑq?4;�bI�ƛ̸�FL<�!��LR�fKG�ں5�,H�Q(<u��˿�+<���F 䩧~���5>|؈X��� +,��oL�⒀����8�l��w��:����A��w��=�b�	�l}��
{a�)�b�
�eF@�$�%����|�17B���ɣ����v'd���]oĺ�J���<��yW�V�:0		�H��ׅ�jټr,bC	��q���׷b�ה����P�nyN��k1�y�>�S�����y���
i�}��U0��r����5WIo����[#ߋ۾G���7��bE�ޑ#G~u���'�Xq��V�_�2.�2.�2&W���nln>B��Z��|"V=���re����E;p��"���sw�rx�O�q	��".$n0���UJ���t�	o��]�y!��c�]YPB��"R�k�gr`1��!Ad���uՏ��X��Y����Uv"�����x��/�j���rf3_y������U�fU�z�=t�-"*ң��C&��t&�-�Y*��U���(��F�=e��Hc�LI1b\��3xZSŢj��֯]ǎݻ�c��'�P�9#�1��K�D�2�s8��3Pk%l��E��7Yc������@�=���Ebؽ<���>�r�v�}ܐ�'UwY!W��lf_��^Ly9����>��П\@��1_�2���DT�\�76��S�a��2��@�]�6�H�������ɡS���vS��x�F���c���1�R�[��X����Vr�qg�?�T��[pr���}����P�.�S�&΢J(��H@l�9+Jr&�G��&�6���ka�nD�?��!�����2q]ĸ{,z	���j��<iM��Fˤ�1d�� dW���(��W�����^�O�T�W��~�!�ݿ��O��[ob�}��������@��'$�.��j���Q���[ÆU�B뀓H���-SfL����f���r�Ur��-���l:�C����EO�)BV̼��������I����H���O��nV��y�ڱ�k�oP�$v��&�����{Y�Ī;4�{��I�]�%�Jb��y���Т�#��0�!�j� 5�&�1cm��ϋ��xI0n��]-���W�pn3��3��;��6����߿�w�ԩ��=�/tXeL��e\��O]���OP��4-*w�������+G	�%�f~�Y�@pv*��� �B��*������k��j3�Z�����E	�c�,A�{$��V�:t�x�#.�V^ې�f�����q�KxRT_����7	�G<���ַ�8ߨ��K�j���R���T�w�C��w���J�ڙ<}L��Sg�J-4��(WT���Q�O%17=��X�nY�;A�W^��\��x.��Z��Qń��"��H��f�o�>5�:�Ϫ��)v�S�F�H�B�ZC_~�#�v��N��ɣ�����cg�X��}�����g��+/#�<����~�UW��"���#���c�	՜�k"�&�r(��{J5�/\ץRS-.,#��P���OǗ���'�GO?��g�<a��f�sq�G1Gf2��Ss�<]_���NWg#1�I�Q�vT+F�7�1m�}�afbJǒiUe%�Z�X�44��0\����m۶m۶m۶m۶m۶�w����;c�/\��ɬ<��!K�L�z����L��>½��	�j��ቻ_��*m�ğG��*i3�sJ���tm��	�oxM�}έI�%���8�"��&�2u�}R͛��׬^G���5&q��W�5�0'V��B�r�Q�d~�� �޹Gj�����|�${��7�����o�OFZ7l�����ᨒ0������`����a3B�(1"`( s�$���1�C�gIk����H� %j�s���"%(,&e�w)0� �*鐞����$;^��Y�"K�{��ǒ���!sM��E"������l!R�tz���%(�`��/�m՗������k�?��PD�CԎ���b;�q<X���wt�W%��<򐩦�������E��9����J�"�w�\d~���E����!i�ո�����*�%fr5���B�ӡ���Z����ؘxz��c<����;�гZ�L{K�AjGk��ԑ,�S]���~ǓD{�Τ�����(�& �>򠝻x��3��� ��^ĩ&&�l�%��)AnD��_�}5v���F�����s��eU<_7p�1>���	��\�p������\�ڽ�}$�~?t�͵ˬt_9���(_�=Z���|��5��Hd�c�.�	��3��/NQ��ِ�;���o�L��T�*Oe��q�������3UAw����������������c<2xu���7O̯M��j1~_����>���~ѳ&�\��K�Xn]kb^��|eM|��u
�6�J)ݚ��(p�,ݜ�߁O/K������i�{�Nw�R�7�j�D��9
��-�li�������
��m��(�X�5F*?އ��iE}{kC6!3�e���:�wd��}����ų������|�[�����LS����P��UQ�R�Ϋ{�1�ǝ��n���קϞN�q��jʧ�Ǔ3�a��Y�Q��C�n�^�v��ƒ���b�Z��������L��r
�5���z��k��՗������i�A �8ry<�;X��2��k%�-��n��w�s�_a�.�����F�vG]��7��4X���b�臿���F�W�Ddq��� -ĉyI�X��֌N�[��>������8H�h�
�"XW��1�ح!�t>oY��HOLV�N��uS;t��֩�aNu���0(���lt2o&}R�%��C�&���Ў�i��"p[��C�]ֹ.����n��A��".bc�P0�7��Z�l����~>�j9q�_o����/|"�0�5c�z���w.1JR<j��S�Zŕ� c^�5t�t�sN���Jrױ�BwtHq�QBC����_	G7us��q&y�M��7ߑ��Fւ� `�Ӫ���c'7:]�k+ 1��[�*���)��3q�Um���)_x4�ؠ"�Jީ�v���b/��[�?�U�W�i�WD�=��^A����&S�eM$Mj�n((k���z%�Z�F�n�P��Li���aڒM���3I��# � ���2�.�#صmI̜�V�+�0W2c��$
dfv�8�����㾒j��s�v������uv��+�.a���x�����lI�/������٦��MKTψ1M��'b[=S�L����o��wn-N�6�cHK;s8g����$�7��M�_��n��zk|��(R�m�+���<A�,aF�@�V�%un������-R��*�%�q�� o�8-K���P��R�=�?���ќ�!�Hy�hfD:�94j�s��.Ӵ6d�c�*C�J��T���F�d[��� *�rc��f]�4�¹�-��O��v}��#������*!3u<?�����O��#�.|��l��Þ���� ����ِ��;�<�5����_s:���Q'ɝ�����ҹT�Fp��勆����p��8��Z�WĎ��C�&]��ʤ��
�O>�=J�ftt6�D8��c&v���(o������ꬫ�[�=Cf:!����5�{��RO��ml��1�U>1ȸ�x��po^�7���ZJk_�{��:J����N��z��tbϳ8����(��t�8WZ��דOLǗd��襸':�s"(˰,���`�1���p��ې;?�Ѫ� ��i}V����C�%W��ey~��������t^�%�vK��۴C+�g*�U,RǋGo�,�����w�h���D��H0G�,�^��CG�����'ј�5�yQI�`�gC���2Eo��8�>�]Ͽ�������׎��?�_"����ѓ,�?|P��"�-ٳ�4m��T���>����
��▃t'����4H�T=e򹢘?S������ u�~i�ȵ^���g(o�z���h�\��P� �A�@Cѿ,���"]���Y���|���`���DR3��a�+��x��T�� Y���]P�Г������l��
����p�^�<����}a~��á|��־Hf��}��0�O�tNw�꜒眽rz���A*�V������l���+N/(@�'TcY�V7}�7|�,L�����3�*q����\o��u�dn�?��$�طv[�9�Xڴ�E���hj܄*l6n$]%�w%��D�֊*�PN� u�Î��!s!g=j��z}����H���XG�����6n�*3�ڄ��(L�aI���I��+n���G�r%F4�z�.	��@𢡄U e���D��N�$nw/������,��Vi�������Rg��T�0�<����_����w<��=D���<�wN�x#�e�!{ga��!XBbDq�9�0�"fk\�m�u,�n��픖tڎxޟ�ژ���n�0a��v�ԓ�$/�F4v!)2�$Bu8/J��!>�t�HԎ��p���t|�{^8�J�{�Hm�1��t�Z��}ؗ�D��m�]��|G��~��(�pc�Mr�E�{����d�m~ï�eO��1�y�K8�,R:�k���P�._
�s�]���ѕ�C�@�{Tkܣ�O_�|,���UU����������\.��������H�����I*=1�����:������n��88� )F�M2��=�p���A�|�u����������!���"p�	��d4utSm1i��縅�$��xB�)=mג]eM�A\e�3��h�G5�J�#���j�Tj�(#k�XҢUoX��b�-UOx��mg�t���r��6�ʪ��'���p��ʂ�l���uVD$�˷e�*M�d�Q '�t��,�Y�li��V� �U3|��J�ʈ��z���U��,����[�zo4��KA3w����S�[=��24'J��lAzL�|� ���8Rd�;9���}�{-�W�g�xA�p%�^��1*vNuU�e���Q��$JJ_�`��zv������JT�-�;V��?`B������)��N��~G^U|tQ�b%�|qV|A��%�L+	B�Fpt��b.K�	!!ۿ=���z��łجA�x���ǈa�ީ�N�9��#�3��g�+P	U�󅬑�Il@���V �pL�QG��D����1fp�S	N�DfPW�H��2�`mP��8ꤩZ��Lתݨz_c]L�)�9�S-��I�}�}���u��о������%���x��ئ�xoN�3�D�h���G�*?�rlv=ַ����IX�JA>�t]�Sv��Y��)G� ���%&�9n��x:fڨ�3�ˮ"Y����㿌#��W}��}��JI��DI��U�ۢ>��%�M�d4�,�s-f\�B �D��D����!DE~7��/���EbE�7�v�@�2=p�2�;���]�+-�D�m���*:ޅ��/m��5%�Sf.�)2H�
)A�DZo02v��}F�>����x����r���~�o����ۥ���a��?�����Z9Wl���z���+U��#�k*{���1�B�$�񅡝WF�9�M$�f��/�l;�'���R"	��|��' ��f��6Tc1���H�#�;~H�Hrf��q�Z&w@��=W�p��C)gdd��ZK�<�u^���8݊#_\�[J��������+Ep����7~-z�R�/ڳ\���w��Z�*W(�V��!!��{A�n�gu��L��DF��:�a���/	�$H�m]�%D��qŒ$���ߨ豲"�uّ%�1-Ѩ)خ76#V�k�i�}�B_����<�<�ې%I��� ?vD�:'r�u���j��,���eɢ=p�-G��P�Χ�\�M}�f\U�}6�*{���,"��w������N�����n	_-�[��nR����o\-]��Q��,{��O�7��D��,0������*�IN�L�,7p_m
A��c �;�V���Cu�m����Î�[�(R8����4.�N�׈FՈ��5y�S)cQ#��H=�H�]i�h�Bz���F�u�F2}�U�E�Uh�����v˻rm�,���J�D*ky�DVڶ�zEy�}sx>���r���^�Ӏ�2��a�:���"H'zڭ��4VE����.��"e)�w�
�o��;�k�
Y'�ґ��i���7�q�c|y����h��U-1/�e�	��'����.~s��~G�Z^y%�O��X��#5��٭c�k�}���^�Q`s/��ϭ'�Kǥ>�Z/%D�o�߿�R�6�mq��kݘ�������r��$�
��oV��W��2sJ�#(/�7Y�#���S�{�R�O�����t��/��9k��������g��4�n��6vv<R�#x����d�4cA�1��(Ҩ�=;��	��<H<"5&��R���a�+wuGXQ�@d}�8��U��8x�&"�6��qI�dB��m\���&�)���lX�X���D(��b�֧�$ǖD̐&I ]ڨ6�u������+��������_g����k�N��w�З���2�b.-�O i]��M	r؀!
mc�0��ѫ��A�Y��0�(X�&l�^4��Q�ˁ?��Cc_6a"y[
�vG_�����v�����쏃��W�+![�I����x;�����ں�O�+�_ �u�����c�V�;Z�Xq{�B��^Q*��Ɉ�ɖ+��ػd<U�a5����_��Ӏ3{^(�����������7�磮��qG d�*/n�Ū=��;���P-�bC�C'�Z#�Z�{^X8��8KC|<��q�c231jRU��шv�ĥ{�f��{Y�Pv�at�s��~��V30�aN���0ygd�Î)�'��)���` lq][W֭�"�ԭ���P��'���L�By{*ʽ~�������]����}��nmq�{��O��<�D&�dB����="���Ar�%*�O�s��׌r@F:�)�I���}�V+~�-B���L�]��N,�H���#�l0��1q�Wߔ���AZ�OT�01�{]�x�"aӂ�΁�DFg׆���ǩ�Ѱ�y���&D#>�;v�5S�G,IpO\�\ɺ����|w��6*.8�a��s������i����t?o��=Z��,;_ר�	��K�!�3�P��*L(y��������4;������3sr~Bs�_eh��t��Ӎ��T�[b�~�����Y`�N���v�D���D1���rG&F����m���!�QP�6���U>��A#�F�b+R���l��z�P\�H=GzDOӾ�VA$�gƢ�SO�T��5�H�ShЗ��X[U+��W"�
 ��Ȟ�S��Io�b��}�4/C�P����x?�QdǞ�i�ӛ��z���Y[����p����v�ܩJ����Bm�b�	�0j��MT�m��5��NY�I����8�!����e~-�Z,�x�ߤ2k����K�������XOV�\��d���w}�]0���d�y���QW�w<ח�x�,��΍���m�:����#_���nǟ��fg�6/�U����#�D�I��/�%	��#s��8����;���뿰�IK��Kz�.���%��?@"uU�foARrh��'o�����u1�%�J-��-!���4D��cR������F�O��r)��@I�c��}���T#��E�-�g\h�G����Zܬ�)(�����W���^pm����-6�J��t�[���Ϭ���	�f�?��Qx��́\���~�Κ��9���䯥S髁@`���p�!�1Z�)_���n�7�nc��� �xW>|8���G>�ݣ��o<g�>E�Ԇ��T�#R5�t���;V�lu#w���{Hҝ��uR8GE8Þ�T[���޴i��!���c��n�q���cH�#�H�I��JD.��wd=␕	g�}����k�H�����K�5�N��
k�{L٘��R*V�ٮ+�ֻ/�^�$��ak2�S���{���yyYY_����_M���©�d�|=��������AΎa�q���`�g�w�>)C�a�g�!Pl����	e��FO����k<{�2���КX�/�B>�&�h�����6I�������>�Pq
�P��T~Z !�d�EФh�"�����$MH�'��?DD)jG��BČ��hf������^oO�Cy�:a����q~�IM�i�r��+E�HٛzW�[:�HX 6���@Z��
YG�?�ߖ5Z(�������e
�U�M2h�9UE��"yy1����[�g��{�S��;Qv9�����@��\%�I�؉����7t�;�/|ߪ���;^���~�6E�q�x�f����y�R|��h�����ШF�� ��7B�R�;�)/~��*q��/���w�J�8�J�/X  ��p�)_Sٵ~4O����t�=�vDQ�{qr��W��<!#ܒJ���t�Ay'�}4��q0�Ve��<�c>a#Q�(s��>���z��@���9u�E�؏�{�`���	�	p9
�aՈ)Ѫ���0[Ϲү_��"��l�{�Ec�r��5���W���{��c�����1����t}�P��m�?�Zm�+�sh�+g�G����u�ǎq�t��7�+���Ͼ����V� <]�k�Qe�����o�{���*%B�d�H�{�j��uD��ld��0�c"O#YLr��5r���3�)�U*��T6�!�:��s!D��Q��G�GWBd׽���6�WO�����8��5��<������'�C.�t�2��O:\�@5O���b�s�FM���66S#��k���?���E�N�s�1u2�L^��zm�2g�A�����zT�p�\��}��ni�9�j��֜��)N�� ��3#��	��L�I���6��
��nb�
\>�>A3 ���,wA�
K�ʲ���0q��X�8��Yy��Ռ�y��|m��bY��b�Tǔ�,!V�
�^ߥ�r���*�(��.KR	�,B��f��eF�7��p�o`�I���x�,o����Ş�wղu�g��t�L�(������
�~����(x�A�ǦͱQ5A�6���n��Zu��qd\�1�D#Yk�O����k�L�_I����XT��6{3p����-������z��l�"B������Zvۍ��%w��D>��Ӥ]]-��?p卋�3��Dg�z�̬m��B�QY��YIb����[��WF��Wl�q�[������L�?�%��u��aS�ʿ��)���Lj�-^r�|�h�eJ�����s�� �C����DZ�T\@�GN��O7���q�gLx�D[���EN8��MVBY����kXۧ�fl��6���K��ш�}Z�dE�Oƃ"�=�~�kX�$0th�U��E���#��v�W���9��8��?>�����{���5k���g��%кI�\�{�u�&��mz/Sp&]�ܘ������.Ǝ-��b!��:Q8�$���^�N������3�{��?���O�H�����*���Kh6 � �ݫ�~�������d��Ǿ�I��`�VL�11�=�{�~Wz��E׉��6�Y��񢝹�A\���5U��%�  ��f�0�u5y�%U+4��}g?�c�s"�d����`^&�@�,�XX���r,|���-»id�Q��u�6)7^eP�g�0(ʖ\Ra��W���V��z�#.�Lb��ț��>[�	���l��!F���T6,�D�y���Q똧��$"�e��?o$"�jzn�u�%q��{��j�}��MJtܭ���zI��v�~�����J[��O��L���Ӿ��wX�^仜�Oo��w�~�r��5����Z�(�alCh��$�)�+ ĔbR�I-;u�Im"R�󀻅p���Ӓ����=:&�G�M0�<�w�s����܋�E�+���(��K�2�Ǉ����U�����G�$�V�A~e#�� `{���o_�i����8RՖ���­�mg@�N(���I3����� Y(���'����^M�p
Ƴg5�R�0茭'���!�JD��]�W!D]Q�#w ��������B>W�Ia�䙁���]
�B�C
���M�H��.�Y� ����b�`,{=�NEz�.rZ+��2H� Ֆ�����5{��7��>?��t�{l�Я꛿J�7���%Db�����*-4���$y`ʓ	py&:.-�:1�5�T���6m�������?y5a�xy��|�nس�X�n?�Vzj����]�&�9����4SQ2�t-�����k�Y7A ����*_b��Kf��6�Γ(3J8�Z��遵�4�T�v���>ЩK������2���^%�'�X/G?��V����j�v��8mZhLjR,����?X��m������^��-�Z�`�4VNnȀ=QZ��A�����H�e�l��q�����c��I�s����ʾ����9��흿�_��$�;1}��C��g���h2Jt��e�>d$aY�3�j�ͳ ��Ti����$`rG�+a�O9�
f��$�oQH��r�-�cM�G�Y>��v�(���P����~� ��Õ�Q=%-�����?�WzSУ ����J��ZE��W`NBG�Ye1�1ܐ��B.+lT���O����c΃��X�)����y�a�M�uM�?1�ԋ߄��d_��cn���p�9s��b���֎t�~R�!��Ō�+���D>@�yBZsϦE
����	yY�<q,��lI��� d�HjY.�`������ ���M%m$�f�� 6qtT�������Η.W�2��5P��U��-���M'B��[���Ի��cl�\�UIJ�?㏙�宻$�y�Qi���_@�����7,켾��bWP�$�݂��5�8�c>��V6�	�ZW!�@��R�d	;$��n�b�r.4��:&Xp'�.RP:B���c���삼`�j�ۇ��!��R�HQ��s"�ȍ��BA�o͆9Hs�$�!�N��#�0����?�J��S��<��<����NL�`�jګ�>��%������iY��V4j��4�S�n�BBk��,NpZ�#1%1r.����(K�?Mi^�EV	D��#h֩�L��+F���G�����I@�����E���L�P�:0ʘ��Y��	�Ѽ��}�^�g�������?�]
v��f��ɘ `=���ܠD;4�E��`|��Z]��}�,�x>R�Ǟm�Y�J���Wu�n�Z-�m����M���.h��9��8Kچ�C__3l�|<t͡@��P�����Rv�`)�\��i��D��K�8����؁Vi�3� ��n�
vg�o�`�غ��ҏ�׼X1)V��G��
�ỏ��r�)@,�;��;03C�)�K��y���zg����]�WY�(C�f��
$�TdPya�)���������h�q��~M�O&6f�d����V�ģp����ǥ�?-@��kݳ&���K�_ޯ��/���P���R���0�T���ಶ�s{���⺑����S\q�e��B��ϗc�	�_�;��o�S�@�J6�f* 1�~������_�M7�F��L���2�?���HY֣	/��wĒ9�`ݹ�W�L{�zx>��l�ڟ�v��PE^��Q�_��B8����|)��T���h�*D���G�k ]�����M*�Vl�1' �o�u��?��o^�����l/7�7MPm;��/G����Z
_�Wl*�V������X���-�"���,2�%�M
��ֹۭٵ|Q���B��]uY��� ����y�l�t��*�X��PH􇄨	�Vm�Ho�e���P Ŗ�+Q+ErK箾9M�	5�r��Ĕ@���A�Vzz�j�+Q��z�Bݹ����k�
Ab�T1�Ԕ�,��
u5���}j9��$����K��Zi��O�	M�DSË�pÎ��X)՚:ۀ�	6r�ǜ�o�
�X��[$D�]��<F}v�Q,��+�<4����r�C��į୒�*�i��^0mVVR��0�O��s��`KF��y�%S���'����ワG�/!ύ@���`̱�AADZ��t3ND٢�>1��)�Z����F�:�I��O�>~��(MfXp|^q X9���OwL9�JG�p�����Wi�������P;��q:b�2�C��@�䖒l�"pFLx��(-��p�w�!m���{��DP���O�(	�@��P�E��U���t��U��G���ZT� H"��W�0�n�V�Y������px�4�d�"������&L��0�����~ԏn>�.XR��r%���&	Dv��ı��yA�}�������0^:�C#::k,|�����*]�,*�����.��;M�T]te������	� U�40�K���>i�!�3\:�&�� ����X���ϥ��_r!y`0N���Z�N��.�v]�,!4]����&/�#�����u����g����.�4���۴��3.S���{�x��g�2_Y�$S2�")�HuE��}e
��FVt;�>��v������}�Uo(Y�񩪫H��& _�Bպ�eV���%���ӧ�5P������n��MLN8y|Z�k�Sϯ��ʗ�U��xT j���-;��]
;����`qn���1�Z��s��_{����Xx��tQ._�t�9��+)�S��P}��"�5�z��ʚ
q�$����APT ��X9�q���*�JN��;��t��l -�Q��6�˒���J$��&]�&��:%u�R���6I����ɿ#̄G���>�Sj�C�{W�5�<IǃCp>dt\j�BH�Ū6�j�ĸ�!5�$*w��"\-�1`��~��� �UƗ�P�j�}��u���-	����Z��ְ���K�{<sK�����z6+��FB	�ہ���o�&5��S}ÇR�.�n�~`����q�^g9��W�7<8��}%�H����;�çU���%�"�ve<n7���1e����=�?�kj�hck�Z���dk��`�{;Ny�E;��)�!�Ec$�l�����Ǐ�u�T`	�e�(lm��ڭA�n�V/U������ E"��z�N�gc�^�Ϧ�8/�@�J���j����8Ǔ`.8��VU�����h)Oh;�]��u���	3GO>������E�O��3��n�TX)�#��A��V�E"C�/}�/��^�og��H���|���h���J�މj�e�6�����6	P_q*��6��нl;+��"�������X^�4Id�-�R^��F���"D�U�.A��sBH���9���y�҆A  � �y}��O�"��Oހ�hX��@����M?=0z���o;���2�*���F�2�_]��AE��8�m1�"m��"��_O�#��g 5;w��=,�^��dĎ#GS�n��$�ey�h���m�k����F�-ⰰ0�,������WWl�Urhh�}|\\_H�~)]��%���_����`��Q����M��c<�8-�A؉ۓ�����x�՚��Z�s;`��k;��@X�:1�*�,��em=q	��=�3"Ŧ+I���aI.�b}1.�J�o���&����X�H'Y�׫]�;/JHH�XqN] ����V1A���%d5~R����"�x���d���
/�i�X[�o]��!�^Ɉ��X�`��Į]U�(�<^��B+4;��Be˰�o�֭B����HJ�Q}Wâ $���K��&�}D�E�W L�"%���P�*�-��͎0�y9gfp������kr� n(�Q�b0% �Ll4��	�����xt��h!j�Ο$X��zrm%���O(���­����^�<LmY����������0��I� ?�;��p�;`����J��F�����l�p1����uЭ�KG�ђ�7b�S~Dtp�*��Y2e	����S���^ò��s h.�dCC�8��&���0������릑|4y��;-g����OM-�ti	V��v*}>�Z�n��oy8nx�X�0�d�#����� i3���y�;��'챣���BlD0��)�h�G�?��I����c�?8u����B�&E#�Aeɳ�f!�F Z�xz��Q��u@d̿�|l��0k�� ^��85&��M_��: ֯и�(�t0��?�,�ڋ�\F���,R*Xt����#q`�Gy�Y��"��4�}�Q���g�w���̃)j����A |a�lU��W���J7+i]��$�.�c�5� v�l�'F���O����<�<U>�W�$cW��r� 	��3n�:CE�0,�&#Ö�	�P	UGWוY�f)08܏��ٙj{�A/���M�h�����Q`j-��b���t�o�r$:HgDca�Sd�&ڀT]V 3�w;Obm��Plh�}��|`\`h=	e�N�颀��U��'�IO<�eO迵=Z�q��YY��UФ�m�Z��.x�(�g\е"e�TIx��c6JW�a�\��;K�R��dk�B���d����T�at��p�ӣ�|�����ZMp���N���V(XE�NJ�K�IP�,eҫ�Lc�|�$4������Tź�@�BH�@°�>�<��_1��N�tE��3�b]��$�|8�(83����{I�|��\���s����#kj�K�$0<O )����m6���4u<�՟̪���q�ٹB a{ȀL��m����!����t�&�)�_��M��"���o�B�l*��uB;-�E�����D;vT�G�	�f��E�"b�B%��%�Y�f�K��7����֮B-,�bB���x8���Ŕ;w�		Z7	��H°�4�~1$ ���)���#13?̨�l.7lVI����~?��H�d����GAgS7|[���oG�����7�牒��!�HUʧ�?υ�����m�y:��h�E5'5b���������TY���nO;��3�?�ݞ�����H	�<N�@���
�)��E��2'[~Y�9�`x�GeO�ȫ��w� m`}�QeA:�G�ʦa*�NU�$6- ]�T�H2<�^(7�Wk;��e,�E? �F�qI�;i�Y�c�Ŋ|�'����uz��]������8��������&x��衜Wf�9I��m��Z�|��3Ѹ�#�`5w�~Ł����v%bYɷ���}�+�h��Pgg��ז�k�����c7˿Щ|�JC�W�1���ګ�%#]t�kk����'R�����PK���d��?;̨��E��'��?RG����إ��lm}=�;(�O��QA�����Z0��y���yE���46�Z4ߣ;������Dh?��]qTW<eu��L7U���*��
<�\"���ڲ�
�$�N=*���Vs���HrU�qG�T!_z�6�O= (�Ew�?�Ҳz����:��Ȕ�BF��R��8O�@'�DnBFN0������L����;�����OT;��"�.#���~Y�JIƋ"­t)�T����J�HMf�C�o		��9}�Z�2��2�&��=/�:u��OvRk\
+�W�O9	$�7q����
<^[��������Y �D	L"� ��? nd R���J��`��E�����녎pR�fogL 8����̠�n��p'"9FvAV�hϊ��?���en���Q�?�:���
��.A;.9�K��dх���P��ȇѾ�{4���a�'=�z���rP�M
#|�
��J�լʽ��A��v�\�p���3�����h�]�{~>�飘���|�5�2�گ>h��z�����ූfI9�all�
%����n�B��Jhbc�N>8nr��ޚ�7��o����>_���s8��x���s��%q�݀w@�J3�LIb*a�yx���F��K�!a���Z#�= �8H�D���]gc����*��4���1�E�l�����(�>-�!R��*ⶴA���ח��C��8�]��7���u�����E�����R��:׿��u����t]f���vk�y9�f����@�of[�7Ϳ4/c;�tԿ��������3�,��K��[��\�V�ܸ/���!T�e���=0?���J�.^p�@���\�b����������9I�^��t�����RmZ������;]�$T�ULn������os"���ȳ�|E��J�;n&	�(O{��������� l@(�Ä
.2��Z��Ej`RcG�J�-P���=j a}nė�6'B�z�ZѣD
8�
�O1�U*TW�ֈ�R�FU��(��R"2Q>�R�P�,&���
��L����wF��(7�r:�ڞ�XP�	XXA��*x�:���_��H�}_l@8�`7(<�	�("�QaJN��r8�؁�pXg'J������p�E����Hu|%nʄ�����>���E|��u"Xۍ�N@y^?�n�X:\ވb�c�����#G
�:HM�H@܀���&�^�#�������*�L����N�+��#�m5��l���4�r�'C���a;=/l�W��G���P�n�B����A_����-�_�!��?b�|q��o؁W1�X�&��,�0^I5h�f�Z�xhv���8�t�� £)ف=h�>z�f0�E�76�I����??�,���=�jhd����~�ˏl����������Cu#8��}�����J~p7:FD
�5؇���.e����D�ۭۍ�Y��9���%J��2O�里�^?�����\g�f�����?�e��7tr�
�GJ&$�W'�+��a(Y+k�]��f5�~C&���
^�m,�F���P`�bY�G� :e%R�	bhW�i�w��Wa��El���3S��iI���eV�D���h���g���.փ�4����g/�3��� �5�*�=q���U߅ u��\����Q2�z�}���Wܫ���מ!�yxZ�0�GЍ>�n���'�`�̅I��w���i�A��S�KcU��$�~� ��C�v=x��	���y故m��#y�{<������ӗ�B�1|��"��2m�x\M��`�G���2p��o�p#т"J��,)4_**�8�`(n�2涭a"�y�@м�\T���eI�UA�cm�p�!����4]'��L�襬c���s\��JD:����*IǍ�R׶��悫�ᚤ���A�aGUR�A�<k�ʡi�@$�&Y�,����󟨃4�a���(�'�"�{���E�o��y@�а�4CA��ݖiЧ-���<G���Tfʝ�p"�����?-���%�)j��[pr ;��Ú#"�8�5殢�QQ�,^��"Vj-�R�e�P�ø�R&��z��4��<3��U���c<�x���IU�ls��&66���q��2e?M4�@���k�(�����%j��W�C"��{�-�X�^w�(9;^�8X"�Mi#E��R�nA�ຬ��4ЯQ;<ˬN�5b���'��焭�{�?��{Q^Գ��K�a����,�Ř*��DKQ�lj,E�)gjp��#N1pK��@t !d�F[�[�z
h덫Y�JzmCɭ ��{����K� �/8LM��������az�������7ڢ�Z�@�XV�WLezacg7�l&���$��]]�l�`m���d)�#`'���H)���(�J���:�~�������'�9��XPB���m,<�j-L�* ��x�"]��W��b)�х�픱>�����懆׎���HoDSWp��r�����֥�!��<�O�������j�`�8'�ub۶�4vN۶m�j�ƶ��f�����w�����g�^kf�Lj�����2��e�A���3Ӛz�p�l{;��i�+ ��X����� �-�7��Hz��>�|�]TX��q�o�G�[p3qQ�J�´��`��%ȓ]�)�Y�Y]�Aʙr)B�O�A����SdF��ҧѻ�鄇���E�>}��39)��.�JI0\# ��Q?�ޏ�]��{
���v���V����x9�R���˚�'��<�XH�������/,r׊��*������ �s���yr'a������b��oֽ8�5[��V�z���;B���Y��yR�N��[`&��CS�[Df�I/�Q0Vo��j�Ǩ��&�S&��C��y�뒍�g��.X����O�p����2��bX�%��ׁQ.�q�輐�M�����=�L��ڠ2���֊��hx�&¼^��>���>>`����]�%_�8�^Tϧg�xY�W�#�#�Gx�n�g�)�^����Z��D�B7��~�&I�B"�������X���>�ӡeD��q���Y��!��:�6űvx��1���!��KNі�@#��?�Ǆ1���#�6)�
3�h�[�eu�K�h8�/�W|�����u~�F��30P����s&��e��̺՜;R��}�!@|�^��C7RS�bd�r��]�@��$u�]V��k��Ef�*�{V�J4ͶK�
�uA�(d3)��[=>�>����Q`n�AZ�7�٘�jL��A0zxrzz�v~HB_0^��&���;!.mj�=A2��?5�������8�#"H�|�����}<���������N���:Fy�Z��K"�9:�~<9i���hu��"4�]j��=�$�#n-�Wc�b�_(-[[�<�hh�W3��C�����Y�;�疿��o}|�)8�R[�]�;Ka�x�}p��w�]�
��f/�0I�5����4�u�ӂ�2�'繁���_��k�xT�q�^l��/L&$�/2��0,�4���N
8����0��[HT*7O���KK��`��_O��/�%��8�*TX`�����ZaX{��^��P?�ϗ.����4ǟ��J�b����ٛn頱��dN��[
��G����A���#	�#[�o�g�%�gT|����q��t�p�sL�z�cZ5~L��~;���4��H>S�����P�@d[[o3�u6����lMH�3Y4N�9}���-��Z��e	8;}���|��G]��uTukI��4����๩��"n�t��!~#e�����\#(��i� ��)�C�b4K��i,TL>_��G�"�̏�I�&�� U�h�J�~��"*\o������|.x�����4�8�&��W'�;���E���������3�^�Ĩ�E$+	I�/�ǆ�`!�f͑=�^٣CXY�/N^��c%>�\��7)D�-J&K�
JH�%\�C��@�f6
���yj9���%�F�F���_�}P�`|�	22L�jf��]ۉ�	!�_UD�i�U����_�HsĴ8~��ߤI�MqY�W�c��?���݅,���;o�XD5�Qm��'P�b�v�H��/Ppa�I����B��LO�.T}Zn��u[g���?G����&M�A(��sZ`�ľ b��f�h:'W��K���QRB."�_�!v��M�5 ��Ӑ-%̜�V�.t����8���c6���}���UkD|�ڢp"�װG��Y?�t���ap�l��9�/�.HIFp�C�R�b.��K\��	^�������oL� +�ȋ#���GW�}<�&ۺ�."�:�
��:Z��i7m��:�������4M:����ѐ��ː��suǪ���'R3���d�W��V�$m+�C�]p��e�Ş6��{�x��y���oy���m�oG���C?j1�₥��a�7�+^��`�湙7�j�� \y���L��[i��Gi.�+��D�"�a�������1RЊ����؟ ;��֏�T��7h����QA}ۍ	�b�5s�͎^8�����;~����ն��(���wp ��&�2jd���)>�n��*����킪U�hD��� Rj�tD�b�.Ym&�n��zQ��ÆUqb� ]Ok�r������iMuL=�Uʝ�����'� ����z��k�1"Ɇ��6,�;���&s��V�`VѲ�4�#��$-��k�T����@�QS_L�����7��#�<l��Ao�ȼ1i`����L�
�&z�e���ʉXQ��r%Ѳr�j�j�Pş��T�S[5���{_���͚�]A�]	*�%O�,
��R���/`�v����ַ�i0b�a|v�0����� �0�s/<�6S�.�ԬQȦ&�G��1�%W���( D��h�|��Jaa� �DG2
Θ�aeg4n׻���?������~Sü�� y�Ȼ3���
�҈K#�E�mE�o�����|93O�EFb�s������3�XP��6���[�*��	 a�I1-2�7��4���=�E�S_�V�`�JV��Ŀ�.�k�E�E��C�v�ZO���n?E��س0z��بW�`�[}�>��(��nMdLy�@��!m,���X��j5$�^8$z�P�\S>s�Dm����] ~#��Qd!pS=(~ I_�K�
#��'�D�t��61�P�v�!Z/n>����Sg�bA~�͝�]뚼I ��8����V�x\���R.��7���6N@�G���M���^j�"�5&��Pvz�t"��sZ�;a&�>��`5Q
x��UiTg���×�
�R�^-nC��v����Buۭ~_jҥ�T�4+���ZI�Ȱ��p�Z{����q��_���g9���xۻ@��2p���.�-����VD~3EĤP�%c3�CGWf�D4t�y�b������O�7^�Fx����_�����3s.�����D�������r�[��&�	�+	UA9��6����@7��x�q����[��	���E���o��s|��҇*!�Ik��|@�	�1E�(ۉ��X�3��<�^s�$08n��ZD�~lp��7 KD�b�����k֣H�j���������57+�h�w�Go��6I�41EH��x6��0��wXJ��)(�*�s��x�AW���{<�֜�ܠp�8u�`f �Dn7�Z���l��zPP�����	�"��ؾ��J�j|9&��H�:&G ���"%�V���9�>S�ޟ��ʸXQ���M�)(	�`�$	6ږ�<BC�R U�(�UB0�x����ŵbb]�"r��bE�R�?2Im�&ޟ>��Ò=;��F�_�Kt��  6t^.��1�Di�U�`ܧ+�f�����B,�P��j ��;��
���q�I��}��C��1!��n�:�$�M���1�M{������V9�D[���qs������G[Ri��
c���b�^���>:�k����ݼy�]=��2(ڸߟ�g����[�Q������1��8�26����� ܿ2�T��M�{���Qt[�Jr�q��tY�\�w�e{��0��;�!���ɗ��ϻg\�"���[+�_X�U?�̃��;4���N�^6�"PkX����n�
.�Z�����.�Z�=ӻ���F�W�P�N��>�7JS	0E9�@C�\q��Q�Gq��}�t<v�:e�y�?}��S��Ո>[ZY}	Ư�����۷����ܡG����'}��M���%�re�wT�e�X�$ ^���1�7�਺����8��H�(0v%�bPa���H�*{�IK�_6�T���2ٵ���)2�;������d%�;���D�I|�x�c0Γ�`�CĽD{�4'}�h͔Ж���)1)�J��'7Q��;%9��x������(e���*�g�ie]�Ԧ�vAgک�Ts�W�/'��C���&�=���Ũ
��)e�e�CS^z��*J/ƛ@�bU0\��\Td��TW� )Ch��ƛ@���L��d1�ν�h6�����;��2�	:$�8�f�%R=�vे��w_T�C�3�t|�&s�󭪣����L�'��7qǅ.����O�p0��@L�N�ܡY���)�;�鉮�M:)������Ԣ���!o���q��ΘHϊy��&���rL�;K��j��^�\E�aȍb�Oh���\��-��j�$s���Yv����2���~�W�q��27D�Ѝ��$�@ (�4�����%	�j��v�cs���Ħj�'YH�'o�sHC�u���U��ڠ�ɐ�C8���`����x����|f��ܙ*#E|H|0n)R( oT�J!(\5�z�!�CFW�38�ެ;{ˬ2��+~�;�_2UX-aE�6.�<2]��`��מ�~��Mq��"�L�J+��%+�nϠ���.�^�����cjN>U>��N�a:��kUY0�� �Z���/f���2D|I6��2����Ҟ#DPG_���� �����vg]���k@�"(�J�
V_���&y�L�l/Vx�̑�A/��=dm3q�5���I�#p��t���x�������3�U�Zh�?�ģ�q`�>���#����=���o�s �,_�q�QKc��jV�i���rQ�8$��������+��E�x� C0�6�T~J�rZ5��q��-���b�d0��>CIB�kY��%�E�a�Orl�����u8̑�zCU����'/��\��23d�����,� O��X�׍Ӫ4�$%K�<W�bY�arO�o�C?���3�my�3q���sF��#	'���#)�b�}�� M�$P�
1��G�����t�E�ȋ�^�V����\�:�ipq�vX��Ǔa���5r3^�Ba�b
m�0Y)��P�N�NCS��u �;�U�/81���;����b
�U�}����N���0i��a����#�	�L�I��ި-���.g�Ju������ Һb�? ���e�&;X&n���~[������?\q2 H'ԇ�3\�f��̹��#�{�9z��M?ٿ�7�$�[��lm�B��!W����b��?[�� ./�Y�x���/h�x�%zBO����(T ���So�ww�X��k����A˨:E�k�NY
�$7�)h2���R�R��}KZMu�����xP��P�4\�		!	��FRͤt/? y����%+?mm�?U��#}����6�O�$��B�>p��D��Ъ�kqw�U��Vh�'�`��~c@"�zI�Ml*��N3�X*q��x�6�Ɵ�{�xW�nN�[&@K��X���0~��kOBQ�[��=p"��ѻ}1O�̑*
۽�_���2n>�:	���d��,����f�v�����p6Ǉ�J5���Z��/�1@��#p�魎p�D^�ۜ��g�����Nx��;�/r�@!��˞5���:|E���;��mT����<a����{7|rrr7úQ7Ĺ��z��`�jSA����~y��Aְ$�(�1@S��"<�Ђ�s!�|��̺r������r�e:��ދ-X1�.WC,H�6* 0���F&YŻ3Y�Q����Q\i�"!�$Ԛ֟�'�!�Ód�|[Ȕ�X�3����Fn	IL�Ey��h�4�6��
�ц�-���II�m�Fk��ybic�{��eӚ��"�pr¤��`e�k۸G�>D���s�^�yq78Q�`��K-��"\�#�	�5`A�7[_Q-��B��C�m%W����Ȓ�y2�YM�ҩ��(f��+e֘Z6� e�aE��e����nw�w#2������~��n=��-
I�ue�+��W*�X�-*��@��!���EʈL(HQ�}�t��H,C
vw��#����/� �yI$�vl�.�8�H�އ۸+����׶�A�����f�Լt��G��qaj�/<���9��f���#{MyMD.�$GI[��DI
�r������ce_Y�ء���v�������f��)�:��~_o1ȃB?�!n�I!�D����$���&\U��4���(Ė��|[�Q�B�OYE+��AV��Ϸ�nj���ߟw�Y�Bo�k�,V$C.�#o��"��ح��E��u�	g�.�Ώ��zF_)��Ε�����B[�b�[|���[�E|�BUA����,��.Ri��6o�K�J~J2���\�
LZ���-[����RB$��Y�qWf>�v����4��!1��{u����3FK�@�@(��ODe�T�i(�}����}2`5�4�o���i��o2l;�Zr�(��-Q���tw��(5����b��O�\�4������C���7��'?a�π��gB�H�"��V�j�����	8��SP��2JYf�F���<hp'¨P|�r6����:�=�pO3��Q�,n�P�Ā����Jǜ,'&nVgY��WN$1'�&	&?5<A�#��<�x�D���o�J�
��@�,R'��q��߮VG^۫��2UX��M�+T��r�g�mw�l�--�e�����:P��	�*NuV(��3J�Dtk:I>�KI���SlA���v�4��_�0K�<�L�8Vn�dԂ�6�&p`��U�F�5��dOq���Ee��<���p��qҽ-k@:�E�|oӯa�3h7	�T�fN���݉����)BW�Q�Dy���1��ϕO0��Ӵg�Lћ.K�#L��	�P`@E�0���2��#�)��u#�je��WQ�,�a�?��	%�t:��5|Y�}L\&z�3L�c�T`37t4�݆��T%"��Nq�CF�f����=�ߣ��v	����[��l��t�m���B�>�4�B
�|[��kH�F�:|膩Ǌ4�
u�Dkå��U�Հ/���"�:�7o�-ǆ����l���;\|��S���M�:��B}�p�?�x�f����u ��j�
��SјUn��=)�:u��unP�\�,<�a`Nb��z/��h�d���Q���$c��:Cll<��EA�oez�Jq)VK�jha�F&vRx��'UC
�ː���f(KfT�	SZc���4�wz^f�A�LT˺5(#�6T��G��x9u��讣&p���-�R��7�~�eۑu��ib�{	���ͷ��oǙ|a�໪���U�J�����2oH�S��i��?�A{aM�0T�T@-�BBToF&�Q{���wrv3C2�r?g!B��s�!l"��7[���s���ͤ��G�T
%�źhX���/QO�0���,EA���.�UՊ�@*�����_��[�W�N��եs�r�/����O��zL�K?}���~:���:��?�q���/4fbm6oih�`�hdd��|�(JU%��G�9�h&Ϩ�,�Nb�t��QDk�� �;�BB��ܷ��kc�A<�TlJ���2T�<\u�TKqQ���>�d��&�\D�Lc^�Pw����D���Y��'��Q���Ap�Y6�i�����?.u9܊S��<���@4o=_x��?{���⭝b�WB��<v���M���8��_7���/'���������˘7�F+�o�RxT��10'�.�� <x`�P*�	�OUK#O��p���P���\iKE�>a�
��=� iqtƬ���|�Jא��Q!����@
e0,��p�aW�t[���S�ؤa�)b"j��4��
{�B;R�4���s~c6�����<�H{8�|���S�����ݒ�?7&��z�����F�"&�h�1�d���?��?�=j!��~���|/�w{cЯ���G�r�m���:�&��A��E�*������r�ub�F^wx��j�c���r+��cO�L���ȧ���^�<��HR���5��AS�E���~x��xr�L�ɨmbSX�Ѝ?�/N���$��cS�%�)�T�}稨����#�	�;	�N�m�@������t+݉����&�,��=�^*}}��RCq�V/�Q�f��߼�dN����V`PYd~p@�wc�%���_�v�6�9%��˹֖� D��bQ��)��n��|r�XL��0A�^��*[�E�<�S�&3]�M��}���}����X
��g�6)��ۧc_�hz�.�=ғƢ�V�&q��`�{�O��N��'����<�9��뇴�]:�?�$�o�~��)|kZg�HK]���Lku�i2�ON��:�B$f���?��wF�p�I���2#���dxF�yۃ�{��c��>ƌ)�SUP��n}}眓�_3u��]DF8��暬z�j�Y|�4���i�O�˔�F��_RB��=�3@6�H�w?
�O}��T`�U�l;ESQ9M������:L�С`�%�Z�m��Ɣ�Do,����4�I�i����Z���gz6oo]��vm儴�R�{�j[~Tɧg�آ'2'��������1*���ll+��"� �@Z(3Ȝ���I��g��
yoPp1���Js�)�~���1i�)��4���Lf7b��X���c��	��-�8���ꖹ��xG44�%�b+U)����H-�]���ru�	�\�PL~��J����#{d��"G�1��X���8"�y�|���|V��SV@J翦o����a𹹏�~�n8!��\!���x�:8D*��z�� �G/k�k|Nj��F81�4#�������i \X��~��G�bXc�[^8]C��-u3���8�S��ׇSЪA||��t1�&=�Ǽ����T	��U.�tQPJqj�O�)��Q<^uv.�0�����:]��jH��2����g��V�o��Cx������t#ԋ��˗<	L�Q�a�1����ŷ8j�XT �\d�3����Ph9H�6d���J���H�_}�S���r�3�T��U0��:YP��A�*E�Ւ!�A��&_��ɶ��ҵ��� ��&����(�/�nވ�����M��$͘EP��*FkCc��Dp�[M3��N��M�b5�aʐ͏H�G�1qh�*����֕�b�<��������3wўo�If�._���z��O��q�am�3��hV��E�o
Q������B��E�3�����!�����|��Q����ә���� H��
e��B�G�8�p([�D˭Q�(�]G��"QL|���F6 s�t��*�����x�.W�Yr,8���o+������גђ�BJ ����${18�����U,U��h*Sx�FU܁�Z��٢�9���	��6�pų��z�èG���ZQ���{����kc�?��s� Nl���RHǫ�1`��(�u���/��׋r�aՀv_���@�?��*��Cz�`	�T��$�d�YE1�:7��Ѵh�c��S�ޑb�O8�zf+�|"�(;Q��]k�bq��xF�ՠ����V������~�pKp4o��5����U�����^��-ZA�����&H���?P7z�
PT�U�|���g��-����ݒM��D��o7��V�& �p��1�C�;�RP��^���c�Y����,p��5���ݴ���`�o�&�<�|9+I(�x��-^]��]��w)�q���2?�F��*q<:#M�<]�a�����C8�g�F6T�M:�o �+F���«��C�G��t߫�"Q�RWW'KX-kj���9���K8��8�0��J/�T5�s_�q��í�Ͼ�{Pb�Q|��'�LL��c����!�I���ǚ��
 ǖ :��"���|���&j�S�3qWFq����w��&~�Q%<[H�%y� b�Z�b�Q��\㝌����-�r���>�������IP�����j��"�"J)Â[�v³
�O4K�Cx�:����	��?�3Gc��kf��Y�:������|sFc��� �r���=.��v�B�C8���!���*=�����H��|��'��^����97~\U��(���ű�^��5�B���I��l�����al-�WKA&'��񨪾7Dµyw�xΖ#�f�a�oY���N{-�9M�2
���� �}��=��]���qy����·}1�k_��A�{���E�S���D�S��0�G=�k����2gS��	l��U|EI�0���A�-H~Ykm�?L6��|�FYT�t�x���Y_�o��|�_&��ߩU��?/sܼ�P�Q�Xe
�<�E��9��^�)��q!��y���9g��f�F�_7��;B�>1�)Ј��٥��1��#�ZA��7�С�*���f�T��
�L��b�R$��x�9`�Ѧ�j�aڗ�}O�W��R������U��Z����ǯ:�Z�L�Za������ݪ��L̃q?k�,{�Ej6B�t͇`��!��ı7�%�HA�P4n��<U3��RSAK+�� �B՚���"�:�'�6��n�8<{g[S�8$���4���dV��������w���P"���N��FWt�<X�0TH���f:yE�'x�}�As��(����L���H�N�PB�sl��k���p��&;�A�(�̷�k>��� �����e\�Z�xQU���r�8*��V��oD��ח����t`�3T��Kx��T2�޼�G���[�\{*�紉{�#v��U���2'Fs��&��������g2R�_�;yU�.揳���_[���F��ˈ3�F;L͟=v��?��Gb�K�+�࿋�v�o�?t`�=��5���N� ��Ĉ��}�?3�l�|ƪ]����۠򿲚p&2�;L�<�����Y��[��i�A�
e�h
�T���ATW���BB�=��G�=��P����l�B�%���(�Q��L�rmI򻇄K����_Χ���7�����/i]�,��|��exJ���'00�c�)�M����4��.g�l8��/^�bP ����e"�������mYj8��XkcKTo��l&.�h���4I��!�Gލ��(f���l�a��@���O�s 7>}�*��!�F^�j�>��l��X��I i�p�J�P��^����3��Ȇ��&ݗ(�%{����o���U=�4���BTU~�Y�}.�� oQ+�mW����Ց��i�i�B�
c-�$�H��i�~i��	F�*L��SC����K0����9�ǋ�6��z5Z�4��`��$�#�P� Ҹ�.9����O������;�޽4v9�PQ����W�k~!��a(�@`�*
�E9��j_xAE�4�2~�"8������i�	����ef���!�>
W��J��gD���U��MO� �5���3Pu��"�5Wn-4rP��5v���0]�!�\$��{W߾LY�DG־�1F�,�o F�ż)�5E�1+��E�J�0��9p�r����'�����\Xo�e^w$d�?�fSD\tj�$.�n���`�l�a4�~*|.-�3)�9�g�ο���<�,�����a_:1�q�������v�ٗ�9v�Ma�7�!3+��LI3�$��K<v�3{�UK�?�Ђ|DjF�Q:�8z m�����kܿ`.�nɡ��<��$��*FE{d��%m�<=_�C`Q~9y����mȱ���P����^NJ�v���R;��2,px<NU�}����ش�`�"�lv%,�����z��3��-��[�J��6�mA���u�f��̿�F�t(%�uZB߿H�>�?�w��UʠωE�읾]Wz�����oi1�_m���e�kx�愰��0Z���-p�fl�d�c:B�с�C��1��Apϓ��\����OX��n�
с������ΐ�PJ\��B/���xC���z�-�zq�Ǝ��"d*P�j�Gq���>�-[�s�n���\|�B���P�Ri)}:d�H���{v�>'�_�P�N�a���EAN�#�_�mWݟI�==�e��e���O׾vⳄ����%��[:}��ǚl2�*5�{�O�w�+�U������K�n��h�&_T��	�訶O#���z|p���:�����(��Ӎ���\��p��I�٣�����W"%��3]���1j�PqZG�L��aF���ݞJ7��zO3ߠ�F��2�6!a�:�������>�Z���"����Zm��'���s}���0�%I"�����A�J��j�a��Dۮ-"!2KR:�^�X8X�;�LtYt4^����d�4��c�^�rs0J�����F�C�H��[����{���E��E]cK���kKf��
	�5GwM���SùiWx��W7��J�j���+x��w������Rd�R�$���^]���=t��)�!U M,G���R����j\/�(s{��"���l0�:��_��簆��0��1ީ�����������<�g��/�=q���o���QZ�UB�E���{�1���O�媃?d��V�̂XX�]����ɨ��� �P��:e;c`��Z=�K[�.�f�D
U_{����rcR���NŽuM6�>r�K���'�Ҿ��R����I��e���B����Rb�"ϻ(��?�;) ��=X�#O#�cf1q
]8n�C6!��������Z@��|a�7bJw�Aѽ�r���y���W�aco(�	D������ ��n)4daW�#�iws�ZW�l�Wd&��9�LCx`-�
�J�Y5;=Y60s�Gd���@�~2L4@<�3Hu ��0��Y[(�x��Wհ���O�S�`���;�4/9ڜc��ؑ̉�m�{��n6�9� ur�FLwJ��h��-��ϙ�=gI����
����TlѾ�T�a�;Ѕ��j1UrԝB�c厵{.ԭ���g�3KFkb��7�Riol�׏x���J�g�T?��"�ݠ|�3)��:����pV#�TC�d�%��ԨJ'���V�mb��M(�2|����ަ���*;/���[�� 3ʰ���8ޘ1��&)�1V'8���JC��n6��j6W� )�;��]��	�o��G���� ��[��cm��VP|�V1�(�ߐ���|��R�{�/]Z�
Fo��4;�����i�p�[��^�uLW� ��V]`m��)�Р�7���8����
�^�AzJ �g�Dp��);��gY<�lUr����}ɍ��L�k������u�?��K���Y�Ԏ$t�FS�S
�.$���_33��h���k~��v��!��.���;"�vX�~���߰� l]����}n'�ệ���+���/VV5�ɢy�� +n�zr�~g�0Xb�nB�GZQ#��,v���v�����̭`��8i\�R�
U7O�R:���-�x@��j⎄g>�(��1';/n(J��/K�F�}�H,��L��Ka�Ld<hQ6���+̫��^�B#�[�_����B.�R�(��ުʲY$B�@��D����{4��hњ���3�,I7�!ȌW�sNrH�/�0k��u��V4�����Q���A��;
�w-�S��H�ė)��I�!?\����B�?_��,$/�ғp�JC�-�`N��H��"6��`]T��m��iUZ/��0�<U�e\�{H���Z|ff~�,�!y�������V��[ў,(ǔĂ��-��nF��?��K=Ǧ'._���Kb���!Z�H�P"�L�w��������ud<#�owIQ/|TЄ^�,�6\�H��*��L��Nq?����>�j,k�3vzbS ���T	l���
;,�&'a�DgQ�|j%��鬸�ExS[Ɏ�ll4z����t ���88���]_�\����-���>�4^�Ƴ�[�4	,J#>��|B�JC��ֶ��Z>��ց�s��\�����6�Mr��Tld��$]YnJ�}G��k���SJ��p��Cu�Cb���
�=ݘ�@����m&+� X�,�,%�Z�?J�m�GX�M�VcFErj���C�tJ؎�����B!��h��Z�iD~��g:�GD�@*���@w�IXU�ͧ�˶�jڦE`6SC�H�H�p����C�G)���/�٨z����ޕ�4_;���Sw����lA��:���~����L�uZ�̽S�����X��֚j �;������)�Ȟ�	�7\�c�v�v�V�L���Apj�%#qΉ��\x��>]�u�Q��g�͵`Dq�GW,،f�F��������/�A���<�����j�K�jxͰw�[�	�u��8Km�����������/��r+�8�:����?�)��)"C��0U��U4�*N{w
+�AQ,���n�xj5��<%<%|~�)�Kw5��i�:��@�#

�4���;�+�� \�@eF*8�h�� T �eJ��讷�����X�-�X�����O�6πK�Lp�~h���y�z�?�/���Mô!
�9
��0�%���T���"ߌ�$0ǈ��sm�8j�;|��!*L��F���m�┙�.3T�g��,���}Qٹ��b5��~�����W����`DH�5���ψ������V���}�?,#�"�oֶ�R�G��$-:'q9�$�?��v�B���%�9˭�lwإI�K�g�5Ҵ�6>�sN��eǲ�=�8e�u�8+Tgdjx_�32��c��cb�%���kN�Sy$D�Ѫ��?�l鵺�nH%�'�o0'dBw�`ʕÜ!7�k�G����cJ�����lN��P�O����x���*�~zE�����	�����&��޴��������Hn8_c�ʺ���{zr� )�������x5�	�����S=�ɬڭ�RK�wӇ{���a�h�Oh���4�����"CD��t�|l73��MGլ�&�6g�	�)Z�|��_�PudQě�S3�YG m�+���%���-�>���)~ ���s]D������oS��vV/�=�Ce�0qd?���L�5�Z�v:���� ���[x���)V��B���/���i�I��s�\�P���J#!������6�_:�;��w�B�-�ܬ8�ܸZ.֦�b 
*l.������~}���ye=/�Z0�|{��`s~���jη�G�d苼�����}ۿ\�W����2�2ҕ3�&��3qP��q�-猹�2ȇ�Vt~Ea�="�mp��^�`	�@X<Ǵb���� ��Ozz�=u������e��.����T�
�Vw�]R�)8p���7�n�q�\E��Lk�N�&�f��܅�?��δK�*a�b��b\v5�4��h�C�n�x�!4c�4���z�EO��Eb�
v�R��_�T�T��#Ѽ
r�~�R���x�K�?�G^�&�*5�M�����S}��,g>c[�̻�r)H+U ,8nY���87�,T�c�xKLz���9yX�h�B'��(�����t�,��v^'��ڽ�|��C�����[�bh��$�bwVi���۶u��l���}�q�e?W��K���ukL:VS3LW�Z~T��
Q�29�@-�:<1i���_&\NIX+�[��v̒��Ŏ }����Me�#���3�p��\��jNS�;���M3�}���!\;j��a6���3���-w=y�o�O��;ΤF_�����_2|�I�[��&W�������׺�� ��ak|S�(�ҡ�5L(�!;L�X8�MBV@e7о�)�(�����m��l������n
b<���=&Y ��`��]P[�^.�(�m4���"��4aZB�����)��{�j@i��n�r�J��oN�-5s@�XF�b*�~l�G���\GbCY
�*���}
��S��Kj�9�bAJr�P*u926��_��Փ�sD��:OV�C�㢰����5��ʎ&W��t���/�y=g�;����eȢ��Z���9�~>�9|�%���~���O��?��� ���6�5wF�ߗ��Kؤ�#�=�:<6���"0I�Q ���pJ���śiܠ	�o#��NF8�>?O)sɦ4Zrٰ�8Ş����4��3:�&��!l_IA�ќ!=`�O�鯓�)���qC���f4��c�98�ޖ�R���l�[G�ނ�*8S��iL*���$���Z��G"���¸���a�}��~U������'�ϫЧi�{
�a��#�W�5���]��N�XEkN7:�Xek2���O�.��8�<	đ�qAS`sv�ð����.m���l�f�q�!Jv!~�$kݾ�f�%;*��!uU�����7�%FV@n������/¼�9&�,n��v�!LuqIָ���bW���u�ʁ���Fѹ�[���0^u�o%{��7;�PD+�/�,)ϲEծ/��4�S`e]�4���;�ضmk��ضձm�c۶m�I���~���Wk��QUc̕h{�kE��p��m>�����a��1'7+�������}w@�8Y��F���}E��ΆR.V�t#����h�>�$
����,��-��r�K}$6��|&'y��˞�.�Ɵ��I\l�v$.b�K����`S0�����򕤡I�<�J�%J,R �\�3�ʨ.a�GQ��q�b`���R�t�~R
�>����}=D���\�=�2Og� H�;O��w�f�$�H���X��:٬�bqD��wǺ��brb׫(ie�ߜ���BI�Us
"#�s5 L�߭+�2��m�H����3�ﻇR��M"�*�gL�����g�d���?4��T:�٠2aH�@]�Ot�ﰞ����Z����x���T��"��fJ� ��a����b���5;H����$B&9UuX�߭��:m�P4Z�u����:���Q�<�l���Бmyȇ�f���|`t����ث���:6	օ�AD��~C�šP�a�`��N"+�d_�����Q���FҨG.����A�80"�2��'LriE������㹯bqk�--M�3Ú0[�`X�:�{��ΧZ\|�~ݏ�O���p;}Btuzd����:�6��4�Fk˙����	d=���\b�X���hȓ�rX�.����&so��ݴ�'L(C���.�uF����¦ `��9&3���dg���KNf��j�u��T_?𹄷���+�w�֛R�W�B=��)��G&PЯ��7�%��0��4���2su���0���f�x�_.׌ٗ���Y���33���V��F_����_����?��W�����EDW7_ش�5Z�ٯU����G[5:Gr���?�4�}�f���B��������mN��L�Z���7N4��������Rrb�Ŕ�c[r�9��6�uT�kq9��az_e�X��g�>��j��<�t��M@��I �e��]>Sn�C2��[.,����(�W^��dv�҉����[�w�AZ��,����k�z��%�&������gTL�>�8,����4����̦��E�H;� �{Ɏ�=�\�r#��� �8�� b�����3�]�7d�,m7�0�>�>��z��D��P��aU������1�S��7 �����]`�w2J?O__w�OJS�W�N��T�Wbb!%2�zf�x�z�q�����|�b�D.�J~AG\��(�al���l�����t��:<��g��tR���a�R
���g(��f4�Ң�����`X|D�R8Q�%���'��g��E�4�Y��/�5?�%��uk�cZT(!��໭�U�$O���~C!��
�_L9yĹ㚜``��$?S"Uq��i�j�(6��lX�<�\X:�GқCB���o��kT�X���d��;{[6��}a ��Ԭ�V�s���;��B+g����AhZup#1�UX�T%��(�0\f^�00��h_Q�?��̨8m�W�*1�kJIv�}|���r1����ޗ>���n���8�W��d�����.@����9u��E5�yʃx8�M���%2����o��4^����|n��7�Ԕ�!�|^4"!���8m�Y��_�Pn���k����B��.=�L�����bΨ
���0"�E%���)wY �sJn`��{N��g���!G]���Ңi�\tkۍ�o�*3/4�����'+�0�]W�M����HjTu�J�tq�z��AQS��bp�!�gw���
������L���2׳u) ���N�@iJv�k����,�$���=Q'���_}�_YK7m}ڸ��:��K��]�1�� ������A�R>�ܢ_1>���6�XP��i��/AE���>$nA�����y� � ��"���v%N�Ω�����?���';y?������H�>$��Ώ�|¡�\�An@��4Ԥ�ӑ��$U��7��^l=�-:��e��y���(;O�!�m�S:2��3(�(�豩򫍖����:-)Dƽ�,����{��.!�T=�_���[w�%�c?�9�%��fZ(��CS�}�X��\���A1T�~���B"B��a�@���]<�(��7�TV��Z�N_VV�N'	�(;���OxN/1;��0�SmPhZO�%�����O��0օ!q��9w;&:��
z; �dx
3f5�x��k'įdۣf>;JNBZ�0gôGn��a���1e7��9�(�������Q�޴��|zdd�xV�uN�����A@�C�1�;!���3�� �3cVa�oᆚolW����r�[7*�R��(`�\�TS�T�)�BR�q�����)��K�(9�T��Ti���5̎��(f���n���y���� ��n�cm1;}=��3��Z��XY�t.ۀP+"ǟ�E�Y��}rr�NIT�V>լu��c��a+`�WI*�D��a��])'�s�o9�:�#B%�S�
���ւyL�ֽ�Ki2-�M���2$�	��t~^����E��T��iX��G�V���ךF�1�R6���nz�����䙆�Z���$�[�����~ �_,WC����sl�� X���� تG�5�O`/uw�ҽ^W�̝FG�����m�z�!!	�O5�_�bA�5$Q]Y4&XU�x�-�TY��F0���TUU���E�eZL}��4~~a7�¾���A����h؉=iTC�¹d�\��@�$��H-|�R: S�C��4J�jة�x{�]��f�L�~K��������'ԡ>�ӖRt������KA56;����@\Zn�(s��>�(s��GXXXvN���r���&���Lρy�M������C�D~��#D���z��G�Z٠z���n>�� Z�WQ��Tr�����[�{eB�e-'P���۟�0�dhǇN�&^��0`�?������������G�1`@T-�h3_�z���
��m+6�H&g�{�}1v��?�@d����3�f�Kr����$@РN6{:�'��@=���<@�,�m]��d�?Q\�p>/M�&DX�U���p>@=��R�ە��R�7!7�xs�C�>N����ꦴ:����5j{�*�h�|l����DX�	)4h]%aP��Q��b�z�A�8�u���L�6�}yec>c8��޴���������Ԧ}�4S)���p\�7�5��mȱ7�&�e��?�d���M�}���Y}ő/K���~�����a/�٧'Ѓ{/4��G�e�8��K�����!�ktߙz>�P^���Vmj��]ȖP��%*����Ņ���P-`�6��7��>9���߽l�gj�M_ejB�%I��s�VT2-|L�iiӷ:�g�����@�8��V�uƕ�.׺�K���>_���;k����N�#Ɲ��K��f��H�Q��V|�(�ND�A�O����\|�̈́�!�OѨ:��f�"g���䠚t$2�-�@�@K�:��'�ħ7a��B����‎DSgq���CC��}��;����1]M����* ��A��%��膦=���U<�u.�`d�.:��o� y�{�c�q��ћj����/n�y{���k�X�uW�g�BKӟ{�e�g��^<��s����z}�Ē3�_o�~�^�AMq:�Z�\�� =-��7�M��H�גf��y���sr|��Gb�%�t(r6�.���TT)"�&p�����l��ö��z�B��JD��g�j�iB��em�1�l�W��jG���ȒQ��w��#g{���4%ItA��$@���@&2�}*e��X���azO�֪+��7��)����P`z�B1��;���'��-��O�/�Z����*�#����]�(ui�^C0�3Ji@����Ƅ�fM/vvX]$=,_r"��q�{��B[
e� $���C<W����`q�>��%~�̑��lp,t���wy�k��SfY�5t�ϸ<�C?�����}��2".�^Y��h�ꕊ$�;�cJ��8����y��`�Z���� �!�v'V-�|([��|�͟�r�ev��c��a���3sxv�b��24�T_s�7���۔�|[���5�w����|�Tfveg�[��Tf�m@����OTA�E�*��Z:������]�̂�i�n�_����� '��R���ف��R��y8��7Q\C錌�E1�t+G���U�w�$������b8�����Uڪ����Kf�omKo���4��]pn���C���ɾ��3X&\���
N0y�-�����|W�JR�����z�x�|s:���)��z��b��8.]��F>��v՜�KܝbQ#���ʆ�>C�B�p���������4�g���&iXZ�#��D���m���P��mheQٜOM�9BN�9a�E��h	p7��ϭUH��<�}����#�+o�/u�]Q�&�r�Kf[x3�H��l#�yɏJ{�A��f%%���3���������$4���M���r�Ҟ������1��,̎�?1nF=��G�2�6h���޵�N1�+�9劾w�e�ۥǮ�Ru�5�N��!޵��� m�͵��d~C/��oNT�Zt��'��~��[�֟hO`=�-vD�@�7Q,�@7vC�"7�$JD	�X[(!�p:���"4)���6Q eă;��<+���ϐ�t�=�'O9U�VG���F��`�@�i_y�6�W"z7��G���a�PqA���?gDE`nS�/�gx��H>�0Ms��tWΏ��x���ĉ4{�x����W��P]�4�C~��W#�����~��Y�p�>��X�d1N�)s���\�?]Z����;J/g�22�4�����5ޜ&��Ym�,�1�ƥ�8�	!����:�'������z��.E%F
���jSd1	 �Dx$��v;�&���r=/!a[**c���h�e���q��vԩm:�/������i��p�+��3�஛Y�Li�������$s`��Y]�#�qf��
�s|E'a�����WH4��R揙S�3�����	��5���$�<��5��� �k%Z�4Fb��! P��ej����b�K۫os:���Ȁph���R�c1�^� zM�n�&��Ā�GN&��ܽ������"g��C�RO��4�s3[o<���B�ӭ*��JiL^�`KX��M��t@NRH���l�AMYPI��;VR��=�7c��B�F3�NP����V�׀4�-A��-|�6j��X���V�g�����j�>pa�L>��E������I�]_��.Ϙތ-�	- ߦT_Q<���>
������I[G��� ��$W��2>C�q>���D��"`y,�_�oI%-�AJ��;<���:�-9`D7r��~;�������� j$N�0�O&^[���կ���Ҟ�Y� ����^�[�a|��_eN���A���	*�����.#�M�cP3��u��o�F�pd�4io�o����T�o>��k��E���I�� �^wx��e�G�����:�ik���B�ch�C� �o"?K|`�mS8�fK���v���-��U��e��X�1�9�_�f,�7�� |[q����k&l@�D%(��Z�GQ�����^C���;��9�g;7i���0TۥI��I@�Jp��*.H��d�X�5"���p%\ |�IPҐ��6�SL}wy3ӈhoh����6jG�{�������֛�[�-���s4=�v�=�M���;���S�ޏ(��G�< �������|韛f�&��].x!�6�����B��5v��@�y�T{:;������	�Ƌ�yme��D%��k.�&�V�D)�8g�q$g��ʦ�8m &�eg��QWK 9��S���
R�v�[��Cf�}�L32��D������Eb�#H��CZ�Hj�:	N�z�sx��3��x���J��ʊ������g>ZO%k�S�',G&����;��C"X̥
�z�e��U"E�nc���Z�懤�E5daڋ	EC�."D�#qi�ŷ-۸A�;���
�`h��?7�y:Ƭ�E1�[� 2�80_"����@.�w
q��Z!�0��2��<�7'��i-���;G�J]C#�����9��˷�e=�sT\����U����H� u�2��y����8$l��M�&����kBs8�a5�E��?e9����K0����{cI�g(��g��a���%���5PhP��3�����CW��
��L��@���2A�P'����N;����E|���J�c����i0L�w�_b�%�j[8��.�R�0�CN8�t��˃�f1�*��E�њ�u t,ZWǲ�a2QQ��+=B6��4S�|~���f�f�S�{Z�Ӳ8���ڵL�̮ẽ�* \��-.:�v�_^���Q�����Վ�m�鼵�O�HL��տ#����5m��#V��9EA�^������j9]���aM�>2��i�/D�*>鹇f��J =�������/J\�&oÅluAϥ,˂�kq�pt�I5�n�.�B�}�
���S���=��E�H�擃 ����a�|�)
�/Ea�Mq�=��������ZX���w7*JF%�D| �q0�,/_>>6q7�uR��K������f����&LHv{s�#%:�!�ʏ�u�)����R*�*,�h9XN������N�!��1*0��Sm���x�	�~�����:S���	�T��V�H��p??Rk>(��$J���=I��+q"�̓��y��TG䣏�� ��mWq�O��}�9��ef\��GN<S��A���&)$5�Բ�����c���F��oo-<�s�b������v}���x}�f�뾆��?54��-^�۱N�,}���6�u}��߰z��yHKrcF�i�EnRF�@�9P�.fr� ��(u��!�-�O��pB��&6��]�m�P��LR���� ���OC��ʟ``��_ϴaB{�RjBgx�U�-p����HΞ���'QT�󁵄��@�E��o8d�=�3�q�|}.}���AV|�Y��A���+D��g�"f
�,O	6��Z�o4\aⱄ�]��U�]�3�>�/�϶EC[(W������u(̷��{=\#�d�:U��>)���dŠ�
��L	~�D����#ؓ!(����V:ES��$��ǣZo%՜��ӧ��I��	��N�J�����?����M�]-,3�5D���x��Ԯ�h۩��ړek�\M�y�.�]v�h���r����Ue<��d�a�)$-q0�)U���Sʨ�4����W�B�,�y��U�E��tp��s�w<�I��|e�yVL��Ӓ2�0#02h��Ou-�BM�t�i� �X������(�,K��#���k�iR2'{Lꔨ52�W�J�����R�g4�Z��8`�G�(?�VI�<�r�hK܎��x��T=���}��W6?	P
c�4�»d�Ү޳�'|�nJn��*��=��)	����_���\���&��n�zl�:s����&�0�V��k��J�>1��p!X���C����,�f�Tk�7l����׿-�_jl���[�������lP/��D�(��\��a���2�j�w�d[cYoՔ@��0-;ۉ����>�ݼ�4�K�d�R��;�`�2�� VER�K�7H9HH�a�Lr�W��;CJ0Q���7Ń[җ����s��*�pr�B�������7���ֺN�s��u��T���d-��=b�r}���@�T���8^��=���?F��6Xm�6R�#̢j�,����L%#�8�x��>GK��>���˧���v;RѶ�V�*.�Mx�]�f ��FS4~'ѡ�Z�6(�2ӣ���֟H��bK��[zȺ+����	N�<��*�cwB�V�:޿�,,�_�Jm��&[z����Jջ���β��È��I�Z�u�6M�����׳ٗ2٨�Į"���;�G��x���1����u˃x�G��0�w��9�{< :�����V�a�_��/��)s�uzTF���*"BB�{�k�܁*�Q�i����mkZ~߾\a���p�PS�B:-�*�+'�G��KĂ��  �	��W�0\����eǝ���H-H��ᩪ��=��R�q�f��7 ��kzh\�j����Z.	h��?,��S3�+��Qe�ׅ[�9(�xA�U�X,=m��9���XQAˎʻ�TV�{�rĔ�u�+��������Ź�P��}��/b(���I2��[;�q���
�:�5�} |��\:==.��?n��0h�p�����_���yKŴ�����[>��^�}������\y��U�8�~�����46c�1�:��K�N�xaDBelq,G�R*�lCfC'�g-"�ъ��Қ�v�~d���qhS���.���p��;&�! �( a��d?�!?񐦄RlE��j=-8F^ج;�£��3��<Z�<�4k>�.�	m�J�~'$@]y�e!�l�5,غ?�n�j��X���u.l�����LF���T�H�-��������9�� ���5�\&e�n��Ldת0�~J��Kq���2�4YT�� a�T��8�I!V������5�K�&��9�T5�RW��_��X�R�l�w���:�4�'bd��m�{t3�<��x�����U����ph�?W�X#�l	6���T�(y�C��\g+������G��B�U4�Y 8YW 4@`>e�h�9�ѣ�ܡt>_�	����Ȗ���4�Q��yӈ\��_��<|������ۻ��Vo��x������C�8()�O%uU��5SQ)H��K�OL���"d�^^��ʒ�I_�8��-ia�������+��.�CWn7��Mܶ[���~]eɠ&�
UK����
5\5WZm~�v֎"�?��p�B�8(&g�:����ǥ�������)��}�lc�"#�r�F}�ч0*��Һ�&��g�/nТs���+����^[࠿8��ZYd2�[�J�Gs��Ǜ/
*���G���^{��f&2��,�N��������?��W���Kv��:Q@����N��� �����5x22��BCCod8�2]:�e
"���gK0(qX�ս*�9�?�0��oC�A�`@bo������&;���|��ZQj��u�[Yo@&�*���|1�-s�s�5D�'�0x!hL��#�\2�$���Aà���o2 E&Z�	Q#���@�1�4�n��4�Sg��z�C~S�Gm5#+�
dҕ�{W��aJs� 7��G�D���{>��wSo���|��	�?�-��Tq	�+�$��� ,	&�y
� ��@iXhU���=V�����u� ΅{�P�6M�R���j��x��`��|�=ҙ�
s3�6�H>���t[�!����H	�%e�l#���ćs8� ����4�G+f�	�i6f$�D�q6]��\&v���o�y���,}}��j���T�ܠ��k���9�7QM͝wy��3	���;�񷌖���{�(�ca�崘�~����������L��m�d��2'WfX��Ʃ2�_�M��qy�E<N�6���h�b���):��cWq��%�%07��C���Q��@ddt���a�O)�^M%{#t(]�T%~�#rcDA�l��ࠟ�;�!�M�'/���NU"��#��T5� 5��l�CTY��i}��d��{�  S���(gt�u#`+����vQ�%\�k�h+Bqɰ�j9>�z���Ş������[�ޯ�3�7�_��Yr���G�ϱ���/66P�7,q*��w>�#�o�l)����t��'������B������j:����Y��`N���NC�v�r2���������l�H���)��c��w��uiA��'v��0�V����AO��B�u~.*�e�[����Rky�(�#�m. H�H�{B��C�!�*���Н(��q���_Q�G�.��ReAz���R���R�$S\ƯF����]kL�\�?�R'�'&jZ2�M3JX��x$�?*f)W�]���t��>a��]r�v~Ѯ�w�r4������A�8tP�4���>FhkW�����Pϝ=��6V	*c����X��UAK�ͺT�b��چC���b$$xK.�"D�'��e>�c�S��t��;EV2���4��i�o���?��:Q�O~�rΆ]5��V�֮z��-�dZOc�c`�hL ����P�G|�`=�h[����by{�*�6��|��8�7z�l�)���c� b��|~���THC}���y��B�]^����6�v�2t�dgn���[0�)��E�M�Lvܪo��q����X1@2���a����V�D8�
�m��U�@9A��j��\��7]i��ȅ�ēd0%Ñ1�H�։��{��qa�U�)������`I�������VNbC�Ń�HV����B(f䖾.X�I�| �񸬭6~�$�R�*dDќ�;�
$�w�A9&-�5yԏ�x��k�ĥ�L�j�P���9��S��^'��:�4L���4��Ǟ�~����t���|���j*M����������n<�ٌ�b���m�D'�p5nI���|v
A�s�?����	9�x� ��0��}U�=�( ���Y�$� �������%����}�ࠄ����W\�C�y���I'�|�܄�!b�gø���ejY��~E���oB`�����@Ŭpi����ʸb�ƿ�����kNTB�F��J҉�2��I*i���@�C�#١�Qa�w��R�.y�9�9�����Y��:��ik�E��I(\�l,�7�i�k���e��{�ݛ��f͓t�Os;!�W�� $q�B`̃�{ܲtEĠ[c���4�8�?i'���.3�zL}]>��Ŝ�XD��$� ��[�h��)�o�9�1n��>�Fr#-`n�7?܈�����1��3?P(�|}���=���"7]n�c�rk�z�Gxxy1�X��^�{��J��^�L�=�y���mN���X�����oc�ū�"a�&R�@�����解�kO1�H����O�J{^��^�v��F�h���f�&��V�I�A��(17ʷ���4t@M?ea��(�A.��Pf3WT��俜�e\"�܁4�-Yܡ�wn�T���Z�+�zvB��24o�����lbX���V�'�9�~D�xT��q�yb��t�}�keY�����0Qs�&!�41v;��N��pk�ݪ��p�m���}=��V�q�ӊ����v��x�������n���_�������N	*��]hzjj��FX�Y=o3�ӒD55la^���5�&]4"#䖣���}�!��&�fl ���B��>oOD��;��ic��=;SBұoP����K�<�Ȁ��e��"<���]|���QB�TڕF���3��	p:xm˝h�����'��/�~:Y�/zR$��ٺJBसe"�aP�]�Gۛ�U`T)cMt#�{����}�@�xyh�qY�WrXC�"�U�	c�N��zɨ3��BP���aZHS7���;*���	�R�A09{+�h��J��`���|��O�DZ.�����Z�. �=g��8�������9Y�l�w�����=�/_� #7�}a�P)N���NVe��p=pn0K�3��󉼏���>���$�@3�&�y$����==_�dU���N���t�H��ARC�Xq�B�+,��k UR��������q3��trv7B���y%�
6��<��Y,���;;��]a�B��>�����p�A�'�ܝ���(C���C��piE0�_��z���
�R�>6��-H@4�>�8��WΘ�R��IvϨ��QY��<L����H]n�I/7Qjq�s�����#eʟ��c��{��eB"�����2�1=�ȤV���0�b�F9�6d.ē娣�@!�7BC����^:Og����ɮ���߮�����¡3���8x:^�l��ݯ֛ngD>�O�CC2l�q�B\�3��O��#��M	m�ꏿ�TB�����,a��׬!�t���.Kf����_NiG��yͫ���3*01䊃�Ր}ঢ়�,D�$���4�r�8�|\K���8F�l�,!^
"j�����9v�cS��S*N�RH�)H�ا�E�m��������|�'%s�?�_.�)'i|����\;מ�Y���p��YM���K���" ��OQbv��@�W������P��ݦ�ɼ&1�^ Kxjevi�w��8��k��+��<<���
��fҰr�/Vj毊�T�����mW@�3l�.��A��Ѐ��Ƚ�Հd���@����V�`��e�ci���a�ё�4�d�t�w�|�7?z	��0��-��u�E��U��{��af~�4�(0�F�@���|�J	���n���u�F��)�ԦW)]�۷�$G�������]R�E��O<��T�ɟ�]2����M���(��}�g�1��Ϸ[K`.���8�*��?��V���~��d�V��yՒ ���c�W9w&�n++0qa�Tl���\��ȕXr�tH�D�m���F�ҭ�VQ~L{��R���PkB?��'�]��}�pMp�Vq��w-p��$���i␽�U�����N&�9���8��n��	;��C��渑<�����7�i^2j[���<�\��3j�Ɠm|�F
�JN��]���59oՅ�����-�H��	�{"�xy�L;���W�d����LB��=�sx��0<�����fkiNA{��C��@�g^7ؽ_�	�������#Ʌ���B���Zv�.�	=i�v��Ay���	�_�T��W0s����ÞH���
�u����7d(-c�<���iߓ��+��t<�]�'q�㛪�>'s�Z-4�w�=+l�Ug��=�OA�ʫ�0��i�"e��3���6�]��h��g��mZ����AA,�Fo�8�v�T�ᕬ��F鰲s�?�WN/��g|�O����:\���l�+�����ޔǊ����W����"��EIWv�2F��i�����↽^*���Ÿ�>zڜU��"�wGA�ϯݫ��Kv��b�ƅǧs����
���*�Zx�������h�m�P.��<2ߤ�/�������
�
��A�33(���\�S;�)LW@����� :��Cpyԍ# �	>H�꺅���($&{w�N���W�3WI�`?��\#a�Y���A`_q��5�L��.Rx%"��Rt)����g�G�;�o�T�C `U�Rs�9a���Ssa�g��5��A+��Q�
?W�q���H��m���dO�2�E�
��_����D�Χ� ͝�#;��[����������ַ�I�˹��Z"��uvVZ��V��1*�H����jV�｡��nì��4Y�!8�4m�}'����Ǭ�%�C�"H+��FV��^�h�N�{�(�?|D�SV�� e2��:Mt� �hO�9�����S'�{������Jf�ۯ��<B�����I�q���{�:�����`š��PM�r��&��Y>)��~��
����i�3Ss��;�bt�l�'��bm��=�	=����~�.M)���r������xt��)Wj���9�Ojd�y�!����QSE �ͪUimkt�kJ<W��:�q����^��Y����$zE�����"+"��I#�EsY�dM�Y�����c�,5��N��^�������b����Me����%��9x��ٟ�JTUdd��$Y���C+��Nz���zL�Ï2��.88����s0�&Y�=��ڻ����*!M����gƾs0�e��a �'D�ޕ��m�Ps轅1_�ǂ$Ct6�x	����@���
���uJԽ��A}�%���(v@_��<u�#i��ܱ�<�l#�T�'F�g�و��J��zB@}X6[D������!���
�s�t�q�I�m=o�ؿ�S��ا����Ya��5�������x��yxx(3M3������?��<�6I晳��|̑���:?���?��ǁ�C�n7�UU��ˮzwǽϒ����I��"�G}��韧-��a�\��翩����6i)NN�Z/.f����PW(�Kk�gE�pEy0���X��L���{j���
!�B�V4F�umc/��X*
~��C�@`�vփ0R��i֐�G���幒�.1C2m!��%:z �!W��T�X)Tkt	�g^� �h�f[I��- &�L�#��;���=�cl�m7������\!J
��I��
8h�G.`�.7`�D�*n�\	o?T����A={�y�|�d�����XVv���(!���wyK���$N����rbNfVI�l���E��v"%J����E��~��Q����Rir�%(�ǘ�
~�MU5�m��0��b��^��O븪0��Lp`~��B���#�,=#�-y�cڜ^j�!���,-�^�u�X�օ;�nPQ���މ��9*Z?~��a��"������+$��
�ȫ�N���O#e]����k�sK$V�(K�!��a���A5+S� /�v��ȩ��t�ˠ�I��o�KK�&��3H���)�y�f�H�~_��ںoNU�%e�ذ#��C�ow��/�nV8�햝R[�/���I<�g�ֿ�ߒgpMU��BU�]#Ku�k�9@�Y������Jh$��V����ל���7����o�$�Z��X_k���h�6��z?X?����5����n:��<{���]f����*��]���LX� �^�6{9F��0❲8�'��i�Ӽ(q�,ug9j�� �U�8��q���7����rb�.#Ĵ|(�� ��'��!pQgݾMAV��Ne�:Rו��j.��3x=��$\�$xU�e�^�Ƞ|e�]��Mz:fXk�j��6���W�_�m6�<�q34��l�a��������H�#g~�'�g�g��N開�S�1�׹����p+�8�
=��>ק>5��a�z%���c����Ÿ4l@��ԭd<w3yn� ��˩5���A���s��U��B�׍|���eǈ|�[,�	��4K5�����Jo�)-�uYī�L�6e���(�u���5����~��VG��D�F�;�V�Gb��Z|��F��\�K�`��^5������ �R�*Z�忯m���*g�ڷN q�?���2�����`�Ue񒌀����5JCVq�/r��'�	�aɭ�Xi���W�O2�#ԓ-������3rQ��T���O�����{��D

md�"�d�����BM����dǜ�w�$ʟ3lߴ(���dp,i*%��x醃>7�HT������6��݋#��*��f=�;�����=���z�G�gUV�i����+��q'U���|O��~�'��5M�_M�9DW~�{��4��������x{c�n�}��"&�]�J��ϗ�>��]FA�-��A�%�](�����˘P��?'�ύv�����.��w�y�(k�����*���x�\+�� �����
Bqoq5j�2u�rJU{.=����rU�>���V;A��*(�D}���H�21��y#� )#~	�Q�{�� A9*5�,�=P��5H�ߍ�$q$���j�{���[㨛:�6j'#0A]��Ze���}�oJ��C|a��>��a��x���B����I�q���4�C�t��[C������H��͉��S?2���|�lqT���¤/��GO;rZex�]�,v��`����f|���F=Oc��{��}��>1>�}��ގ���ͭRLxx��-��[7�qD��������v�V�['⾤u�ݼ�B�F�G�'��U^�"�Ӡ�d�1���wƥz]�9� � ��4��gG�#)`��3��8�íU�6w���*y^���L����ʖ,�)�z�:y�()��vTj�Ε�ety�0�oP�%둨�xۢ��6�eq2����U�X�Ǔ.������_D/�akȻ.Xs}-��Tg�WJ�Xm}8sK�&f �T!2P@Clsr��'��E�R�"��n��br�%�Q�D�w�U_Qr!
QK~ƿ�cJ���n,�M���	5��� �ʋ
��F`e:Mq'8왒���A��}��e;n>r�t��p����9c���}N����Uˑl݋t2�gL��3�/e7��ӝҌNB�J4�5x�k�c�;�M��Q)Vف��mN#�=�]�n7���������ͭ�W�����9�e�nm�ζk�k�yg�55q�9�&۶��M�m۶��y���q|�u����Zk��l޶qJN~@�����m*��)�J.����u0�Q�m�(%���Rǩ�'{�\�01X�f084$$�"ĝ�4JO�Pp�G�I�$�w�����0��_��d ��^�ԝ1yk)�RG�~����ӀK��7��p��ΪxM&>�
L`��3��%�ǯG��I`t����x�%�0ݎA�R4Z���s�SS�1�I�>+�ibB�
�J����
�j�.�B��ƻ�R2�����m6Z��3�����B�:�,�0��|���/� v��R��'Y�~V��^�0�MЗ`���gg�P���f*X�N�KK��$G��XցB��D�ᧆ�Q�؞�%���(� ��̼�L�-����NN�}I�̄g8V���6�D�|�	�Jrn��$J�Z?R��P�eS�J�������Fq6���H�c�n�\���u;<4�9�{����M.7~`��D����EgA�?��i��5�L��C<��O�����h^��)���H�Gh��F�d�ݐJ���yG���?%p�~N�$�s��K,�sҨ�o�����W��^��׆'�jU�N�촬��LC��rB��n�j(#Z�^�H�"�W�+�E���t��[�� ���T�K� ΀���[�k�����.��M��*x�l�R`�W\S�#��C��h��u��������b��-�j"A�筩��.Q��dV��ۜZ�7x�{ь�vym�4z����?av��.�q�aj��HI���@,�0�n1\�(��?c~��@Z@ڗ�)��\�2��P^����Y�i`����m�����ú/�/����w�&pi�^�F�Ǳ�� w����c��)2"3P��z|�kM�>�s�A��:���O ���۾�Q�`�M��	��]�k��ݶ�Qo�Y>��:!��zy�����I����E�KȖѧZ���ܗ�&�'���zi�T���%�m�	2)1H�q|�y�TU��$������;.l-�$9��h}�9')ɍ�
�2���)��7�hUD ��킎�8��>��	7
��R�������2e��yvs�L�������)� ��D�P6�˨n��4l��zH���(>c�Y�p��p�. ���e�Rdk�v�>H:/���h*o0�L-�qw$��I�,Ɯ$�2t��VB��-�?��;��o�L�ec�7��Մ��:�PH
�c7t�
��7_aZI���3�r�x����1`_�n8/Z3�p�
"�"�EZ�?q�x&U��>����b�WrwIn敤�����i��Dz0&}��`	�ڔ
Q�)��|Z��r�����@���G\B0�P��p�%A����Q�Z,
X���)**:����	!�y�A@@��q{�w�o[��6pubg�k����`���p�rw���ntz��tz�DEc���8��[���3=dp��rȬ�ߤ���n����,�n���gŗ�$�Πo�ۭAx���O�)@���y`�O�����#����9�KH74���Z(�͠�5�ܴ��YF�+E�yM��wu1���X���zM��K�i�������s���4�=��AB�">�N"��gI����S�����r��ں�vP:\���>�x�ߍ:��!���?n�����V��ۓ�)��QU�����@�wg	9���
�n@6�
�2��6�DƠ�ɘp��֋��B�}�u�vi�W�u,V
|���7��L�Nh���D�����RA^^o�R$t�9IP̋~����
���/��,+��?�����"FZ���6�����~2+�i|,�6�n�74�x<��&0��a���&C�4wrC�sp��A�a��4��O�����Rj��'<+	�$Pt���fޣ��2?���ϔl>oE�x��f�z�Rc�?pB�y�}��S,��î�d�,3�1�W����#�����/aqy`�H���~v:Q̣����b�k��Ji�Om]iΐw]��G�d��#�8���s��$r����`M���ٳ\4(�AC�@~�NEA~��a�Ԭ�8������L����dPgAA+�AG9v�^g�i1n��je�ZZ׍kY��~q��QQ�-�L熵T9��$��frq�q_I��4r;�8<��B�F�n\-�����<t��=��8�=B��� �����h�R>~����Li�:�c&��s���w;�'�Tf�aq)�2r�c���V=�^����Tq��{��@q;�!�b_��ܑ��b����Rn��d���u#��9�|�q��8�4���ʋ���15���������:~��jM�����׊��y�	��߃k0�S9���T�}-�Z�ӽ�)���"��S�}���!z �e�ܭ%+����h��۪V��T�hx��D3��� h�C�(p����4)+0�����q���+�5/Ζ&"pD��q@2�S��o�ɖ�I)�M�r���H�a=�V@Z�q����{)�H���?Fx��\W��-aF���?��G�#u�x����Ɲ�ISs`�W`�-ԿSIxj4�F%{�ŔRC_���O�X�T��bP �ͥ;t?a���Sk�&R�Q#��?܆���~�W*�E�ɣԸi&),�R 3�M�=pO�of?�Y%����-���v�����p��`���������LIDZ��H�/����ؾ��r��G�՗ꍍ�q���5]%�5_�[��{ J��>R����G���>�e`e��q
����>�����f���Wl��bEu5��b��te�.sn"�}m�CTM�U೟R��|46�ϓVn����7�.���e=��W�Mk�"��[{
��H�h$�����|�6R����W�u��������_�olŉ���^�d�t��H6N��.���@pI��,��Vm�w��xWÈ^�CᬐJk"&ٴ׼$����_���l�l�NeiuBw��.�l-A��DŚ��W��L�K\�l�/����a��#������J]�%��F�N�Ӷds�N1Hy^�"3��g���K�4�)W���;�X�=�\��j�(^�6��a�$�,l ����|��uth�:�4�Z�?�R��	��z�~>FЃ���tv6���a�R'�H���U쮹��%Ɉ=X�����𛇏�������d
ē�a��2m�Q��IK�����٤�%�n?15h�y=;��^�*��%F�3a��bˡ�-o�����.-���&̦�߻�f�D�l����:�
afb����Fu�o��7�F9�^�dH��x�<�?�BpͿ~ge7����O���̶k�{�����/��(W�Ъ�������K���:�"�9x�z��xې)rL[�P�_�Z���4ߖ���r6�O#f����?%����[�#\ߢ�h�t3���֔���bRj�I��Jz���\SP�q� P߫邸
QM�I@������0c�cPl`P��&T�]zH���(����p�4����C����#�w׊(e�Lod����o����/��5�V�O[]"�)ay�jθ����\��]�X���Wt@�.�ؙs`�te1G�ʾꈃ����kpl���J:�U�V���7��֞�ˣ���+�-֨�_�O���+�I��>��2�N[ɵY�:����<.0��έ��*��U6\/�X�p�./!-qP"]�R���Uƣ �F¤=?]���?U��z�����+��R�D8����ݡ�����W�:n
M2W�s�Ws��[Z�RB
͛>���#s����Q���
��[�"@������O��0g�8�eI*P����y#��?|;7�B!	N�Su�ɞn�f$���iq�L_C�DA��������iւD�z�,6c�to� �����O)IFf�[�r�=?;�?�u�6��R3�?>�:��߳��0�p�l	���ޒ5����?��P��v�dR[��*����BĶ��
�i�#0P
SL�`-�NxK�GX>�����(�###1�ѹ��̪����TA��㞦�\�x�@�B(��ک�}^ٴ�.�r��k���|YٞG�P�N"| yL1P�H�dp��������R�[�3
��0Z��3$jw#!����#;E�g��P`:�#�Shv�'��{��r��cླྀe�t�T]�I�j�Iկ������rF���o��g�����p�Pw������`�˸�C/k#QZ��m�i	���<�\-{b�����3��;wɇY����4��7i����/��͗��.�WU�VqC��pJ��������mT@
��MN,�>B�0lZ��|��zy����V�jzt���g�WL��^w�(U��\�bd�B����":����{ȵ�����OI��fmt��~y"c�FD2;i_���o��k���<�\~#W�ȫ���P����P�TD&�f	teή��F��s���X�Ng6/Bt��*�pn�U�1}Vݭ�pL�y~u4j�9�$f���G��,���:�~�/����UR�d��`��x�^�����п�\��z�@O��_����~¢���Xp�t &r��,�F,\/ d�e*�ozo���?4Y�ذ
|����.�8j�Bc�-a��3����*��K{�t�����j��{2�~��XJ���[`�y���Y����]��7����S��^��c�����SM��s����\����Ś�e�\F���0��F�k�T�k���Z��`RڣGǡ�z ��/<,�Q��9�/"]�kL @ �n_a'�D�����Ѕ�^V��N�Mu��[ѡ�~�B"}�0S�]F��$�κ��(�̱ʯ�-T �I���d`s�*������w���sy�k��9Tr��>AB���߹8 ����sB����j�5b�2��Zr�fK�uv\�t?U��Rȸm��z?�����Y����c�Y����qڇ���͈.(��E`2����pL�[�#@�r�P�\�w~,\�N�1UI�ϼ�n�8��e��T�98`&x����:�I<1n�RGC�7����"�4-4>��#+~ѐ�.d<_34���AgX	�� �2��Y9��${L�56��禾9�9Lg?QbQ�WO�/Rj"��x��.�kGo<�E���[㑚�����_���0% �G�� � ��1��o��r&R3eB1�#��#9�h��Dsp�d���,��$?�9�29��>� �
Vt����1ٻ���y�(tz$��L���ɘr�Z���/A]_��h�j��j��h��|'45I�K��B@c���Q(�u��bٖ���@�ȷ��$zژ;�-��T������������uֻC��2��c�?=^leTm����#F���-��{۵q���V�cq�`�3ۤ�⢴���������|�Ƅ���0��	���������\��y)�uW��ZX�F��	�,��rѷ��'��f	�(�]L	�X"!����R�M�15�`���\\���B`�����:�v�*>�Q�:�E�TQs\�`W�I(���1sy
�I����n�&�^�D��y5���n�3��_)_�]�(��(pFj4��,�G��j��;��#j��5��.�������5��@9�B�uN*�JS����9f�1%�T�z=���0� .�8+H�}9i�h�7�^��a4<z��)oG��T�X�_�>"Rٓ����S�����2�fSD��~Z#r����s��A�*JX�`�y�H�9Ft�惻�⎾f�zO�n_=�k���w5�G�:�$��<B�˘
`0>�`^af��T6�à��9��o5�SUs�"*��
��)I
�~�tDL�_��Z��|�v�d��p��݋�4��B�011cQ�rx�oȥG��Y�apJ^F�8�&2Z0���<�]��AoG����U�$ǿ��zƸS�v�g�E	bH��ptļ����o�goOW@ ד�\����p�#�x�g��32^��=N��D��}�g$�?�&�i�Z<�:jj�qp&��Qx�+)��5%��:��zO��ah��fۡ�Kg��ϾA��-Ŷ������Vq���/�O����zC�?�����|�	)�^����t�ЧU0��'���AY�fYъ�WR,��TW�|�;���"xF_nJ�Q� ��N[NBeS�?��!~��ah>E7N��@qz�|"<D�uf��zf��W�����T�o�a����-�y���ߛ:��`\�g�w�R��^.��G����^��n�Gx��bc��E�I��ڃ=KO�{�U�JG��U:YA�]j��S����(�0���BȽx���M�L�T���P2�WM�D����Ǒ��vg}�a�'�5�U���k��Y��*M6+:�+�
�KE���6x����;�e��v���!(�ā�uR#���63��G׮RKL������ԁLi�Bߊ�<�2���T�0k��	lN8�����
\.	5oxK`�fiv�تz�^�HG�_i$�V��i
	py����w�e����!��n2�Y�hR��?��ox�#.�7p�$���}n��NJ�l��:z��t�{�����l��iB��o����Oeh�࿓u��^�2�
v>-�{Nf�9^��`>#���>�]��U��GSBvk� ���,��5l�h����w𐝪�P�E��P�}g�$5Ժ"�����A��[~N9~?3��61�E?q3�s�|�\u�J��g5:q��oʴ��(ȕ�ש����mB��d���w�S�������Y![u&���$�5��'d���;��[��C=�R�I�M�Ƴ��p�+��c��SDJ9���<EF����� ��D؏0		����ӽ�����	+���&C6�Vd`*����B����х4��˝$�oV G�����'j�
B�-�ܼm lo}`e��0w8=�~�k�h|��]i��Z(1-eU��;e����a�c�����f�<2X�P�sim\��W5���D����w��BҝW��>�F�$�Ĥ(������\�ݥ�14hb�T����e�!Vٮ7�=�ɤ0��)?u��,�F����(����ĩP�R�����`���$��J+���˓�B 7%U��㤞p�&�=K&��'[�m��qL�h���[{k�W�~bH_�J�5�;A�8�ְٗקU�pr}�L���3����:��e����g��"|���A����*���K"q�Ll>�q��+f�T���MFK��Y�{�!��(�T^
�^�r������<����%��E,������b�)'5-�Ƈ�E��.?�,�fw	��5R
{�vxxԷ�bq�D5!�oyyY3�H�����d~�>`oi/� @�N[������3o�JI#�HN j��yh�܋������hL,evT�uѼu���e�|�1V��|^�qy�����qQ ��h�9�I�����	ʃ�Z��"z��#X�h۲�ȏ�A��\�;��!�XJ:�YrHe^���hJW�h/��J�]K�m��,-��5|{ȃ�,Y���#Eqp~l�?-\RM�l�$���gP$?��~d�>6v�2�Mfe���..�� U�mc�o�OlY�k6�Z*1�d�h�a�n�N��gC�+��b/ˉ4����ƥ*=� �l;N�o���h�5�!�ik-U�Z�<0��%��&��
ʯ�0,?�,�Wټ���r����W��G�Ym]���b�����Й3�h�7 ���7���G��=&%��rA1߃RyU��-�"�`�"WMyw3֍�)�DIB�����t)Q�&1�������č���\�x���R���t���m�c=-���0���ת��cH�{�<���T�2ߏ5K�Z�u�K����K��D�[���f������zJ�J�L�~|��A�>:[��k�ޛZȹv{�����,�&��Z@���-t�:s�S��j���!�q}���LAQ�ÃǦ!��N!}�W��̜%���"�L|O
bE���kxjj
�������x���c�MF*��L|����u���F��<��G�/C1��UO�fk$*����6�ƕ
1��BU_�E���S�<tek/qN���V��,ʲ�h��`sp�Z[4�D��",��~i&k�9� t�_{�+�V��$�*��H�����	����h��
��G��6�ʠ�Cl�)Q�����|��u�"�:C�!��'M�)�_���3~+#�[M�x.~&��ؠ��c]}��04��s-<5��Q��|?��f�:4D=��AIq4G�
�ZlJ�a�����l�t���GXS�Oz�	8#�WJ�5 �$�X(J����1x�Zy?����u���=��̪ɗ��w3i�~Uff�Ͱ�$:����L�ç��T_���\G,#V��M�/��:��o%D�g���,,m#��.4E��YR	<~�q�ϭF��&T#�f�Wb6$E��$��%C���R���E���'O�þrjzwN�1jV��Ck��HS<����!��/�(Yz&F.��@b������W�P�-g��eeh���D��K��j�҉����d�|ͮ�A���߿4�e�����S̝�S�q��릛t\�-��.@���y!�p��0 �����c㤀?��Dv�@��!�|F��-+�ɕ֢�]f@=ѕK�G^#�:]S���qĜ��|¼=���?MWX��
媺'W�������$�[��Pt��N ΢�q�����"��h~2�3�ȋe%Q[�����9�&�
L>��*06���,W�#3p|�1<?�����'�7�]�������i*��	b� ��PKԌ�6�fDItW6��"����X�nb-*�@�|D��b\��c"���H�Q(XM��m�Z_��@�sp�>#�Ӱ�+<�T��a�!�{u]kB�y�P���8c�E��y��aФ�K��*P�A�r��d�Y�)iK�er�Zh�6�ֶ�)#^�sd���M6����޴��
RN�i^���+�z�����V!���{��8��w��V�	uUXx��/1���@�jx���ƕb5��so6KmĐ�:�b�����l�>K��|�U���u������z	�{;���z4!�$K�+�{Ow[�l��`��f?��%b��^F6��H��s-�/���m���цۖ3Oz�Ӧ�l��"���ë�J�*�N��T�}��R��Vj�x���3�]����I��P�^�<cP�*~.�Z�T��F�}�8L��|p�Y������E�~)�o"�Ʃ��">�r�l:�H*�v�tk�Bo\���8�dӊ�w�j�+*7�^� �	f�@f�\T�b�W����.<eG�d'���."���y
-J�;Uq&ki��{1'�8j7{	&��F�J�U�K��eWC��D��Q�����6���|�@P�!MA��"���L�!��1��������FT��4!L5>��E��yW=���"C�*���$��� ʣ��)��H���1��`~>�0��!�p7���N8�#�< ]g?�-x|�E}������@�{#U}ͫ������/���a���x��xk��947Rm�Q*oap����5Ŗ�e��?�A�XQ� ��R�_�[2n��A3	�F/sp�ɖ�t��d���P�):ڙ��+�S ����S��z(�]=(\WRT qQj��"��u�!*-��Λ��k~��~���\Qi$8X���FY
��dW�ΰ�#K�e�r=���Zns�R-׬�ЧUG�T�c�W�H���lɷ��t`��q�o�e�q7�I���!�8��n�~���#��¡E\4��l�@EV<�"\���b6�R��� �X/�+�3I�vDM�¿;/R�5i��_IՑ�h��͘�ڀ�͆�L*�����y������o�f��f-�{^�G��(��y�=�Y��QN��T���i��3{�@�������@�v�bcJ/A ��uN�r�xm��ߨB+�`�q<���~⩏�h�4v���F�,K%����W�Ƿ$=��5e��W��[DX�T��&�ȓ��4zB<��M���(��Jyuj��6�̆��2�U�4-q�\�/t�2�G簡��%�:�(bu�)
cNԶ�C;Y���.��0֜&mG�z~SM&��qsg�D�.~�0�|�/���|(2����-��M�#B��߄{�"+WW��xN<�8������$?<P����[� �M�[�hJsh�y*�[���C��~JC��`���|��x����F�q[� ƨ���&�SI�99��$ۿ�HL!��Y�I��,�u�
�O�I�e#�x���(���վ1;�F8Q9�~�^N-6� �6�
灜���]����퇡p�N���Rt\}�
����)�ϥ�%��]�WD�^O�1��,�%q �2����Ѿ֒�܅�`�00����z���v�����6��oiF������b��"�.y.����ܯ����6q2�OE�  X�p |���Vp�bۇ�2i�3+��S5��ƅ�P:0�8�2����czH�pi�e��fa!C�R2��:�.��B�N��5`B�XP=ḧP�u�S�l�?~�/���ot>cf�A�a[]`Zd!Y|�Be�$������	��a1�M@�>�}�ڊsqU�����������k�{���Z���w��!٦"uv_>|n'�/'ON8�N۔m^u<���_vs���d� `��k���J���q�T�_T����ſ��������洢Fj~�N)��zmB��;����U-R[��j�Y���I ӆ�0�pc`Ma�������v�
��|H��L�h"n3pS��)њWlO�14��*���������9����B61W��{3����]�/�j����͔������{��ӧTό�����K)�p<�N��Y�Ӯf�*T#<�視�yI��%������P2��h[Nי��ge;��d�A�.��!6"�����HO�s��pG�<������!�#aC���J�w7Y�.�Z���f�V�J$S33��V�����⟻M��?���E��@�k��>�X���������0����3�l�C�{�2����<<�"�J�]�v��E�e�5�[ˆV�,�n��g`�%�eO'�?�O)ڲ��<5���'�Γ��pl�I�J�3���s���D�G0��m� ,>i���Wo��J��&�L������E���#��\O��)&ý1�V+f�GM{�s�s�BA7Ρfr�{)���;A�]q���N�;�l������μ�3RU��K<~�s�K^�yI��&��r��s��m��8�y���;R
��&����,����T��dՙaR\��4�m�,O�)8ǾJ��Y�Z��H�b{�e6�L����e0�r��LVd��e����s�	A���>yD�Q��J�a����	o�s�(��C��j^L�HMto���]h����OZ%�v��%�!��� j� ��x9S �����}�Y�O�<���iF:�z�A���/1�M�Џ��?�]lX�c�� ��:��V����#�4����]���x�(9��!C����NvA{���y���os:��~y{�Js�=ݨ�������W�v	�f��&y�����~2������ma�U����-�(�;�����A���9Z�B%sb����7ySit{<!�a���+'J!Eծ���|����e�R�2����t�u`��*��b.ǽ7�];;�4?�R�P@��s���7��61�y�����ѼAQ�C�ܰ��0%�]�xee�!Ԁ([M�TH��ׇ4�󳧽�����ƃ��oN�AK�1��i��<鳄����Æ[��$-�������N�w�]�ERڽ)�\��_�]けyQ��J�
�K�?O3�Et,�\)J_����e���aبE�l����>��Y�'Z3�2�F��U!���A���,6@�/8�D�YcY�SŤ�
.o�W{�'/��ֿ��V���[O	<��8�(�2:\8�m���O�a]�-b#Z&ר���i2���t�`A�v�=Jԅ�a���=��]���5̨]����>�2Kso%W��e�2��gx�?sD�r�Y�6 ����^���N��꿸9nL�N�����~���{(�xϾ�%��?��O�����/��_�L(��ʋ���j�z<����id����l�b�\wа4�?���������޾)�Oe����`Pl�<��0���ϿW��� ���h��O��b��R�k ��¢а��H���ԽLڽ���yA3!�� *<����7�l8:Ce�5�Hm�g�JF�ڟA6�(�®ra�t��2�L�رgz)��(A��?Q6;@�χ�*&���H]߿���?U�n� ���Pщ}(�R :�O���7VN�%� ?u��S�bH�Q���s
��WK&-�0_��·}ΟY('IԾ�Ws����n�Eii��Mb)�U�����.&TX�r^6Öcm^ﮦk����2��zŐ�O��죣�� �u8�T�yQC(}�xpeT�u߽�a���۔����|���$�Z#�}�a^�w�F�+�1"8��i@=�^	��O�:�G�yL	�<{%G?Jځ|7Uȭ����?��A!-}Z�� C=���M��|����Gs��ItD����
�������2�"K���%�K@#���k�$��5���NiOj��7�Z����JR�}�rt�����~T�Ңp�l�m��ҍb��ٳ����·�C�R"=aӱN�[����UĂ��X���[C�U�*����ϡhB��@��GP�'Z��'���28����W��e�|���}-�$P�t<h��r�.Vo��+*�i�%��7(6W&ѳ�
�j�e���F��Z-�k�k��9����f1�l��z.�2���;����!$�yj�q�!�,,�u[F��i\XQ�5#�(P�[(8Ϫf�7�T��a*(~��)M�!Ok����5��m�=�ʒAX�ԑ�����P�_�<>(�e� s�6:��#K��5�U��`�w7J՜m���)��W�G�w�1>"L�0Χ�:�?)L�gN��V�Tz��W�!z\E,�F��F"&�)wXd����*�eʬW�q�S�O���EHAH��.�z�,��t�84�	2!�ñ>�_�8m�i�)�s:*Q,�����p����s!�EuX�� W~@u��bjfgHñ,�v� ��IyҜF:��j�^vr��r����S2���ÊU٭E������W��_:�_���Uc�@�D]m_�RB��e�\F6�߃�9�{����ߛ*Q��E��Q�/���wƄ|4(ywԿw˺�����	6v�*k��ٽ��R�QC�.# c����<K��b\��B �h��vri�����M>��[6R��7��	���(��{�W�g���nwP��3�-����Q[؊�[०��������zW6�揨I��˘�_�s���ƙ�
ʚ��W���vB;��I&�11i�0�>I����4=��S`�M� p��J.�T�~_'�� $t�E��/�&���X��Щ"�S�K�M��5��t��S�bZxw*̟�R���Oifr{�����cրd[�0��fN�o����mu���̹��w�kY�D��+���Ջ�,�+�����[Rq�J��.$%�������	�̈́��S0��\��sC���G��7��&���T̲Վd0H��뷨�Y��_��d�J�o�3%�kW��2\���b�ɂ?�6�l)X-V�E�D�Lsc9)��4La��A�7h�B�"��3l;��T�h�/��@QL}g������o�� ^i��2ٮeG���ꔲW`��+̽�ϟ��Ѥ*#�RB��Z�}h0V��ͺ�K����YW��|�N]<3^�Ҩ�w9�8�#"��D�����	������hV ���ă��U*{;a�ʅ��|S}��(����7��
Z!xw;�U�����u:�
�R�����܀��y<�eY�-V�m��� 3��x.ِ��3�	���U��<�_�_]�4χ/���dbA���T�`��p,���SB@9t���s�i]<�)^*��DPqa�U�۠" �0���Dx�3���}>�����<5׃�"��%"����]x�<$�Q��<�s�A�oǙ0���p�+"��j���ww%\�Y��H�QQ?=�cP�&5��z.?tHG�����J�4=ĳ��Hc�,U@�J���Ww���	������Cx#��oO�\H��6L7B�V�/�u4�F�6�B���լG%�w�����ʱ�-�7��W�5U���օz�VjP<�d���D�G�,u;)|�����`��<��b�6пU�h'�)�}��8���7��n���ⷯ��ܙヨ�f	!(V��Z�B5Q'����ܰ&�g�EQ�ܨ�z��X-�%���p��KE>��y9�K��7m�����x�ko�峌����C�xG���K���ͱ�=��A��Ŭ��mem��Vՙ҂jq���/
�w)��h.X߄��L|�d*V�Im	[k���~Vo17������ד���o�L-g�fX����'���9��p��������yT��4/�t'�T��Sx,���	�S��g�R�O6�|�$���Ҩ�@�n|�5�����T� \ 6��g]~�3�ԛ���w���r��!��r*K%D�1?X����K$o��::V�/f�7�C��64�τAU�LJ�>���T|��
)~�Y̆H1�ۀX�<v&�L*�$x3��H���ҩƢND��<��i�*��)Ș��ʒ9�#7���>�|%��2O�j\G֧����l'��Xe� �8�
M6u�n��q�y:�?��{�m-�J{��AkEA�l\@��$6NN������;�^o|BX�Dt�7�����ˉ���}2�~@_���+\�� �<*T!����"e�ҏp�JJ���O�r���(�1�*-9\�2տ$x���4�Q����*?�[��n�H��̧u���f߯���^�K߀bQe9���
�y�pt�%!�X���eL>�<PW�s��",�se��X�un
yaA��]���!삕6�gK��9&�]����ͱ�Ϻ|psVA���F��rW��?���P���YZ�J,��٧6_��*
n"�"��^)���7��I�K����ܮ�Ζ�%�_
��u����MK�]��/�l�������FߏJ;��׻��^?p`zx�m�#��U�}x HHe|:��\��XH��:��@X8����l��rC(���gg\`'���l_���-F� b����x�D��#� Z�,�����!`߮1Ɓ<��.��zp�;$�"��җ����s�66���Q���AV�Ɖ�V��N��A�hl����:��r�t��v]�s��u���G?��h���X�쀛bZ@e�s��X0��y�N���wU��������ys������SO�7��,�#�ѥ�CW2|�K�G��0��O1����i��y��	��f�ޖ+b�k0�Vgi�ʲ2��'M!�F;$i���c�@Ϙ��Lrik$�؆��,6�'���)ɠc\X:_窩f��ռji��&hxH��6�ck�3����C��:��7e�5�;Z���6]�`�ݥ�t��N}4-�C������9��y�k���,���-��(�c���?�"�̠�� J�,R���bn���`�l��|h�y~Ngr� �7�=� '��*H��:��?��X�P�>K^���B٤g(����D�B����NG�a�X<���G���z����;��@-/'��-cӱY������Z��)�5��T=�7�=�w,CT���
�<�����R�d�c/�VG��G!}�B� XD��(����'9�ꇶb��>� i�J��õyC=�d����r ��؅�N�[;:a����y���:�#�=��4e�i�|W���xL�X\8;^Y���%��T�c���(�{5�iq��I���,M[B��+tu���*�i�%��qn����/I��(��j�5�T��ߵ88:��NΠ9�JKfyf��/����}��T���蟨N!�)D�+w��APdAw���4Z˶KUz��8�ou1�� X+y�HY���W��k.��3jZ��#Y����DL11�7C�����;8)�Hn&��{��@�#=��DLw�9M�bH&*�:m�
����:��Th�Pzo�z�}��g�\ِC�1w�t��8�7�o�C�����!�U��N�����j�eq�-Xpw\�5܂3hpw	� ���w�����߹Y��WuUuu?Ð��#��;��Y��g$@��pg(A�Q�L+����z��:�!F���>���}���ʍ ��c��t�����(��q�y�������85��au�S��Q3���.�;�+�jU.�T�4�!w:�ϣSl�l����YKO
��"�6�T��[zf���z<�g�s�T
�W����_�*�s�rs�pk���U��G�I���%�S�����VX$H�m���{w��< :.�P`WG0䍿��&!=�9,ɓ�l��DW^��~.X�r�a�t��g�$U_r������^)]|$����ӝ��͢O�^k����^+���EoB���tMb�xy�0�3�v�����`G:R�۹c
Y�m=--�[m��d�2�Bf݆A��������2������["uQ�l�A;����X�H
�j1���8��S**��4�,�"�L1*�j������"��<y��X-�P|x�?_r�B��R�ݢ��<"d���ەf9��=
��j�R��T?��E�rs�~t:����t^RDͽ����9h���&/[�Fo�������#�U��`����< �Tgɗ���yf-V���o����,����H]r���0�~��K�D�u�.��^��Y��İ��w��L\f����7���B��9rⱸ�Ø�rF���g�.�=�tҥ�.��w�J�Nѓ��2�3+1��b�&?Qd(� �.���9.�z���~��.�z��>
�tJ�UV�{��5�ד�㓇�������U��s�d�Ǽ�:���/�:j�P�A�pq|�ϑDϾώ��dz{0m.I륯�7j����z��0����#��0�2�J��JX���p9I]|�����Ͳ�Ƿ�����?��-w����#w=/{3A�u�a��Z��u�b�� s'逰0'�o
���9��x�'�� @���*��IR�A%YtU뺲��TB	��������5�=�����b�T��],A�U��d"x�% � ��MF��R���ʾ������y��8����3j_q�R�{���?���t���Mq�N�<v�rA�M[\HW��~�x��/�*�'ʄ����h�t��%�.ɧ�����T���a%�t�ҩ�Wr�h�@�0�Q��+���D�"����~���d ��Km�����.3����/�<<��<n��!�=m}J�n�%�`����W����K��'3��Ƕ:��Xb^;�������Ƽ�(4%_���0m8��Z�ΜQe���ު�6*����"5j��+@{���"�~��X�u5�0/B�����@.�U�����x��xԲ�!�-���K$f@�8��'������|��xы�P�`	X���h7�j1A~���8��!`N�ڥ��7,�0���	��z�[�����"��,kD�:�N���t�
�A�Ir�&����v�W�1e�1/k�@��iw狵��j�������S토H��?r�T�?�jT:B������3@D%M,�=���g��6�N�?�N_���&Wl���m̚����I�LLF珹?����Cc��-,�c�S�?����$�Uי��eA;�����;D��~q�ȡ����a���P��0�,�7�`W��{v��ߺ�5p��F�Q��Z��o.�}"���كW��Hl�3Z�!K�ǯ���g��@B�.�Ǘ�:�U���\��)JQå⏥��K��א���i���4���c���S1>�he�j:(`A �Q?rJm�����g�](����c?Ӎb��j�ۯr�Ʒ��C7�����?��A)��P_/=M�v!��Յ�\o��r_����ڲ�Hr��T tV�p����O�񲞧$lXQ�0+�rI1��9�[��g��Gg����6��@�$�4,��y�y8XO-	،���vG=��D��ͩ�E�z,��a}V����(��G�^2�/��a���.�o`�P`�Nj�V%�T��;�TRV�e3���b�d�+K~��I0��Z2��;��{wP����ڏ�y��6�i\����l�	�Z���#�U�.�����ǝ"���\~�p�\I��
͋�b��.�h�WcQ��YK�c�qE�\�,�e�/,�^�og~eɔ$�J�a�ߍmD�fw�\t�GG#���{?
s�|$��昙a�k�u�̠Mv�"�����ySY�QCP=��ǤgU��".X�tI�gw�z�|�	���o��>z~��</����DT��{{L9�yR�;k=���~�x۲�B�/#�U��o�����ު��[r�ң�"�*��P.ߏD&"9/��.�y�%?�`�N�dy���cJ�n�G��	y�%������0�9���ǔ�d�$��B턐�G>���0�v�
�"PH�ty��-J_�pW���Χ�H.�%'z:I�'�Q*�-š�+�B����+?M�C�|��v(l�@�|��oN5>��k�5,OO���f��%��3(�^@A�C|[�*fU|��*�g*���E�s�s&��=;E�ã?��P8��Xo
���S�4��A��D��X
eZ�n��ĳ�DE���-O�EƎɧ?x�}�O� ,���/��j�̘�����)4��F���٤>%����S�()����U;�9#���sc Λ�����g,�'�o>nk�3��â�p |�v���+�X$�L���;�e���e�V�;�>d�ܥZV۵�4�������ouy���	�K�-9��,�%�0m�����,>fz����鳓�.,r���ɭ��y��g0����5:��ӹ�l�Sτ��C���I�����s֌��w�O���V&��	��頇ty��B�c&��-�tw�˼�BZNY�U�l�uAuL�i�����#P����vI���ˍ���Od���K�?l�>��ٶ+M����D��D��^�^5e��Cg+�؇:�|�3��3�bG�$�P�8m�� ��T�.������9u��|��H8$����Q��/��-7���ԋ���P�j��Yۋ��Q'aK�����r���$P������U�VVN��M�*�
x5Ο[���o_ʕ���jU���洽)A:�X�����Pm�I�z�b��#�bG5��͇�i���_D|��s�7,�A ����LԤ���
��I�C����6y����0��b�|<���u��U| ���i�	�6��ǜ�Op^Y��\޻P7x�����E,/�=(��c�׊�:YA7�ĶF>���9)�oIb��	QT_��g��PM�.㺵�ZJ$��[׹�鰫�O����LI��a�:���ֵ%g?�6��?«�Xhȧ9m��
�FF��$ڇ�!��:/�B���SR�P��f��h�w�рRry]�79�VI� @1,�dV9��܉J6G@��e}�^gy�V��(2N�����?�kk�:r�g=G�U!J,�S��og������	s,G��3]q�_,V�T�
��?���g���Ò�|;�����f�^��ENTz�Q�st,
v�T���+w����>�]���V}�~��dz��S�o���@'H���1��3���/�z_�G	�?&]�;���ի/�|�`8��w ���ԗ�9�$K�����7���+�[�Dцs�qi+�؎qj{�I� �#-�e�� (�#�����H�������B~
�#���_��o�Mbf�n���z�u��Q�T��q�O���j,���!BIA~�;|�c	��گA!.Kx5���Yx�7B?煂#�˦��g�>�)k�g���љ�/����uu|�n� Ar��ߚ�����ԃ�;��x���N���1�h��+�]���z��~�oӑC�⍀2�Q�Qd"?v1�3�NA@|�	"t�߹�=�\h�,�^G�8���踿c���WLȢ��z�EM�����C���Y�]�N,=rN0@9�ƺt��;�s��$�`������w�U͑|3~�#L��)�����M�,&$;7Fm�3��&WCX8���C�xg�ġϖs8N���"��3�1
��{{�Y#�׽�]%����$>���mu]dɐ������Z�!��.Rb!LI��b�;YT��b6�N�y�ٙ~���嫇��pһ���A�|���:b���ط�<XdvK�&i4��c��M/�wf�$�-E�!�ۘ��`8� ˁ+uU�S��ݏ�}�Z�"��L=g���9��|C���lICS��_�sޖ�d�m�V��u�+�9���I��8p��@wj��#�%	�?`���`�|`j�=��9��4'ˎ�QYY�~Z6��A�O�雟�Ds�2�j�;?=2ͩ� ��z�o������c� �����N�5�K�u#������ߨ�F��q��=�E=�¸�p˅�D��
�� {�%���yτ:��">�L�ך�Ë�x��mG�r��-Mg�_h�.����G�t�����������8"/B<<���0�CC���\�R�]{��ٿ������U4�;��?Cɘ��O>��꒕f��t�����T�fU:)�)J'�:�K�\O�`\aUr�'d�t$~���X( �de��� f����HK6+��Q����&���
��N��_����:z}ZU��Q�C���C�\��'&��{��g��ow�4h��c{F�1��'����<�cm�\ݿ�?��_�_ �I�OX�i�@F/3-��z��X<s�zB���;q 9%���}�:��b�* j%�#�	j�;���Tu,Yy���=| �"�:�Z���jFjm]_B�yL\mbȦn��qr�r�?�jd4Z˭QK-�-�Ӄ�r*N�p_z	�3`[�e`���K�6/X*v��Yܸ��=��1d�������s��FX)?y��s�6�qB������Q��d�����K�H�ٞI���|ϴ�*H`%�3.��"���r5' '�җ�wJ�V�I���U*-TQx�cc3��j����B�E��\:�/��!3VıFd���K��&"��;+�_'/��)~G�	��@@�,=al�z�G�7k_e:e��bmY�D����wˋ��L~��I�ph�%���*I҈�0wK��vM����7�S3�ӟ)��#��L\nV./�Y�+�%���É_��}�T��u�בN�Ι
�@1�[�g&�R��04�?I��Z�!V���%�V�Y�%iIV�A����䷞�Wm���E��>��[K�n�.�Ѥ��L\bc�cq\4��������w�F������\��nf��_+��t�玘�b�D����E��z�04��_�c���>L}}	�UK���b�nDz��!�NB�e�PfR�(x���"R��?�F��! y�K?D�4Zhy|����vw��RdfN��o��qK�ʭ߼m��w�^��L` d��g��
�3W�U�ؼ���(�g)?���0���h��8�JR�`�����7䒳��O͞V�Z�ZBC��6\xt�������5WֱO,ֳ�ѫL-3+`wj5�/gg����ؗ׵-�x�}6�հ�W��P���E��KU�3�L'{�����{-e���0�&��t=[�����Y�(n�?�C#0�RŌ�kD8��Y�(��^m�*��z!Ds���!bfӤ_"�O�4�y���K��N9:G�sI�)NT���۔fkx�,��߄~W�����s�YHZ�J��u+x$'8;�&O�"<˹�d�;q�2pk.�\�	�<���ý�6�������VX����a�Jp}��*9�� VF��b���O��qV��ɕohc+�V9��?����e��F���b�a��R��t����m�fĈ���/h#&V֡g���R��Ʈ%�����b\�;̥�c����;��rh�����<��4�j�ʅ}�\��^/�Nq��C �nX���K������zM��I25�q����M3K�jz�U3�c�o���G"NY�k+�&�lZ_���ˋ	�o}����Εq$��RVf��;�V.�f��d���|{��6���KlAZ좺dm1>�Cc3�7�1��Z�Ii�#���s�v���̖o�*���AR���ɇ�c�q���!�?���\�ʺO�����Xqi�Z�]��a�~�R����q8D�2��r���&Nbj�?M�_~[D�r��ş>�Y���Q/�~���n=��e�%����#�� �0MH&�q��ͱ>t�e��*��0���`�b��V=��Y�"3*Z��\F5GR�KK0�����Eƶ�l���Ѓ��Gr�Ǜ
��9�-�L���2��&�B�����л�]�Uؤ)#���|ut�:�����L8F <jt�J���9B�ve���\�~�����SLL�{bc���jh=�?����F+���|��IE�/�Ny�%�^ u���˵9G��U�SL�*X(@���P�74�'���F�c���)^�>�Hd�P� �i+0���n�����ʚ�-`y�Ь�,���g��iy�;� ����'�;�nh����ۈ�7��ē�بB+�soi[�+_)�g2I��������ܳHd�lk֦מ��lt.7P���UK=QZ�����Z�������0�W��y|��|p��)�tQrHy5�Ph.��V��_<;zBp�C�^ 0��t6k�m:�1�Ք�Xo��29��	�v�X��Tk��Q�H�)&�I�RՏ��ܷ�|��2��xҟB�w���\����7wN�kn��cH����
W�/�H'c�hI��b�tly��Ӷv?t��ly�7����Y�$�R�X�k �����?�|�_�T(�8�(.�
:���ں��{�5�+�j�J: �B�&v�1�0���lu�Hm2a�W�1x�t͕��������lH��A&�YI�]!d�7��k^666'4Yr�����/���_�m"��NMM��W�,.J<��z�[W��~�8:o�?��룆Ћ��3G��t��������m+~��TO�� ;	Y1[
�܄W��.�u��\�U�B�1�Sa)��A�A�Ӝ�����	��~Y	��ʂ�~�O�l0�b[g��6��OB%�ӭ~�,&�*
]a[%���LW���ڧ�T��:qG��J��"�a���G�H��)�+\5�XT���og�N�:~�YF�������3��ɓ�'8_��ޓ+�<WY�z�$����t���'4���_��>�]�����\#bb��R�&����F3�_u���anl':�ff��i�]a�P	�K�녉՟����rhe�}�s=�Hdk�"�]nH27/�tt$��+���yCl�N��Dz� �1�!�m�/�߼W�Q��"E(}Z�D#��T���U� �;�^ec����䂸�J�]�Ud����>=�1���3n�"���N���1&d��>�}v�`�@��dи`����L�����r<n�ޙ��^�E�4�x`��|��ޗ�)�5f2����xo����e=�ng+��;;;�+�*��*�+#0�F��vO__g�J�u>5}���f3h��}d��m���1���D��7?��2�v�X�fg	~�0���yN�� s�ОH��w��d0{ �3���p[�`T;�B�<��1�z��jי?�������A����DA��R������%�|��I�N�X*�����:��7��o�Ͷ3���!D
�jө�&(1//�����\$P ����5+���(!�zv�e�����r�w�\]�qЗi�&����.T����9mM)��K��4����~N"���]>M*s��85y�Q��'��#M����T@k����gR����jBEf�"�Z�:��/ob�~��jb���-g2�!�|���s�-�V;������m�x��;� t�����|]!�=�2��Q�L�c��� �}U��ͭ�>���R������r5��_�ĵ$(K���w�b��.a���B�,>FI��ݗj�z!@�#0l'�nW<tݗ�$��*��w�e�D�< K-=�=p����j�Yb����p���- [D����>����`��	x��+�ޔ�$���r-~���F�0�ü�<k�³5�_''>U >[s��JL�KOٟnm��=����1�4���m���Fu	�[�,�!!!Jv���#1�_����<����,�G������J��L�
%`��W��k���
�����P�-c�U���C��U�Xdغ&�|J-�)dw�����*E�4�+��@���0�d��D�Z����wq:��F����"ʜ�3xd�q={��t������U��(�!���&�h�,�}6��T1Q�Ao����%?n�/l��s'a����L�Dכ���i���z}�{k��1|������_���� |E�����<��>B;�Űy4E�ps
SU�aqD�,룉��7����8�]F�wq�+�D�b���cG�ru����p�3_QuF��T�V��%���c;Z�/C�jԉ �iDK�������#9M3�>�ns���	',�(8���!e~K�u]tl�7��U�ֵY{B�[��w����+YY5�d{�@V_`��;с�kr���W|Q��y�����*�i�̓�*dE��K�%���%͔�&Wh�Ƌr��*���ͭ��B���)E����DFÓװ�Ty�5�Bk6E�-"�r�Cˍ��a���_,Ѝ.We�Sk�/����?1GP���[[�+��x_>�~V��ΉD�q=.���H�d�)�r����h���ٱ�A��b�D�N�GO���	��d���!&�i���v�g��Y�����:E@��kӃwA�C���'5�C�
��R	ZdE�`=��d���f"UF@��~�&�p��o��J�"L����W��̪^��R�(���W-�X�8Ρ���a'՚(��|������
\���H�z�.����-W��?ߧmr�Jls[%ϣ'M݅w���'�'�Q�Bz.S�>%M���pשfCPV��\���a�YB��}�s�"�*���Z�c�~�+r��A~5�ռ�}.ca`��j��Zw��ƕhN�O�������,��ƃr��tf�t����e�o8b�s��	���QM Sx�hhuz&���i����c�����2�Ox��Gc��ୖ�svY�e�T�VD�B���Ŕ�+���q���&��F�g]�tԋ%���T�����c[��
>�`�����*�9:D%H!f�Z_��������h���uV��޹q��W�/�{�j�pu�7v,�{EE��r5�{�X�dz��B�mՖ�n��\�ˠP
uװj'�V'�sR�n,��j�t��H������:s,�[��,��:8w����W:�9�}���Z�gx�i�uV]	����ɝb�H�UWA�_�
F��r$�)�s�#�U�f2�B�Ԣ�'[��-�Vi	6=��V�;Y�W���l�)=�&�=�C��M+菛�0�C9Ma	��,�F�	�n�u��i�G;�8��nrB��k����M ��J���X��39X%�
t�o����2��g�y�{�V;��:ЩR�A�9!Р��'9'{r�!!�<w@��"t����7��-��J����J#Pֻ��y�Z^}�@�"���/�em�0Y;��táB;�/�SS�Y������G	���
p`M�Rl�oJqd0 ,�f)8�B��Tn�HWX������D�,"�ٗ �a����z�LU霶���L���=���AJ6�H�_�g�l�����C����{[D��Cq�JE�R�����o��^En��!��1-Bz�qT��Qas�_��^.'&G�$��?�oh��uj�*�Ύ�o�U��s2ƻN�-��ݢ��\|�qt�����+�{���Q2������C]L�h����y9!��4� ġ� �2Z���+1�?CȁX����AJ� ~X�WRp��B_/���n<�eI�O�aC �9�L��w&S�N������ʱ�5�ǟ4��+��D9��ٝs?� T����"l*�b�]c�a"f�J��u�����j�O�~�j��m;��8�,�9��Β�G�+l|��h��c����{���dm:Uj1�w1?3��:߼T��v!����s��y�p�����s��NQ�19�]��/���񬯌}H�冝dê������i��:�����������lo�����^����@j��}\���5��	G��⯑Ii��c���Yz��@�Y���[z͸ ܣA=OK]��m�YW�w��������0U�Z�S^ढ़�٦�&~,S9|��N׺VF�k�_�	r����R��"��)�l��<�p�� Rl켌�����a�/�^bp����L�s��>�SfW,���s!��os���R�zP�ngO
�"��1��4���፝�h*?��������7U������l�N���:X]��B�=z\� ����k	�I���f�ܬ��@���? �eC [n	�ʑn�hr2I�GC6R�o�VC������L��ͪ���>i*)q��q���d�-�Rn��P��Ӧ��k�$�(M��rk>��m���DZ��2q8X9ӿ�����c�����}��FGD�jn�'!��(*j}�"�kz�H"˱&�)�1�_T[-d��M5��{�7���I����^��2�@DwG5��h�2���Pm*�!7l��[B�|B{��ТLk�� ��x��kљ���~�)N�j��ßq���`��HJ:J �Zu�\Uꏕ�}��gQֵy��S�7�����4}-˹�9oJ������ S�����{���9��~l��E,x`A{Y9�ۨ�w!�u�k��o'n���F�R<�Ȅ}V�_�y�W�ֳ96߄ηa<���ׄ��kBq�dרb1eڵ��}�J���n�2'���$���e�@,h���_��%_�x�P<( ,P~�~s���*�ܟ�o�R�_���뫄��J�u�;V�҄�ܡ�?����io.~���ރ�bw�S�&��۩���R��~�L�����ǋ��n�������z>���D�c�o��_S����q�53򊃡���@�����߳%7R����=c�����S���*7�b�y%��f {�_���>��x,7SI��+g�̚�R2^�h%S��t����kXL�`~>1�	�NT�e����"�?�~?u?�㊂���ՙ.3�T��˱/@�[��5��u��`������.T9k�Z�S7J��ω`�+`/�8�KlF�?��MTJ6�95J	�ῑ���.^`TT���"�N� T�aM����P�U��S���I]�y���j|s�)Z�V3�#y��p�O������% `e�m�vTZ�^	:��x���]7޾�P�����P��V�3a�SBݏ��j�#�{_�B5zO�}N�?������d]��YƔ-�\�Zk�*l]�R5�s�(�bHB�T�|��5�B�.�f����@��_:ܤ^�zB)+#2�$*��'�MM�3G-ي[?	(#��}���ʥ�sފ���J�9¤��{���
�����- "b|��
W���s�Y,�7��Ñ@�{��G����X�%(�Đ��M��5\WX^6]�lp��z¯>.�,��Α�<y�o�|  �bw78K��|F#j��,�����n/_>��j�H�UOo��#k�>����3/��M�U=�� k��EOb�`�f���:
�$���ϳ��Y��0H�d�c,B��Z5�B�{b�>��<T��_�`�B�'Vk�~�he��؛&�s=I�r�WIʙ�]�����v�	!���<Ǐ�>*LQog�:6]@��Ks<�%o�����z=�*	�RK�_`乜�F}A�9�5����}�
.||4и�Z�$�l��Q}}�W�ʤC�/{�$��?�cJ�󰉯Q��X�]v���|+�e�yib���־���?��ʳ�y���z��Gb|=��v/�����*��X�=���=�B�Jv�r��h�:�K.5�����76[���V?^w-����B�]�y�E�v��UT ��O+� nA�{	u�]�+� �O��M$b$�U��ş���'�H/�x���ټ�h
��)A����fo���Y�,���c>,��3��,.Ƕ��9=UFIE�����FYT��W�Z�3��fo���SNM�o��^}���1k\n�}=e I�%V+W�)Y�bsi�=\��|�|���n�k��ve�
������ �
�:��Ipɨ���?2u����F�<J.�I�����/������ozܩ�8�U!�2��=Fp����f���FLi#��m�蠋nī�hRA�q�*t0ç^P��񳈥 �Z�m:�4yVy��5~z��C�+)�3Z�br�C%�z@/�F5Pl6T�#]�H-bP�&!-������2�
.Q���,5@*��~�Ї"GW>s~�π7uQ�'�%�h������}�/�	Z��7v6��y�
E(�T�3|��R}���ޘx��f��i8,?Όt�sC5{��0��q-G�-�a�d\��?N#���^����ۯ�43B�{��ܛxzǅ�z�s��,qo�tQ����M,^�U�$�>��7��-�A���:1�e�h�Y��>�r�DdX{�	��?�r��a���9���T;���������x�z�/�)[�|��Ж�Tؒ�n�բ&6(E�N��S	�%�&z���|=3�r���ʅs���RP|O��b z��j��'ָ�
���?��<lY2NZ�R��`G��x���*A���+b1����C�C//믄���.��I���n/��d�.��������oO܉ɧZ����O
��oW�p���x����;�B�Fy�~��{�i+T�Ɣ<_�J�8����ɫ��S�G�s8>�n՟�~٣�/�[���J���*+�N�|դ���/��>��'1W)�l���]F I�ʌx	�`�7�4$��{�b�pY���0	�ڗcJ�������	��S���f�EG��z�
W燪�\�� K4�K�(�nu�	m����E��{�o�]��a b9�Jn<B���wq���v8?��	�B�҆�_��ۚ�����'�}�U�0x����9~�v����-��,�9��[��{�����/���Ș�ʙ���bfo�������k��-��7;���Qu�SU��eW�f$��<�< ���0��LOj��^�@�[5-��P\�H��u2���W���n冗V�ZYT̘}#�j��A��X�n1Jn8V_�е����T�)#�#_�I���ʕ"��A̩������sxjⒼr�Β!��1�ߠ=�����ׇG��Zƺ�D��d�����K܌V�ixx�jv{y�s�j9 � ��%���������C����?D� [2b�OU�s�%�G to�7�Yod�=�P~��df�Qb�6сh҄}�*#E������ W�����]��z�[4`�-���o[o��j��hE����ǲi�*D6pv)�%�ֆ)[�n/���~����eԸ|���\�
ߎM&l��_^�Q+���𰥹�	���.Tu�M<�I�� ��䧳=�|X��.��A�PKzϰ�j� 3��M���^��#�W�WԹ��un޷��s���3V��z�4�B���|����b���F����@#G�tl�u��ԁ�Q_u�ex5�
Tvn����:��@��
0�>)OG�HW;4�8����ϸsſ���#��[�"����[p�~U �
͝��OL�wH����+�2� � aMUx�8�Y
���SU�U�����L���U`֦�쬩��{��wKU"b%�k�=�+k6���^=X˩�1��U���3�t	?���N�=��k��MzP�h�{�I�O뜱}7/30?C��D��W��P�*i���e���68Qŧ:o)��fa�����5�-<eA�7�����q;��d��ǫ�a���Gyo��>�=�H�M韸gaAAFe9Ŭ/�"M9�+_�?@��������_����A~��jCC�R]>��{8�Z .�t�Stiv�Ã��k�S�&r^V �^�g@���蕋1f�Q��J���e֬��C���9*�G���Y�a%��-��56]�C��n��R����T��_���w��=p��c�/�����[�Q�����]�ʠ�0|�e\g�d�g�_m�?�0�jӸ���C#�H��Q���7d_�N�!G+��Q�$�1���Cdhp�K[��Ls g��މL��|rP���9�G����,{����i=N��m3�o�t�@��!�@71����O���c:��6<,M$������pJO�4���,�J�d*Ӡ�������|��*a�P=��{c�8��AWIg����c
u{U��~�3DH�2�{=�{Ͳm�Te�p=
�8��
d���˼@���5�|ѳ6)���w7�W���
}FP�b���d/���L����p-[�T"#���~�������G>�,�W�L��j��~���8�cb���~kP�R��ʕDI彺|��CK(F��a��ׄ3��(C($��Ks�j��ʆs� >0,�-��f�83k���'MXI�Q�ﱺm����k�ґVD���mf6����K��M��f��Ev�A�����/��&$%}���̥�_`�?-�="�)������C �ޏ6~o"���ާ�����F�p=��V=�����D��q���KP3`��=|����)���C���i]�}9�c΀�����G½ȭ8�Ĺ�^p�y�|�zչ���Ӟ(�P1ȏ|I�/GP�+6t�am�A4g �^�l�%+��C|�R�Y7��ӧvҸ�Q%ν�qz��C������S���!<@Т��y�s*/����g���]G�%�O�@4,�=+{�)��_��,�*����֥���Hi�d>���k��@��u a0�*G�{W�}�V/��0-g��dzW0M?5�7�7xN�K��ҷ#��k�)����	����/y ���C�/3j�v�OP�J�[\���u�m?\n;�c0��:��ѵ�<�J�}s�D�q�&<�,��"�du��࢑ΐ&1�5[���]"�nIj(LONb�	�ܣ]�-��h�h� �pϰ���V�Sa�^�+��:W�6o �		�*j5Ĩ�q�
F��FZ��]s��r=�y�����V����β��������%���0�M�����S�e�)X	��݁��UMl�o/�?&��]����[�3
�e�gn(5MM#�������s#�d�%^���,�7@�:���ƿF�%�}�2;kܓ�=�˶���Vmz1���QjP?�n���)�Ϛ��wgad(�U�|ty���+D���0��U,�|��B�DZR�Y��𞣡��}�&�ecʹ��8�)Xm5~�D�%�D-E=�s�
`�E�o�L}@�qIH*�l~'S%"�G�u�_d��ZVH�MҶ)��^ǓNШi Q���	���鐕���M>K�Q�ƥ��&(�.[�u�kr���s��pu��#�$kZXī�|�pP"!�NܯFVLV�H��M���m*��ċ}���֧Qߞ�>�:!o_L�Y�!2ސ�=�;��\hD�c�Kl(����0b:P�^�3���9��@����؅�<B��C~��Tf�U#���ٌu���;W��K�عh��%:j���_ޙ�o�}G.|ه-�!��E�h*��U�����B+z�H�,hiiYҹƤ����/����au�x�n�'3����y:#A�s�oo��&���2���'������p!K��e�D�>^�_ܥ)�	�SМ?,�}C<" ����m:�7��O�.iӇrP���?f�M��'��9k���هɐ!g���վ�:���@+n�O{*:�?��/3.����ƋU��ea-���Q���a���jT٠&�]��Ҍ��lj�5��S:�9�g��lL�'�<�r�����-�%[��r,a[a�K�h5JB�N�Mdz��{�S�f�a�1�O^���b��Q�J!�ㄇ�t��{q�I#��:Y��4N�Z�ۿ��ڛTCYz�]�;y~��@]���T0�Sd����@7;�g����!γ:mM�uk1���gS`�7���%��T=1��ȓ��r�Y`���)�6���Q���A�Dۦ�/��]4|�%n�F;5���^i"m@����M@)N��^S����z*��蟘~���\g���W�fj������u
I��$����Գ`��h�xar�h��mQh�v�o轹,ݖ5>�:��P�uoWkҏj�˦5sjk+�������:��ݝ옍���Ic�ܱm6��ƍ��ضmm�ܞs�o��֜��\k=B�c_j�V�~�zۿ��{uF�%  ��;�%���D`��J����j�:^Rj;�h�P��F��fk34h��X�J����������(�^��?G��nj�s��2㲺�ⴅ>%b|�Q���k���T[��ŔNU����x�ū�A��:�/ɳ�kr�  1�S��j���D>����F��<�)[X�[^��P�}�5����a����gG2[���X�/NA��C\�1���@�(h��v��=�>�����6%+�k$&�Yъ+I��fh�����h�Dv��O݊��N�s�;|r�ԈY���H�����z����u=�Xh5|�����o��U��8��N/2�^\�ԌQX-! ���@ �`DX��~��5���� (�܋�}�f��y"L�2�J���
!�5)�4�@�vvz�b�(!=�E��BĦ�����i�����p!M���cz�]ݧ
Bq¿!7ng���c�,R���Y��U��� � 8qk;���l	'�ɧ��ٿ���ev���a~�sP��V��M��Y�Qk����I������G��9k���2W��Ӹ�����#�]�X�8�Q�d��n�����F���
�8�N7�9%�h}����o~���z8��������HJ?��á}�lF���b���`6Q���_�/����ȕ�v�:M�������\FM.A�"ɣ�����`�01�!��R�J��T�R�QL����v���f4)��3(/�W�Au#m�$��J1B�	��_*B� �;`�j�Z@��.W[W<�U�͢�u;��\���T��:1��#�U@�v���
�����@�yO�#���W�s�h�nN�w��F��E�t7p��R;��G����4���yתLq<9��Ų]$�'U�͡F��H�R����� ��z�����nc�Ɇ|'G�>�0��E���>��S��N�^�) �lNA�F�0A��A0���򱽦k��6�H��H�\�ޤP�?�>��O3 �3�Xְ��0^ʦ���7i�"JY]^8�;�_��7��hx+���<�-�<U3����y_F�-��d�lL��qJ>u:�����:�J�6�i�b&7�m7�VK�z���\=)������
(��
�|��1x:[,s{a��2
D��M�����_�_;�4���{)5@���Nc��8�u/W���A;��dL��7�u�ry6w'Y�O�Q�ތEe��/R�ݒ-P:��Uk�8T�I��+ꆦ:�*$�r���UZN��s,l$�A{��!�&�}����t�f+F+��#��l�xG���ܫe��k6�i�$�����DR�0V�rp�'W�F+���:���MU1�3���!�@��Z-`d�x�S#�5f��^ۚʿ9q�v�3�	T�I����K/4���cT���K�
L�¢�g��� T�J2o
����bp�~�M�7�h����)�����`؆����1L������#4 ���y��b�6�^RQ����ur�6��X��F���`Ɗ�G���rV���	ṷ8ɻYI���e��d՛��U%���^�t�M}��d"P�H�,]j`�ϽU
R=O�m8��g\�Z�"��>g�u:rB�LR�/7�4��<�H���վv\�^�N��~������$����h�j��b��>�+�wW2����7SGv�Dxx�jmWy���r�d0���l�o��f�*�`��n7��C�hf���vP�{���s?��T'+;;E^<�*T�x	z��_ϧ�q�Ϯpl�ā3��}^4��7����e�S�S&?8nⱵ�$���L)Y	���cX,7�Xܡ��uD���[�:In�)եT[� 8v�&ې4����D]r�n�zh�]��	���8���>�\���Xb�ۤ���>U	�b+��[>ש	9.��2���N��8r�/d��H��4�P) �Y�&]z��������yt��П�$��Al�/����N]{CqQ<�P��B⣵jE���J{�G*=�U�]�]��
y�W_�[�B�t���N��C�Ja���T�$������eh���⤧ؕ��y��z�aS�h��N�����g�E�8�P�ҞI7�
�d!��B�xS��-j��ܯ�a4��S2�-���z���Ѕ4�񾗫���*{߳Yή�	ߜ�o�$��i
�[b<P-�*�;����|F�>>b�H]I0��݄>2���~�K�kL����0s^��~��.K��Dɫ[�nU ((�>�Mz7ݚ@�!"�^�:��(�v�MJͿw�x�]~�|C������O����'����x��.�R��+��ԛe�a,�r��I&���e����1�?��_�i�uĞ����,B�k@�����d)���`>\*�xl�?i�&���%P��	B{����"�y�������pn���I|�����Iiy�@خI���T�2<)J�y�"�����(��1uM�{�so"�.%�����l�L�Q�΁B.��2�N��g��5�E��)#zcF)冕��H>�5��@���}O�,kc��H� �p����۵�״����˧�(X���,��^�ӞoG�I����@Zg�j�K��ُ��&��̰���<�o.j%@��̯�s{���=dh}6p)��c2)�j�&J�����D�u��=1�c7b���\׃���9d-�?�`������N���;B��,��r$�O�&��{�8[��{ �7�u�_�fކ�|�W�rA�w�x� �8xV����K@
ڄ�0��=����ѯ��2�S��+ψ��&��+\���]��T��Ą
����j�h�D˓��o)� ��LJ �!1L��xn�SӲ��Y++�3�a�w:aEb ,EþF_�K�ϻ�������S�a|'��X��cs���Fm*1���8�gV����Z�=ч��_�c��e�}���;H�Q �D�G�}tħ4���$�X5�Q��>�
��(��a���+e����a�?Vz�����E
�L�x�j����,}�d^��}��F�k��T^\�M�L<�@��5<0����S�Ws��J7��ʓR~Mt���B.|�� �~����ڴ�������C�F
�d�.��LhF`�=�ķK&�Z1C�0ds�ve¨@�����)_ӏ�K�e��(���v����A��8h$x��}0��_������T\d��U+�̥A��;��}�?������/����̵����r��������A	���)XX��du�TL|H���\*��T줻��6N�.��6�{r`x��E�ؑ�?�jd��Ģ��l��|�d�X�9�N��?ϲ�ηɮg�ӫ�����s���o;�s�1�����$B��Jhtl�$9�>'������I�Z���j-9T��5��3��1�'�	q';J��O2�/s���T3x���
��)���$�o�''�M�I�2��Pi���L����o�oqj��� � z�c}{�ߖ���xDx���O���oAŐ����-�8��='�)����H̊m&�f�N������L�Bp
�w�^H���e���
���)�B���)�CN�IM���,ʗ�E�3����͇��;���ۃ��P<����&b�F� :m��3���o|�k���G?SEEe��������>�j!�ћ��-)���hB9`�Ƒs�Hq���T�]�����/Ws	�%4���x�߿�������<wuB��p�(�!�C�G_�l�;"?��/���O�ճwS��xGp~A��-F9�K6��З��Y�|-��j�_��Ö��j��҄����a�E����+c����̶]�s"��}ryg��R�.�zȵw
�&!g[��bh�"���unKꟾ� ���D��n��@Q�~��a�}#�,���P�B9/u��,�Y�^
���]7;D��c5[�Vܰ��J��;�J�(u�;4mJ���y&�uD+q$B�8-�8.a�/ӏnV�J?i "�6�̥s�d�����ܟ=�`��y��u�5��Ơ��˨�O7�>��=�D����\�Q��.�ơk@���dS����?±"K�_�����.9�fw�ox�)��4.]ߵT��ykl��'��Z]]�z[�x4P��� KC�7�
 :�f�1L�u�M��nc"�5�dB������J`d��s���Wz�*30�P�_�\�$�`Ɉ}ve��p�$Z�6�֫J.'��1p�Gw����/ijȝ���a��Ԁ -��$I�5��ϣ�|�o�({r�G+�֕�V��(k(ON��#|�G�D��/��/ֵ�ر�f)鱨���"R}n9�����V�i��|�(�P��p��ë\�Y2�`�2M�m�ܐ���e_K�qP}����9��j���L _S�*.�ˑ�P���Nqgg,�7�D�f��y~�%6h���j)��k0�@D�:������T,q88��E�pc�]k�?�<:��EQe?E3����ŁE�����	u|�M���1d�K:��V�w�)<aA�JD*��r��,C|׽�=�mr��u���!�D��i�XY�4 �洜��o.-]BB�����!k����N��%6��f�쨷��^��)�"sTZ�P7��7��5y�W��+��T$PQ���5*	VwX���z���_f2�r����A~�6d��u�K�}ydl|m3�"�+�e�|PI\n�6Y����$��:�ĴB���g0�V�'�

��#����<��#�v{Պ���k����6{f��`,�C0;=����G"��7B�*�[/�G-X@��T��UY�	����A� �2��ȫ��&_����ĸ0�q qY�#�𠈌�<[/"�^-_��ڷ�I���;��Ȅ��o�l?5`�� � �\M5c�`D3�(N����B(�CAy0���+���%���㗉ځQ?���=C�����?x0U�}�?��1�>W��rv�{ˇ_���|�:,�\�/~��yt?�#�c��]���9Р]�������|�E@$�'fm�CVy���_����,T��~v8�"d� Ko�k�!�ǢIp�������S"���3��k�ɬg_���çzE��sʄ�bvn �v ��Ua�=H��Vus�"�VC_`[�(�b�Yo1CnT�kS20��*H�K��Y~ݡu�*N�l *�~��M{𬟱�ȕ
o���h��3�c�K���Ы���9����_�VJE}`M.i��������	x��_Y`L�㵮�p��j:�O�Ks��8���$Q[��e���m�~�f�JF.�*��e|b��a)���"�eJ��x�� <C!�*t%�Z�9�Y2�2s�H9
�j���� :A>�>��8�S1� 7ĥ&��d��h����Hx�,�zRh��@]�X�\W&1]y�{"Q�w��y��t9���h�$]Q��G�xL�пZ���|Rk������Aݕ�����a�ɢ����c�����o���K�L���q��\�X�%�U�umܩ�>k�A��2��� 2�<+�[�O��&-`���>���� ���.��"!��h�̵�g���>՞"��<׌i�s�*�V����q/�;BP��ׂU�m���I�(d�B|�(�'p|v�Ԣ��2r�%���@."�-����V�5z*��������ڋ	
H��X��J��7_��]A�%
�XM�
�4S�^�<�ہ�ƩH���Zީ�-�}t��c~�n"�[�p������PVs������@k��o�h0�󼝑�v?_�#lo��x�n���K� W��ק����!e��r9W�]�P#i����)�Wo����[x�M�f�Y��B?� 3�����4�jյӊ�� 4C{>52}O�N�g��ڕ�K�N~�j���CمRT4T%�&8H_4␪���V�w@�3ǡ����-������]TB���kj�g��|��Ǜ���T��&�c�G��iW��ǈ�Q����	�8��/)W���E|�S���=�����E��ї�����=�������6�#W��?61����P7��Fz�,���8*�u�m�n�}�4W7��"�]>��OW�Ϡ��}�e�d'�p2�G 	s�i��	7��>i��v�2|�=j0��]��05XF�D�����d�����E��H�:��l�`��4�3���gč��s+���3����S�TőLO֫��Y�V?;�H�C��GTf��>�uG���kn�y�Y^�%�����������*��s�3��X�=���ѣ�OyM�\�K�^��	!-��Y��m\\���S�K���y~� �:}���	� b�Z��*�D6����	��vL~�i[�e�o e�5+���aڈ��zɷh�O튅E}�AX��G;�E��JˊvX�#��_$��!�R��ヵ�E"�O�ˣ��"_�K1, �!��&K�L����Y�A�f5pU�A�I�L0�< ���7+��
������'��SY�a�r��f
Q��ʶ�~'5m\}��a$��%���"�,ǿswu��i�J�5�����-v�3��	��2CB�-@�}c��P�O�9qJd��]�?�)�S�����!b�¬������k	g✛
9�Nfp+�]�ݣn\x�,�c�� �A�Ŷ^�ok-���pf�+H�~R�`��%w&Hf��z�	�%Q4ݖ�7��=y����#@!�X�r������4��b^��q�o��@Ԣ*�:x�=#�C�V��(((��|��;a���L��ۙ�F��c���ȋ�b��	������:�񈣧��z�b�Gd,t����ù�����9/�؋�祅!MQ�]YS�Rf�PH�Qa*��n�z鯃LܚGYm�_��U/�_�)W̔���&��0F�ӬsLW��P-/�n�f�ȭ�Ḷ�_��܃�ʨ�GS6`�d/�O��Xe]�m�$�z�[��߉ɳ���9q��N�!s,Xϛ~�*җ�D\��
`D��-wGa��� L���@�xY�(�%�<�V��#���x�c]P�]1Ɏ�F�B�P4T��3X�:oT�N����9�k�%�xjUzG�����&��f�\���V�ߑm��Ș+�ϩ��?J�\�%^�tj�;�TqFIx:o=��
�F��m~N�L����� �6=�����~�nAB?�`�e��Jz�Δ��Z!ſ���b+�g޷͚���t:	��+pؤ��θ�M�>_sf��_O�r����W�F����%2bC�kO��!4���eە6����c�_���a�AK�@�V�ۇ�<���u���lɎ6ӱT�����M/kb�����f������(�hM���h�|���ʇClY��.'1���8��T+��dr��J�<xf�p���������%��m�w���?��#��M?<0�}.�T{��A��S�PX���qT���ϥ�:�hD�1g}����[�u@[�:��슠�y���c���z9@��9=��#�ݐ`��oS�W�b��Gk��塽�L�o�6�������ߠ��%����{DNA�	�:��R ���:�W�#�'���Y��������Wic� �]�:�Vy��PW��[-u�4�qm����Z"�)F��X@�(���x�g@��#�	�5XF�&��ᏸ���:}���*���=��}%�+'����Or�P�&[In~W݃�΀:��7�P�	G' ���ݶm�[a�ҧL}��%N�(#�_�k!�� ����_��Pc	��4��{	ay�UbP���Oft=Fu5�ۮ5�ֽ�m��ԃ�� �T|�EswqY?v�X�ҁ�K���ۑ�hJ�'0��j�-�Y c�ohSa�rPgӛ�@�����5��qA�𤕭7H6ݚ ��l����R�͟Aw苽#�,�H�r��*���H�GQ�SF������e��k�1�3V�A%+R�IH���O�[N��0�@\�Ĝ$��Ag�9�Lݰ�K�%�ڃ?S���{Fs�ZV�vZ_38ð�I;��$tN�2�j:�%��K}f9~�Z8��Ӫ���a��3������.�;��a��΁1�RY,�4�-?�yFr�~�*���/������̳�\o�e���Z����/A��k2Sn#��Q���P��:�y���m4�ʠ�+��Pϫ-S|vI5ʾፗU~�lN�"v�]ۙ'�F�͹J0�Xqme�^�'
�n�f���A��Pz�*_��Z�Vɽ�s>Z�]m��XiXZo��:DE�1��:�{Gz��|��7��	�٬Y�����B����2��);�N"e�������
(��c2�����g�-������@��YK
/6Z�:B��h�`J���#��߻Rc-?��$m��#TD华�p��,��M9��c�:oEp�JS��uQ1"nu&g,N�(v�G����.�\/h�(P�Q{\d�"�6����q���W�3$��L�#�����Z�\ �$����L�/�*���.M������e�]�]t��eUIģ�g}��1+#ߗ��C��i<�?�\f���|��2mP�ܫ�N�s�F�վ9�������T��A���zlHCׅ���c�-�_�$fjƖE)7@�C�w�݇@rϗ�l�ԁ�ח�7r�&V՚K��g@.�z�9kq�?!�"x�L��#]{\�޶��&���P��y�/	eYM�g4Ƹ�
ĥ�m�)�_����\W���� ܸ�`�Y�$]������t@��1+_�UV���Y��L|G��H�n�[��C�OXs(��}��5��-|R܃�����#��qAT?�ͮ&^�l�^�)Re��c��͕������һ���J�����7�줪��������� T�2a��8&XT����P�إo��	ِ����o�Ԧr�;2d�_��[-�A9ٲ�A_gc�P�]���.���)���YV 4�l���4���N�/!�49�j�ܒ���R����a $,�)%�����8�o���Ъ[2t�o�Ȧ0��L,`�����!��k�@ף�Fy )�E�G��~�yy�;�:�=��OG4=(Zz$K	&����(^��{��g�gZ�|�����pg� e/��e9�E�̃c�2����b��6a=���k��>�����Eϭ��Vh�`��JB����њJ`�-q* 1�7���*�MF�	��#��[/U�wCvk%G$Q��z{�kе���Ƈ��ռO��M��`C�{��ҥ��A�PZ�����[Ά�%CyU�3ȶ֏8�zl �n"�Z�$� &c��������fjnO�i��������cWђ����J���rݞ|��|�s�wV��ƿn���Y���~�������}p�~C��c���岉x-���d�Q��}�*�rm9i0
eϰ�ypm�HM�˔H�	�T�O��/NŽk86�M��_��k����_)u��Y%1�=��OG��_�k2�l7Yտ@C~�]C�e�V	_�:v�Ђ�K1�>W	
���г��:���θ�Gz��U�$M��~�e6�k
$'r0�����?��|�N\�B �{E�')����f�p�S�z�G/^�˃����e�A+!ir�}j��Æ�+v3����^o��v�٦���wZ��4cI&��i
?��y�����3�:;�����N9�j�j۲ ��N꛰*<Gd�{��Ӷ�|n5� �L�6���`U��(��*�����!ٍ#(S���9��++�R'��"6� 1�<�����P�z��ϝ�US�c$�m��}tHkX{�ɸ�?��K��l�ㅁ�����b�s�Z�m�A�m�v��0�n����p��������$$����9���w�s
8<<<��[o���J����P��ү���sF^%A�����F����q}��P0S�GԊr'��yh4e�Bb�鳫�f�9hDSW��b2����i��f#).�t;u��D�Y�J��0�hSs�!w��5y��)?=��0�VCB�i7aI}�<�XZ<S�%���<ׯ�Ȼ1+RRZQ���7�y:�7ͧ!�00h{9���O�Z�*�{XA�������"\�h�6aԮ��&WV���U(�1�!��\D�c���Y��S��Ne���n�q�W�J8ӷ�ej��.8h�ڋ��ί�du6�ARgK5G���#�./�r����3��V������gq�J��@_= .�8��>����|y�'L�g�Z<C#.S�&�?"}�3�+<�p䳚o���b{�1q��F D�����r���gΥ/��|9^�\G��}EL$����Bd'������p���">���)��� �º��y�ݾ�x�P��8�]I���ke���pڵs�#P�o�8l%a���R��I�'5�9�c;��x��������BӬ� d4��FI�s,�o�����a����J��*G_�/��iS�F���m]C p���z>�����og�:�:�|{S+ T�i�G��A)@N�Y3�-Y��i�M^���->�'��Q'�׷���'���P|?�?��t�A�G�0\K�&2�.@��U�#:�d~�{�zmVv^��Yd	įf�Y2w)1�@��v��JɬX0��h�yOhS��8N���S�	���u`S��2+�^~B���6ͽ3��Ck��`����{�A�<d����χ�z�eR� ��s�r9�k{�Ք٭���b�e�����g�H��i+:��5��z�S�T��6�J��U�6�I�A�r.g��ڳ���b��;��/\�@���%o��4����F��}^��w��z�R~W�[�]-����c�Q�i�?%'﷧�gEMp)E�lp{w������VZjN��~�L�O��i�5�ўiy+���C[*bw���̂��	���d�Q����iI����kP0�gWI^e�Lt6L�6]��Tb�=z�l�o��Ò�]V��] �� Q-���jY�%v:�HC��j<W*pt���W�p�D�`D�fx��7�	�, ���Yr�6�<�?/��!+`��/�&��i�{^��CF�'4i�dg����f��u�������)(�x�Qy)rA5�5�I�>��:�*��.�{���:2=wa0��W�W��ՋF{����#4#R��$W'���4r�������11R{ۛ���������1@�="�Al�0���U"ȩ�)ܧ1���>���z܀���P�+_|�B�9?�q���rg�'�d�V���(v��VDD%�T�6=�a'i]��rr�3�S�2q|�p����+��(�_���L��O���}]SO��X���~���}*��nV��h��+yAĦ���������NHH�CZ�A�c[2�x&��4q��(T��&����<%E��5��+S�0�&B�E`���n��+c-_���
)����I�;��M3�8^�e$#�$.r4D �IX��b\(ռ��̴��;�y~ޯ-�w�:�'�\��˅���hg�!c#���}�#g��V��H�� Rc�b�T�F��뀲�n��xIW��ˌ�ڐB�s����k�{�ZK��;.L���np;�@�S��.Y�z�N���̭SGx@@4�9�2��GȅCGD�b6wD4�v�xk֧B� ��u@��d�z]dl���Ep]��Gg���Hߣ��:Z����'b�~�N2��2�|F�z��L75-��#��|OCZ^?��E��K\cc>�T��Q�֡���� �Y�i���t� ����&�����b�""�l�o­mP���&���I&�@��l���qJW��ҥ]e����Jzp���>�y��Ȅf�`X�ȥ�k҃^�_�0`�_(ޱ��Y,����#yF��T�|�U*H熱��(�a,ǅ�OZ^��B�8B�^2�@��1`9b� P�f���"�8�6/9��4j��ދ^T�H��L�UG�6M���¶�2?S��$����L�@�>�G�#@M�g�9��Dd!�Z*��(NnɎG�@����������E&���%h罔�t}�/�����~#+���qZ����Y��� �� Xvz��n��)^z7���2��Lr�+ �i����⯠���C�FpU���"����L�����-Z�D:끭R���P�o
+S������Ƌ?��w�/\��])_aS_�S�A@uͨ?�xX���t�3X�ica_�w?C��C�<Y�!�����S�$��.̪�	�rv����l�/�%�T�;BE'���G��"!e{?��~D'���{�@'����}�e���_��G6��.��!}uJ�]��F֠� ]S�[p�ԇ�MI�y��V	����GiD-�͖c�o"��+9�K,d\�U�,��8 ��m���C]E�XC�3��*f���J��_"�Ҧ�(�e_p�b�٩;�.c��L����0��m�}+©E����T3S�8�>�!(+�M�vf�䙵m��H㗄l�0@�H��!v��+�+���M_�
���H:e��,V0��U�Y�ﮏ' �D� �{�؜���=�VDђ���l�c�|���b���/E����`��K����S>�|%� �{ ����6��}K��e��uQ.	�"	(�`8)=�
�ID�+�ed����,�����X(�ɴ�E?������@��T����N���5%�2Z�=l,�9����H��!@�q+*��!��Q��E��r�6�����g�<��H��5�þK�Z�f�>��TR��'���l��y�`�`�����u�����|J��~�ڷM�v�/�R���r�,�1{Cq5�$�7�(mf��MMi�H�Z�����F�R�����歱�/Z~�󧺀�����ц
7q�A�#":<�1�����f��ȣ+��nҷ����dL��a|*!��Vd��ٶ�b }���@a���D�]���*� M�P���� �0��+�����O��?��U��¸�DcK��;%�L)��dP{��<�Hݨ�Tm}��u9;5��F��is�x� ����aq�[�Th������p7F.6��,'�@^z�%J0"���j��1֦EU8
$��%�.44;�\����~$�j5��Y3_�iY�����? _�z�b���ɦ.�%��Ր�X�4Qm�B1zQ����֜� �VKA�H�Ì���x\��ӝ�bH��&����X���!�@uk!A)�5�x�����jmjf���ߟ�@T����!b�`��VJ���׷/�x��(���� Q���[Tv@������'8K��?�W�����b�������sV�ϳ"V�Al03>�r�fN�^��nu�zl:��iaj��:������)�!~�xV�s�Њ\�N�_��f���$,4A�`V*�U�W�`��n?g���T2��,"�,�(�S�¢!�)ۼP?�a�>���
�6|�G*�q����U�a�%M���� Ѣ������zh������xB�������r�WQ�����Qg��������i��r��ʂG^�x�ck�q:�O6��ƭy���B2�Ẻ�T㬮�ܹ����#総�\���W5z겴o�*�^w?� �JQ��o����j0r%I�#ߴ9�d��� �����z�}����8*�U�����ﬞ�Ұw�2G�y���r�/���A�|Z�W��׊
�QK$�,�֩~z�U]�
��y��x�,N[��>Е)����-Ҽ������e&�W����[���y�Fp[��~�:��S��naG,
gc���ܶ��q����a���O ���o��~=�T��Q��}ɨg��I�\Pi�`0��ϐGW::�[��ׅ�[����Ew
�CqL����	a'���Z���`��V��&�ZU��k�sl.�,�X|�%��g�=~e�s�8�(l{N*��Ţx��Rl�F]��|QFʮ�|:�5���.�j�;�lyy�v$�l8�v5���U��Z��|���%�.���zD{���/��x������X�ΐŭ��L�F� }�,]�]w��CA2xG�b��B�c��b.��8ԑ�$A���0���e��O��H�F�3K[��C *p ��y
�F1�!JM�ud�`|�ٱ��!A�@�m$P4/�Sx�4@�����d�����ӡ��:��ݡ�/���]��[3��'��DiA�����{��_Sg���/6%��wZq<��wx} ���B%���`���@E`r�?��=�I���_Ň������r/e`�U%�!���bq��r�iӏΊM��d"�e�����y��=-u�Y�:��H�񾅸Q�tf*�a}+5�xw�S�a�@�$�P�ע؁Jw�.+�8I�x�[��N�A�o�0(:�S)#_�K�@�>oq]SjK��p��s��wz�E����4c�f8���T�3�ePՐ4��l�g
�N1�R���\�?;�Y��އ�*��DBP���/1s63�E��٘͘��o9џc���M�P�g�����^�u�����2m��q4���#�sH�դ����,o0�Q����� ���,��K~���s=\n�.���>�p�o���t������c����^��.���V�)<���E`�/���
��>'�<Ľ>@ҩ;�$�p�@ρDJ'��k�8�y�籮W�����^���闁���?�L=�"3 MW�E��U��R�Kխ�d���Y�wi����;l��E�U��P��O@�=?-|Y\����� p�&��+ggf����*O�*Vn��.��ƙbsP�_�.Ep�s\�2ŭ\W���U~�W/-�^�?z�l)����h����;�N9#���y0C�1�6�x(�i�ŀ>�:��
}��}(Y����C�ƺ�E]��t�d�C a5�|��"n��r��`V��'.W�%\5V�]܂v����-nfD�{��PB��4z�/m��O�u����Afm��V�ʁB���#`Wa։� ���61�?��۹�h!.k�g���$-����U%�I��jI<�[r�1!�8k���:���$�]��N#�����0�M�������Qfs%r,��1���Z�����Ϸ����(v�E��������w��K�����>:nN�����ұ'��, 9�g��w� uÙP�O�7����#*�W}]��$r`T]>��h��&�����MB�Y����<�<�|Z;�9����+��.�?\���?��ϊ.q3�4Q��l}���-miv�:	�T�W��S|sJ��0���Q]�}�\W
���!�Z�~�=��z�F�ȭJ�͒�׸d�M:��K�IOaBQF���Q>K�����uQQ9C�h#4�vꎧ��TU°<{��R��}1��m��o2���J䝬I�*������}b��	W3�EP��)\q8^�^�h��ê����m�)��+�����.'ؔ��מ�۷��O������Y�����[��,f�!B�O�י)*��\���� �o	���+/�8jAi�[�����W�}���f�'� >"��rk��܄�X�OHX���	�L����C�ŉ���cߍ`&��V���]��Lը&j�����5hN���\>�3|(�%)Z1�^��k���	�o{vDo��}1��V>�/�A�����8H�fg���=O�vl||6�D9*z�U��+,��mt��2�3������s����׻K�ϻ�	{[�`��q���c�Ur�PQ�~�������އ���z�ƤZ,T���R�d�~s>X%N��*0��P�%2��3��h��|x����z�I�u�x=��0��Z���9}M*v��͓��;���;w(}�����]�P_�ģ��G�FZ`٨����v����
}��7��F�B�Ȗ�]���(���횜Rq�-�3�������N%��~�s��J'DPUy����pAKK�]�Wb-�IVqhN�����z�zX�_Bg�H:0���Y��d*����[�?�@����І�kP��$��V����a��y�О s�ǂ�ȴ�	�rEi [���'��NgA57v�L�Z���R��
������|3���fre��O�kvH��ZS�i�+0����WWM�(ĵIh��7s��1�YXt��q��X��uk���̮9�����m���_����.B�X�BN��;T'g�Z���~,��&6#=��r�.�7���26N�/3Ṱ�l^������R�(D�"y�<L\��<�����I��q�tdH
�����T��2��JUf�Z.�)a9��V��g����S������:���k'i�8il'�m5���v�$��c۶�ض���מs����_��{�9�k5��)zDw��ȗ��hv�%���q4��,ڢ&�����1Lw���!��U ��8l"�+C��)��h,�F*��x�O�T졽Tк޲�:p����^ �b3jt�O)=w��z9�H�)F�����K�(�(�6�
��K(J���-�vA���ņīb�e.�6<eH�8���)�$�,#�"Q�YR�C����a5J]P�ee��"uV�d�� ��.�����d.&θ�o�f��/]|�]�}��B9a�~���z���0���H ��~z����컠4�*���2p�(�=�#u �ec�dhVn�a�S�UG��b�I(/Z�)����_�VK�6�}n)�|��N��gf�����MFw�M�W�,���[�´_��So�]��]������nQ���ܛ	�kZ��{M�z��|����L���Ւۅ�N�5�_�ZpwW���I�X���E%=o�i���S|���$����0���֗E���%G?r������S��K��Љ�Oz=`6� h*�jY���Q��Ҁ4�k�?xf�Nd���m��r)n�v�k\��3ro�����ɖ�d��Bg跅����v[��eE`��
C:�%[=�܌Fޟ�4n���
^\mg�����0�~��5
TP���Ke �n�B�1�%u9YH���v���@��x�y��������T	���h�j=��m�1�=�@�ρU�}��]]z����_Z�� 8~^s�=xF�l�C$����S����� l���b�R3|+� �m1y���3~�<���^�XBn!� B���> W��kפQ�H�]�?)�ҷ&C~o\Vgtege��k���N2�[E���6�kնq��ֽ���>�i�G��'�����zX���<u���e�x|/����s���Iz���;Ƶ��3��JWD�u��R��!�F(�����t7g�Z����~J���企&�����^�ƊM�zg�qe�"�`�h`����l
]�{@����%�qDޣ�w�#�)�Ѿ���cdB��vB�@;�3�s�^-��n��ˆ�D�,�P��ѝH~�u���З��z=�2lX5�	V�k4���l�e�!/.�����۩�I��g�'ż��BuF����m�x��Sm**8��4J�	Ni�N:�CE���!^��(CW=�2�����@����~�,0�m�!�Su�]+8������2m��Gz��[,?ʱX�D�2`ky+�Z9�9/~�Xh�r���%I�m�Y��#i�̏�>��u�'Xy?Z=����j���y_�����W�J�%���/+�H[XSc�"@`S�H���(2��O�X���_õ	L;��*�G�M``��MS�ۙ��/��V����b�c/B��6��O�"!�g�����2�^.ӡš/�ʁlB԰�"�&2S�����߻}�l�&�HL������,�3[�Y��
0�z���pY&i9�@{����i�"(��L�:%"|W�sM�5D&%���d��J�L���0xR�4��ɗ�������W�Ǉf�h$S�"o0���%ǁo��Ƌ9^��%�7o��cq?^4��%���%=��y;�5�ek{���7����a��5}�5���H~���U9�'?u�E}�6U@��G/`��"L��I��'�N�7�%r,-@2Su�C���p� -�$�L%*��O$
6q�Q����V#��v6N	�|ř�#9���@�ݮ`d*�v��]��@���g��'���8��0Co�]�R���k�9sw��SHK�u,��s/h?`!��ɢ�rZ�[�b���K����]ӂ�(o���L�/Ȱ�x���r�Ѿo'��/�%��5F��x���:�fg�D:o+��A�����X �(��HD������!�?FZ�,�b���U�� έ�1Us䙪��Q�$P�4&ڻ�~E��ws\�������TOR��Z���T�^객���ǁK5��b�>��/�I�PCd
o�`t{�c�P���<ǆ��8���}�����W��a\`���+v�n̏���#>?��(���zڐy��2���i�.�Z8��\*CDz�(�)�3fˀ9�vǮ�HWd��)x�r�{~J���ߺh#�F~��>^�o��V�[0OR�n����/A6��u�@��ߝ���'�Z��(."��`5�Oכc���Ĭq
ađv_��.6�W)����X����P86L�����cX��������'i�8�Q�:uX?0 ��ͱ' jn�����0�M����y��n\]]��0�����o�a�����Ss0����,�V��oz^WOۊ%<C�}�U:L����́���ufY�;R�qG�tm���T'�����ymS.��10,�t�>�D��	�:	�:M25D�9{dǄ��E�	����c�e�T��L�hHݞ3֜/��&�38	��iLN���f�̂|n�G�n��KR֨�)�`��bp_�d�G�23�b9	��{�m�}�h�&����y�н��Q�}\����΃[�ׄ�ر�|>[{p�೮t�׺S��Z�J9E��$X���ds�4�����1t�*bQ9�;Z������G����	d�<�`r�}v�{�d�2�,��I�&ED��9Nu3��	��QxS��~�lG֮��ʐS �t���h��lBNA�?�Dp+a��*�C��.���O|.��A��?.
��6�$���@v@��t����NP��M��5���n��a�b��m�V�;��;���WQ����;�;�]y�ȰMy�չG��_u��]�ŗ��U]W��4(��-3מ�ҕA)�1�sT��̨�J���q�h�Q���e�#� �n�so'���Y}�������l�[���!��.D����zT��{ښ'>��[�:\�9I�}��'����JR���%n�WB+�y[1������.^,^��d���x��f�)�%�~���)���Gn��g�$���a�f��Es�e#��L4�W���PM��N�3��>�'C�ܱ� ꆉ�+0�m0@/'���$~%���m�]���ݚ���T��8�$/����8���EH��M�T~���Z�HC�,�wN�D??�����f�w�JTN�MtM��,"m���\��!��-�2�׫A���I9o��D���L�LbD$z��B:.�x4~�D��f�U��t-7��y{�(�N������MC$��ۿg���C�5Y��4�)f��]n�>����/���9;+���ʴ����h�� 88�8K�q�m��f����+��	d��΀�z$HT5/��^��RP\�2�� �;���5*'��?�P�[��A�|(Q/K� ~�2p�4���;���:���μSO�$�������ɝ��6���Q���$�	¢5e	e����e�V��!g<����I�@��I���q�=A�ڶx�C�̏�������6�펇��8ӻl�-渓9�]�Ъ�-K�+��E�`�D�"�x�Kp"(p����/O��\l�����HD���>U�~�M�2�'���ȩ��(��Rk���/Y��Ϩ�V���(d���ϑP����>X-���N��}��g��>� !�������}jM��f�~����1�X�J������z�n{:���V��$=f���櫞X6K5��M�j_��׎qS'����ڢ���a�L�(O�?#��bJ�k���z8V�ty�T��6ZCok�̍�Q:������2�;�������GS����ʠ�]`�|��}e��ǀO0��qUKg4PB�Y�E����2v@	D�F�-U܅3��K��K���@-��P%�QP�1J��$�:L�qc��'��-=���t����cx�^���b���
�}�8&�؜j��ov�e������>{�$BmTl�Fo����6{���;�-u�X�,��Z��*o.��\FO?�>X�(w�~_ls�P�2:|�.��a���7�Q9����(J�[�GR��m�����!�s0�ۺ��8r���@9G?�O��^Щ@9��|0��Գ��b����ֿ)+�XJ٠T+�|��v�'�6{�?
���G��*�*�A_�h�c5��C�N�NkR�H�f;P�uR�Jk,�V���:���s�$lx?�jV�zu^�И�7�v01�a�$Z4��`��h��:n�Ԟ��[�<߹��h�덇KW���g��v�f�����tyv���݂����5�&���h���UH7ɳ��.�B�~β��'��7Dʕ�"8?rZ$���0�~�%r(����^v�e�bg�N�h�ˣT2緼�*�eB��� ��'��Ֆ6��2t��V ��[��b`23�����������R���v��rX�h�k�R�,a����3ʸ��3�^O!��aYzQeOP�>�J�f3W����������u���qtUҪs�3>m֨H�@>9�'	u26�����\��)D}�@>v��<������!�}G�bW�*@m�Qpŕ,QL\���S�����N�t�¼�k��z������~/���T<	��N��-5FU��=E��?�Շ�/G�h�|>�/S	�Į��Ϩ�����w�(����CC8c>���P��/��da6
�{��`���{{����6Z<�/D�Y�z~[?�~��g�cc����L��@$ྭ�W�u%���gzm�D����'��No�?\p;�����P����.aj�����,�4#�&�G2b[�\�����o�됀��5��~����z.��Y�6�����{�C1ܢY�m�@6�^%�ł��Y��7'���RÙ��(B�n�v�n��d�]��S3~�s��+��ZJ�`�z22m�>gZmM�Ԩ��^�cհ�j��'�s,�G4�i��#���#�|�E���Ԅv�Ҥ�w5~�v��򛲌�~�Dba�RD�f��do�\Tj�k�6��Y�o+��_���9�+��p'��~�s�l�-h��<`'GFJ��N�2���o��!b�����7Fz�9�� ,gK��ѩP�@�`�/x���m}�$4;�<��t9��/iR�*|J���<����6��������O��������H�I�z,���a�qX����k��9�0k<���\�ܵ��{G�?�����邥�(8�y�C�8�8�8��!ʙ�/��+��&����Ɂ�t�F��y�9�������αwg�th�NΠZ!xc�����v&S ŝ� )���m�5s7��o!2�N�8��s̼H�ٰ��u�.��	��x�ŸI��W6G��R�86UOw�S\���tJ)&�qbY7ʔ�e�ʕ�L4#��&w
n����;^_˺޸[o�=��YD�N�*�%5y��2&ϫ�_��,wI*��w�����S�d4�}e�̠Wh�V�ļ̘/j�*r��(ӳT�<�$���%�]��g#adr�qQ@|�!iB-DЇ�r:_�4�Ap�Je����@�����R��4�zX�1j��8�0��l���,��ǧ,��B?5�V���ƃ��xӏ�7��C�y5=}������ ��՝�!���.1rSҡ���N��߉ƛ������t��Y�K!���"<]k���}�`1��q����j�Q��b�?�vg;:^
��qƐ��4v��7вJ:��^E�p0�>��P�H�/nQ�.g�"&e��Ts/gZ�d�npܐ7�j��xGȱ�e����W�f�����G���<Ӕ�9O�N��9��m7�1�)o�n�$�Wo(��n�Y!Z����v�e�JahX�&C��3)��`j���h�W���Ȉ�]V��B���3V�'�Z`������SujnI�di4�w'���V��5�Bf�"؎��T���{Aa[f	:�ʕD�j5΋�߁A��́��=�"����t1	9�������b�� )�@���<��j�B;�-�@��=��2�?����v?5�(�~&��Ծܟ�Ġ�<�m��6�W�<>6k�r�A@@ �v_��	���& x�}�3��\]\�.�q�S�����u��d!������x1�D��į��͍���~h��#��f�����%��J��dNh��	���弫�x(�Tr+o�p�8�eC��!(�z�1�9��?��O�S�P����҇�����8��]6c�'�ˤ��_�Gv��}a/r�.(�l������X���2�C|��A�	�����\p*C$	Zq:��-�5I\B��y
ߋ�����}��Mߘ�5�ܽ^�G�ə��4,��,����V��4Fת�\�*�5�4��6
��'�À�@A�>V\g�?��b4�_	avP�hq罕���W-ё��� ��� Eh���'�:aaa�l�n�����_0���|ԛ�ApP����G�3��I��,�t��':�.7Q(���_�Ҿ��W�vhb��2tE0趫�x/�a�sWg�ȵ.����c��Hmn�㹹���-����t��zE�ㄓ�}x��;��x�{���x2��Bm�^e�@V�#'k[$裸�&�OHO�;7ֆ����Mx,Wb�|K��KZ&(��l�S��G�޷�Q3 ����1�M�8�J"z^�M��D4�vݏ= �{�=�	��n����,�EM+q�����)o�������?�oPn�p8+�_���0�WU���~�Vv�|A[��ωV}}W�ܩϨ�MX��`�l�BI�H���JTf�����q�����=���n�wp^�꘱��hԺg�}�&�ў�N,hGء��P�R*[FՏ�X�~�a"
���3ۯ#�/v����T�<#|�Ww����jaEqa?�%�4�����!�D_�4��(�������;���,I��$�"�����N�kNr����@3�����uu�x��� �q�~Q��=����}����>&�>`����34ED�̟�y���X�64����5�YW�(Ik���fњ	5["b��kƜ�U�Tq{�����Z�>6�/_� �ݢ����-�[f�	@�Ix��� ����ə�5�����S�:�)�T����r�����K�K���B���Ɗn�0��SyP���Z�
w!j�N�lԴZg��7C�OTI4���iž= σTd)�3Y�5�\�A>R-v��7�:��x�u���
���w�uG�أ\rY����
�8�n%�e���Ff�ztI��J=��ڎ���ǲ�E�7�
y�-؉�&>�~��������ٕz �F��o�˓���&���o�oʤ��:`ŀ�)a���զo���]�4~��;^��U��n���g�mj�ՇY��;3Ҷ��.W-�]M��0b`�7����b������ac��
��vZ|�A���}�TR��� ��|�UF$p㭝��~C��{�ޗ�ݬľ���r��eY$��J����y�g���ع���O���dҐvL�	'����ӄ���7A�����$N�:�Jj��=,r[ٺ�~C(��&�6��6��ɲiJ�+c�O�Fc����	(x���ȱ2�5����&DR#Ias}ٻ5U]B�O���<N?>�O��qd�y��l�Vh��v�ܡHQ��a�wg�Ϝq���(�r��*)���K����Q&J��D���WV�6L�)Q'����� �D�l�Pee"���c�-��'���7�1o%���I[�E����ze���m�>Y �����9=��AKD��&�����~�@�c����<�4������U<|��qǟ������nA�l���||�M@��h�w�����/��;?f�e�n�!�vw�S搬"���K�m��������[�Ox�w�õ>�(_s����z 7��F ��:�o����Q7\<w��+��6�5NF0?� p�Dq�-C�q�np��5$6�־�����&����T�6VU�D��'I�S4�A��5���y����TpN?Ȣ�x���^�R��Q�$}���u�p<�X�L�{�o_i�b��~��.��w��$¬��6&L��UO^��r���`��o��|�C�:�l[u�������JRy�hZEl%
qE8����ov(U�$�[��S��B~�|��׭%]dd7��Q;�Q�M�߅PPu���̗"J��b�C�K��f��ah���l�Sf�Ha�rn��_�V^��dW�s�%��R D���[X�S��AY�}��?�T������sd0��������(��|O{h!~}��@h^�M '�/Eu���� �����D��SL������y��gCT���3`a��_ц�(�)8��R�~�\tu����m���QV
P��d��N��x�@AY@�:��3xOh���,)�yڶ���Ք�d"y$�7c�爾�邱�\�����6���2oI+���AE�&��LZG�В \-��/͗ N3��C(n�S�nZO�Sg�O���H@b��7	���� �������^3Bm���^*�g-��<���3+����ղU��������~��,���^�ܗF�P��8�K���4�xG�K8E;�a��'P��O^�R���'�	��x����K@:\zػ�m�S׏�\�����Q��./�t6���س�����zߛ���]�KB���ϋd��k�:����y��[6߿K@cu�Y��$����+q���F�q:����^<��x�-D����C��\?��~�j��F^��zrE���Lo�hs9��Ē�iZ'��̠ۮ�'n�:�X�⮮��`��apO7���]��4�`�-��Y���k|)�'j4��]]DK"苗u�ϕIy��yhk\���CqA<R��s@/,$"n4E/���ȇ������)�_5�"��-��h���s�!1�:%�x+(n2C��=��L�f�rO��̝7�W�9�=6������>r
��.��њ�+T|R$tv6�����f�<�������A�ja�2�$��ق��q�܅/'	�lhb����|��{E�{:�B~�i�Ĩ�K�o�t���z��
2��C����g�&�#H�p}�V� ���4�Nl��Z��ǫݬN�I���l�f�?�/|���n��ߗ�g�x���t�8��Z��I�5�=�h��M�#�C�j <���B	�`~Tb���s��Z��_���yRhv��o��%y����e e��AԶ	ۛ�[�6�3�<Mv��r�zj�� 	�M��!�"M�@���H��8�ﺎtq�����҅mP(��[�]¼<�6#��5�H���+i�ݰ�A�?�=��i�Q�h�غ<�A]��B���C\%J����/M�)�Ny�G��F�XF<�pY$c����JBPC
�%e�	RH�,qTY�DbG	"��^x��x�7c������e�Key��&�>�"�V/m��g�|�ݷˈ�a[ss�wD�`�d��+R!f�un�VS��|?Jj�H˞w�m�U��Cާ���GW�}G7�?4�U�����Gl�J��M'Ow�%���M�p�ѝ��y�����c.�xs��o���,?�?ӈ�Dzh�m�!�$��n�0�;]���3|�I<7��/1��>8=eP��^���X�b��l�M�4�M�O�Ӑ���J8l;|��2�?��V?p��	*T�34���>W��>cH'hع�t�]�U���v�6������5����U;y�|�H�Z��.��;��{�{}��ئ��m"�h�$Mٖͼ�U(Ek���&ڱ��Ea�z�B%�L��TJ�Bye#Zq�� e1&���id�5`�A�E0��YD�t䶚�wQ@\�e?��v���s5���]/�%'_����E��N�]��<j�Ǎ�6##@�E�������r���s�k��pS��������W6<���U��;{×���&<�_��Ȝ�JEr�^ٔV��}!%uu�
w1������ U^�|��PIe8X��$�������/1�R�I���9��d�Vt�VG�r���<�K?��\&�*��-l��0#�*��n�7���(�d鐠��c�4�ᕡ=+�S.��q<�o'��}̩�2ϴ��dUH�>+��ӽ�H�'<u�*�YVNfzm�zs���ujW��</�da��B�d"b�H��>͡��d�/�l����ަ��r�BqOD����9�k����c	��ߕeC�f�k6eK�x�m��5�0�h)�NK5�ٳ��ϫ`崷�kSyA�	(+j���b��kk�?'��z�1�M!:/	���+u^�>*:<�n^t�|?��?`h�4�Y�yy��B�>P弅��0CD�5iv2Y�8�#���p�@Q��Ny���vT:�Z��i�EJy��[I*e����C�9t%���p ������7��{+B�U�]����һ�K�s'����o~�I'W�J+���X9��gt�d��T��̅�4f�T>���K�U�V���cB��`���ۗB"�~���_�5+�'�6��be�V|YF�Wł`�ʟ�؟A8���j��G��m�x�9SeB�V:�$���*��V�B��NJ����-�L͜;�U�3t��W���FFiС�ެM�j��S����=�����@?ZaݚL2峬B��di��+	Ww��6͟[>1o���N	۾�fk�G��c�iܶ:��>v�Ý�G0�O�=�!��O��1����%��궷F��E��?|i���|��!��n솙�  �H^\d�D b+���A!'BCS��L����{��5�T�T�'����q�'��I�
s2ko�$zk��#�L�kA��x����r��_9
�&|��]j|��?,ؘ̒g^�Ыɳh�GfG�5~K^�l�yG@LG1wL��ZX���Ѝ���35�,Nj�Kq*����j��=?4_"�#���'��H�b�?Ђe-X��R�f�U��P���d��kG�!����&Q[���t9�%j�J=�3��6Z���������^�������3�5Do��jΠE���+�@�P7����VQM�dX�m��ry�����h"�4�X�Du�e
��f��`�����R�q�<Z�������b�.b$s����N�͚_����n̶ᩱ�G�4y_N�f��
�0Η��)�f����iX�2��:~�C���!:��'��`_ϟ��Ĩ�R�L���������RaD��9Y?u�͉<^��Wc��:D`xT�yJbR�讀���-"fr��&a�b~���I��_P�N΁���"�]�c"V��g�-���T�d�.4�(��SEA��|_0^�Y�S��B 䮞U��u[��kC���?莤�u�Qs�ȂV8��ja���ܺ��F{��F�h�tO[	h,�Rn0r��!O��W8dAR*�c��iJMs��8��ǎ=�UD�l�Xd��(qΏs�B�[���.����L*�%���p)������T}�n`�{tL��,��B��p���Uz�\�,S@��B[5A�ZI���(g�b�fYQ����թ��)���8�k� ����������$P�4|r�V��$P=:(ʫ��b3�����wTg�"��|��bv�͵k��=�����BX˿���������du��_��a?������$=��r���ZZ�"������쀔CV�J7oQ�W'��O��$/�H~�[��ĔE~��^��W!�RB@r�G<�ę)�� B�'f���p�r2��d{�p�Bf���H��J��^|mW��J��t��C�$)��G�낅���5zM��ZZ�A����δw�f+�>X�J�r"N�tTx`���մ.(,33����Es+�Ӌ1E�yŖ	��\̧�t�n�`oF}e��I>�|FA�^�t���rc��1o)�j�?~�Kvxj�fzj�<?�|�Ŝ�#��dPkj��b�VAq�B�"�ʔ��Y�S6d.A��wH�Vbt��S�5�B8���]3�����$,5�
!�4�ݠ��O�bԐ�;�;/;{��a��������<�
��{(��*<>�%��$R���xT�O"LOo��l���|���o�^��/��¿��."8V0D�DYi��^�g=���������/p��tLMCa�`s$�0p,D`�?"=�%Rf�]���$Zes�����GnYX�V_�/�z	PX��+�5�0E=��q�HXπ/K���)��آm+�$��h��Rа�x��V�jm��&0H��w�dA���,g����5�'gj-�ǹ�h.���A�팶��������$�)�L�ch乤�L��-�j4E����5ʞ�^9?���<���&+�R�;��&Z�̹�
��.[D�(���h�'+�{���h�C;�)�3(q~Wȋr�HDz��?f[��:�Ǽה_�$�v.�YwF�3T8,��?~el��>T\0�4�w#8]I��wv��-C�e���y}\��oW1�q9�f�`���7�x��4���v䫮�y.��n��-��b�*ր"m������}oy�̋��YX�tQ���*�_�  �#��ȕD$���-��{�|��m��L���4�N����<,]�٠7�3��Yf�ķ������J���1[��@�>Ў�'{��e^��7��n�����x�O�x酶�	����N
bJ�V�^y��4	�n��j35_�fno ��)`_,�v,v�)������b���j�+;��<��ҐJ�% 
W+qtPT�-r>^�Sr�+W�Y7�X�,q����\Q���L���H!]���硓���1�)�I�c�V6D�I'�u�,L��{~I��d�Ţ\��:	p�������ԅ����u�b��.�v5Hȿ�����{�����n��O��t�G�����,�al&�ދ��o����V� ��	ю�HR�"�d�����~)�]F;�������D�B����ζ�O&�S�B�Ci�BN��R�0+(���7���R�=�t�����=��pB��Fc4�po�:PcX��s�M��kp��ou�ȳƪ%�W|5m�FՀ��h��b���Ү]y5�!�Z��Ty`HX�U�2D�䔯\�,�=�=�^;��A�fyY����r�r�������K��B��%[91��¨�x�@���欠FY˰�f+g�bR��TU����~��
���Ϥ��̢,ҥNvYQQԶg��*#���1�[�oN"t��j�Dk	�h|t��SB��.qN���!�E�c��I�,;�c�JcF��0��_�nz'�?k�%h�����7�Η���~cjn~������zĮ:ls�������]a�k|q!)6.)7��xؘ����(���*�ӈ�-T�&�r�V�7$X��I8�F��9���t���Vc�������; ��A'����Nj�p�^߉�㰲�	$ry�lrn��yCi�^�&�=3c�3�)]?bP�Y�br�;<��zh��ў&� �&���?�*d���࠱�-�X8����{ۙ)�@RP19��I%=��Sl2����Z�栧ƫTc���d��o"��sQgn"�*�S��}T�;AV/*�-wVLk��>�BD���i��ͳxnS�z��b����S��<3�L�;�6���S.)�A%e������G��g�I<�\Ց�*�{��b��v�s����e�7S{z<ߚ�۵\G�z���]9z�t�C����ϓw��%m/�޿����Q��5��Ԕ #3�9EF�����I�>���խ����а���Fe�%��<.��<H
�D��l�Y�c~j�C�
>(WE=��&`j"��l������� #�~_��$��_S&����� 5IN] ql3�\
0�5��� j]��<��
ޘ�J�Ŭ��B�{s��9�f)QY����~[rd�w�~
9C�3�n���_���NQ����09C�:;:[\R������U%��+�Tj�b���#��U����XO֐G0�~Ӊ�ϡ�.�����_�p��\�WM,�DZ_]�KLCV�/�_���kd���dO��3��y�ҖJ'�~�jY�+���K�;�_�e�G����yE;wr�2/��k���yO���J��v������	���u�������{�f����É<###�G�0����:�;ʱ���+�l��>�'e*SK�� �cu����HC߷���rK򹹤,.6xs��.�M�a3Ќ`uw	9%j��]�!k|-W�l�t[�U1�pv K��.)a v�ǎ�+e����v9�A�-�&������XRK+ �[%�b�4�� �2��Jn�� �4� {�|����� z?�bU�]]�٦�믔��k`U��HX0���V��6����P���#�<�N.���xsT�	j@��z����<���+����vT�ܙ��V�WY�߭�﹧�e����7�}-X@:>��Vd�h��d�K�F���,Y�h"��jH;�4�FW*�&�T>��F|I�\qЦ &�/~�ŗ�����}/$N�}���^Ŋ	��jR�?�aH���|w��bfj�M����~�,7$���Κ�g����oq�_HN�����:�E���,��DP�߿���L����}u��!��6r����s��żZ%�*T�,h��!�]�2f�
"%��N&�-͞��Qr�����K�UK�=Q��v�7���S���g֛nC8qy]�Be�=���Q�ΦA�0P�T�`�[jZZ^�W�ғjBܺ���g��f�l��X=~m1ϰ�T�s|�P��H���e">��ģ	��Jj���3�{�3����7ie���:��)�?_�WyX����g�v!��R
�)$�p6��)o��'.�����Щ��_y-g�2���/|
(]�D2�șI9����]�{=�F�m�䟔���CUQY���}���n�ο��ѻ	����]������#{;���.���_�&�v��1)_D������I[$,�Ԅ��Y�k����d?lx~�x=�W����X��'{B����!�h�}�a�Р�)S�!4��ēۨ���SRhI�h�wPj��F����l�㞤a��>4�̺l9�`���V�6E �?|#�A�RO�=���)�,Դ-��S�ȸD��S�A�s+����h�A�7˅r�`���!4[�,A�@�m�iX���`H=TE�3��s#��������U��֘1�any_��/����'�tɖ��X��?�e~wC�7�V����
���G+V�g�+hi@&�6�&J\��F/떊�u��! p�^B.�4y#�������G�=����z���O���������"W�1(�D���3[�ҁ ǃ��g�ι'e�P\��At��J��W�$�Mi�\�:H�`gkaԵi���������������(J�G����ԇ�W�ī�s����,?8?����p��Xlub�i������8�ل����BJ'�����g�)�������MR'�@/�TV�\:��>N(�x�e��h�L�*�m�O�+AH�j�ׯ�����~#�̦:�s�JHD2�Vj��d�e��I�"wqf~��t�����k���$���&$��h|�%Ґye��B���X�diO��B�MEO�Z��-
����֮�#v�oN�TX����,��$I}1�}���������Z�M�P1���%+	�@n!�Ó�>/gMWi�W��f�00z�O~Y�40N�V#���FTqr,�:\wxl��� ��Iˁ�>S�Z��	XLٴȾ/�z��1������_tk�\*
�dc�4�\ ��F?G�l��.�=��?� ���%��3=�x_/I�\�0 s�b����+���n)��ĭy��ױ�%%uOW2�47K�A�_�@��X����F�9+��+�y��O����p�����7�9�':���,���	W����e�C�a&���}�!�a��#\�_��Do[��8vɺ�,0
X���ݯ��sѳɌ/��0��r�+���Ta�j4e�}X�u�y�pS��e�d��"ϗ�V=;G��K��:ĎW�4g��h�J��!ؠ��,�C�@���u�/bk�J�_�?ƀI�A+��	���԰8��7���}Z�ywrv��qRѴ��2%���3y�wc������ׂ�
��L�鿗��8.--�����Z����^}0��dBWH|��L�BZ8k YM��a���c�D\&>!Y��"r��V*ۛa�T�.]B�	���%�z�����"�7*�� �����B�����||�q�׷�j^L)�%�����/$�Qt����_���!�M��W�ae�T���ȳ1XG�Y��ie��@z�>�#���E4y��E,�p�.qa��}2�P\�/m�6Kf������(V���M6#�W�o>n$��l>d��K��_lj�K�0A�]����V}QQ^)��b�<]c`\kם�m;�m�jl;i�ƶm�nl'���vc�k���w~͜5��k���s@U�B:�kVd��`���`�(���F�{�*G�߲������V�n��*+T����.4�H�.=�3gAX1�Q�����W~7ZB��f,�K9+���^�R�Tj]�}��I�1����|�I����	�&�P�WP�-�����a��M���J��;�_�ȕt�K�a0��V�H�drMwdi���e��5_x���?^}YX^�l4����M������	P}}�H�Z���7k��ks\Π��
y>�>��,J�eՒzB\W�%>��z�h�܆����q(숬i�[�Q�edA׹2�i��}�Ҕv�8f&MQ���u�s�ۿ��>��%�R��;t#Vv�Kp��CY�d�G��{{�c����K�,��m~����p�#Ij��5��l�EB�����G�if�����s�!�ര��#6� ��+�v����K���j�o�-���4�o���C���J�k�4��[�Ʒ��N�}���h�o_����[���e�7H^�:QgR���9�Q.��_����%�y����%d��v���/Nzg ���PA�6��>�Ofr�fdd���A��^�HL���� S4��'�k^R����%h�ަ�r�^��
���Q*'Zc�쮡WE[ ��4�m4A�Bʸ9�����R�Z~��?��:�W�ʩ���Qi�M���jS��ƁT+9��{��i��N��Nwe:�ɚ7ok>~��7�-_���|Q�OUø�놫�yG�-ٺp< ߯7�pU���r�Q6����;|8k-a�Z��������.��<'��|Bj�����I�F�j�Z#?7q�T ���돲�UhyA�V�SԢJ5P�fB!�C?���i���q����5'�?���ü��K�2�\���裮�;�-�b���mHLW��싀�qe�m2떓�g{�"�cyC��@��o�6��������ܵ.��J8�ۦ����G5��@}�	�J�.=_[������C�cO��O&� Y�3i��ei�of�S��h��b�q7
�X�
;%h"P�����5ތ{g�"]]| �
� yiw#, ͅV������	(�:DC��4��w��,C�]��E���������|��\�)$�6(,��#O��P]�QT�pT*�1̀�)��"	Bh�� -ݝB�Mo"�JQ���!���r�J�jX�%�X`�,�K�:?FS�
�"&D���
;��;����ؐGS��`�P�l�%��R�L�V�JI*-v����ǆ8�Z�h�ͬ��D�j�:�T5�5��hiS�b�(@�t�a�*�Z3�����N=E�2��Z��\��M�C���+/����j��n;L5�Xb�M�"�,��!J��S0y(�^7�tHo��=��+��U���1b)�_^�X���e���w�f�Y���襌�!�ͳ<N�\���6E�&���I���X�l���>U����+�"S"����vc�3ENK�F��� q�Qr�Z%Oi������Ie�ҁw�.��d�l������[T��(.��`������N0��ޖ�7k��mU�-��޼��̝Jy�<�r��'�<���S���25��+���P�''��t�tg؃��.]�ް��*j�G�.9%9�D�nNV6Y�X���F�RRDyj}���o���ݭ�Q� �C�Z�#s0u�
i�C"1�Ԝ)�č��u!�Ƒ���y`�#J'I!߾�W���gR���7���U'XMJw�ms��H,�����a(�I��Ԗ��"l�
�9�l�(ʆh���J�yBҚS���N~�'Ө��E�3���p�8�蹰�W�@o�C�T��v�3�F�G�Ss������pyճs�.]5l���%e�ҹt9�sM	w	6���qE2K�vt�-�j%�{�<�E!�6+�A�[
����N�S;��ʾ��Ov���V���o� S]V�[�tn��H !�,b�(��F#�
�+�3@��?���%�L�<�"����T�n����z+r	pN� ��R�i�|������z���D;a�(b��b�K9k�����÷Z��D�$����T�����6 '8��(-T\G��^��V�UP[1[���AO%`6���
۵�c�b�*��MT�ke����ƨ?�i�jt���g�L��d�j6;�k�l�V���[�q/z��!�7ȯR.�Vճ�&''�zX[å��z�*	���j-0�Z֣�h�RƖ�L���0��B��M��*u��]���(g�N����$��f�1���fk��4� *�}j9[^pgp_Ǐ���D��*/]n���']<87ǩ�G�kN�h->aG�T.P������j�a��I�M�AC���<x8�ΉRW�����9����X4С���N#�:�w���ʠCFỖ���_��s.��x���> �4҄|#Ukj
F�-0������E2��|���Pc4(�n���גJHH��~��9��~�/�<Pd<��}�pa��� �ǣ��Y�`�r�B����T3�KJ�d�C�Gc�2��B8�Ib�1/=l�������l��h��AW�$���Ņ0�헂UU�����V-8	�+����E@e��^YW㦤����2�@˼��P5��U8J@�y��������	R �c�rx6�!��
����A�>����?T4�Ve�.N��O�<_�=q:���BS]��A8���Q9?͟D$(���Z���sӮ���~�8M�kw|�oC�[�C�"����Y�|VEה������I/5���� ºq��v9_���lyJ�^�tw��W�������jQ�>=�����D�-��XB=I~S	F3zkJ����!0~���J��OKj;���gcfv#^�O�|)�_�t���/ F��C��s6;/�9�1ڒ���ynyE8zu�};�q4�^�j%:��v^R��R�DJ$#
k�b�h����m�3n�Q��w5�)D���A�b�½t��zI��5�Ȋ���S��g' �L��a{6|蕂;|~����H�7"k#�I� HA[-����:����p\[Ť��`��R���{����Pg�	����2��(���/͠���j,�epٶ�tfk�3i���י�sTiy��0�p=^��<T�لb4�ő]�T:e��a�TZP����b���)X g�)�qջ	1C1w��>��œ�i~T'�JDv����w��:��ʠ�$g��ή>r����-^���i�v����h�p���ڧJi���2��6qw�:��$�k~.85�B��?�`S��oc�'�h���q��{��O�.:��3 a&�ؚT��DPc<B�Yz���z��fw������|;�m���veG�^ �~��sB�t�a}�C[�����˥���w�%�mAǓ)�Uxr�Fq?�*M/�WJ�MS~qj�U 75ɕ9>��q�Z^Sk*C�P~�g��cmo�-�]��%� ����{?S����J�߄�V]KHM����h�^�����_�/s��J���g2�]�`w����iE�r�ړ�7ĖIqm��+%������Ux���t�����7��.�#�{Xe�zy��UZ8X(>^��p�N}���j�O�yuE���ݲ5|���qw���a��������3��Z|�_���3p;��|z[{1P,��ňx!NEވ"HM`��Pc[[	ʬ����������R��L�d�Ƕ��ĭk�QK1�^�vO1��g�1�i�<�&#���_�'�n��I$T��k�OIR&셹Pi��*$[�~�a֝Ǵ$�O�'�����<M�`�"!aD�\�Ń�쒉���s�X+0�Q�;>ĳQFr.H2��g]����,.��2yWDh���n��M�g�c����\(P��b��bl�g��͉�cս7V1=�x���w�Q�D{�ΥWQ�;q�Q����6���e��f����K�b��5�{��/�S[c����S���%�lδk*�'*��S�Gea�a�TM8���Em��{~K{K��I�ۧ�efGb�v���]/s>��F2�?.�|�.�>)'�6~�����)]���N��)0!�`ER���	�C���I^PE�%�lmt�'�+HHH�$�^��s�5��d�+c���a	��yR����R�rJ�����j�;r�55'7���?��?>.��Le�b	��AA�����L����l�C|R��*x��U�$]	i&�������&h���5�0���ii�Ľt�}��Fg�u��|U�l�L.�k#�\�����Q4?�)�}'6�ժUR~*��m�C�&������w�����͂����},vg/ ��Wi�����T��{ۥ<�&�����`U��<�q.'�����3-�T�(�>�MKLV�L��u1a?�`}����ճ��c���Fͪ��̤�{$��z	�ͦ�F!��r�m;3�a���T���F��򖫳s6�����U�>T��i�VPǄNgG��ϴ�����;���0�0�5�`w��o@A)uvj�iM�~�X::P�|D2(mː�^U�W*4G�L1w\�s���=��Eh5�b���~�\'������r^��w�y�Z&��dGj��O��ǫ_
1,ΤF�.`En�̶낃Z�эˋx�]�4��-�R��сBY�X���nu����5!a�q��_�0�Vwz0t�U+�*��u7�����T�T�a�ٿ�r�p�����b貵�m��jΚ�S�|� U��lЂ~��bu��"V
�����B3F��ԣ�˄ d_�1��X���1醁^ø�}C�.z��$=N�#�`V�El�@�9�g�]z�5Z���$���U�����͡CڵF~.���J�B?&��6��>T��C�|���Ꮢ��_M{S����"gњc��OLM��(�����<��i����t�SG��
���,�@@q~�^��Z(wWQQQ�����F2�U�ʕME[coM�  ��_D�̐�yu����  ;��յ����Ce��<�[���������v%�,0n�1�xL�ML��?���Mϸ�c �R�ZE� ��#s�9�*���H�����&��Ǉ:v�6k�����M�|0��s�Y����3�A�'�eT${���]f����������OSE���h�Q�Mz5�K�����.���Rng�*3aVX��` �%��z��6� �_��a0&D��X2�E�7�g���+*�J�0rvX��e|l��4�ρ=�ў�0�X^t�Kv�Ӡf3�VN2/{k��c�g�}}~Ǫ�ɖ�-�;�@��z�upp��G�o�@�ǸQ$�R�{�������%���J5@�	?k�����G�|R�4�T2a�n~�Bv
�%��Of��h47N���s��L�;"�����H)���V�m*r�a6G��J�h*��\#�Z~��ʆd��b�����qC���9����َt�U�'�*42ߙLa�ox)���n��j����yo�0���Ƭb�ł��p�����.0[��+Cf�;��Tj?c�/.�5OS�3TiW�?uv�砷����^�̈́D$.����=N�2�瘄2+���V��?u�����m�׽_c�£5w�\$��>���)��*h��?�)��z.c��5�LC�0�U��6�ʞT\�	.��i�O�Gi�(,6�E�=�1GPI>3o�ڽch�~K-��`�~<�:���؄��\VG<���]�����4�A���3���O��)�U��m�� ��dn�*�С&BJ0"�T0��i�� ޼G�*|��`�~��Z��Q�"����W��\HTeL�=n�$q�5@@��뿞7������luȗ���Z|��ԯ ��Di��9��T
�(�|NV�f�Ɓ��f78��'vߟ3�����J��k��frTqT�ꠣs�T6�Dm�C�J�������Hya
���
��$	��&&��m	��˚M�m?���0'���杧&�!<��;�$X�.�z/C�S�Aǔ}��j�D����8cģȅ8��F�h�!� E��vn`LY�"�V�)?�ǉ�#�Y����够�����ޭ�r�O��y�́+��2��I�#.�Z{���	v7s�!���*/�zF���G�<��r��
�oaZ���?u���C!	\l���?��F��;���+���Y�~E�8<:����_��8�zz��(#��T\��Jv(؜&<9ݜ�љ�%a�h$���E2!@������!�m$��)2*�K,f�JneS�;�S��F�N����INˑ���'����bW�y��1�����W��r֣4-���8��~����)����[�Ɛw�]�wD ��Q�J�DM}��㥤��%�mU�y�G��5���&�Ԟ�,D?��UM��T��>1��ͱN�����P��|��[��P}FF��Wa;����Š��{�i��&�>��fn��v��{�i�EA�M�3%�06�5��@W�.�rAV�w-�v*	d���� '��Kݐ=�4�Z�S�X�0���._{C��sg��V�QYֺ��m�T@����Ѽq���-"��SuM���h7w�k�o2u���*����Y��������GE��T@Q�*#Hn��n��0Y�8����l1P���㯻ǐ`~�"�����{ypG��Q�?b�w<��v�H���+�~eԙ������4J;[K+�R٬�Ǒ���u���"��C�ϣ��؏�~L���s1�<�xO�PBtND�d�wS�OW�(�����rټ�T��n�����bGٮ�n9�K-�>��;�A46�rU+�>�{ʽ1@���D'�"���kqa�m��;�H~c�T<���ya�Z h�3?}`������8�a���?�)���)0'����A�^�T傤`�E�UO��zqKv����!y/c6�_��UX�XFn�wk�Z�Jk�Zn����̗�U��@�7�+8�&�W83��Ó�'���kDnVf���X�=���|ڵ|�_��v�r���O������JOwC��T��"zU+����! �.gCE�b}�W�L�0��&>i��0ϫJ�G������om"Yz���SLVJ���Y�:�l-�q����g�F��U&�⤤��,D$��5�5�3�o�ezXFU=����]W��w��0�B|���Ju$VQ�:�v������+���,����?ߜ��WI,��Q	+0�s�5�)�gR�2Q����~E�-�UH����-f�_f�6��15�t��0[&�I\�k��9��v���C!�۪t��.�)���/�tI�F<~н1�'B"йT�_�WljS����E#��E��%d��{������7�J�}���yY�s���+zj�oYJ�57�7��s}�4)������z��r�ي].Vo����\<�\�!*EB��i�ǅ�����c=]]�(}_~����JT�h�d�XD���	OZy�;_�p��ɏd��)%�!0�dDD���q��D������O�d�LƃŶ���J���Ǡ�uv�V9ypD���:��,��5q���K�+�!��-@�;>�hw	��a�!��y�#��*i9[R�4����ʓ����R�}������P��P!b|��5K5ީ�P����b���E�R3�?�����.h��h���|�f��|����Zn�[mN�����)jлT6i�n,q
���L<��\$��C�y�u�f0E�7*�߆9�`ܴ��t���(�Fi�ѿ����a�EI�ΩDg@Oh��2 aN�1(v��˕��b0-hDU&���qr[�keu�y��uew/�;/X�� �&���b~ƾQN��UeS�ޞ�Vz�o^�۩"T�ӏ&-�2%�$�N�]�cw���z�
�J��e0�mLQ���,�i��
�n3S'��&C�=0<rlY�ӒQ�h"�_@���Epi�V�xa��0'=yy�In�e`���
�1}���t�R����n�'�����f�e��� (1���2��uiL�����G���Б����@��U����,�m�R(���t�W�D��E%Kv��ބ��l26��\���:gm�
���r��ҖȈb^��'�H5J-{} vľ��|��������f�d�I6���(��7Pr�V��17I��<�}��7���f�=q�� �/����������ͫ6�~�Q'��ɴ<�dz�F:~���V��022�y)�͖.�-'_$���I�R��ci�5uD���	���S�r�z|HхB���*+q.���*N���|u�$�d�t5}��Rʕ����`TR.��#'ֽ�V���s������,�"jl����>G�*�c�l��q&��7��/�����iigxkA(*�KLJP�Z�Ƣ8����~��Ұ3n�뇎!l��p�.���<�Q��B��K�.7H���|Fggg1��������Tt� Dq5�~�BZ$>��O�ͩ��19�����֤h'w�
qtz'x�'mMd���PD��N,w���w�_/+V�y�����~�7��/��#�L#�������kOc������Di���y)�|�ݖ�&�<��x�&��[����.>�c����r"[L(|�kU<]��QW2F�ք_��I�ub,��<�����H(-kza�B��:�{a�p PVI���ݡ�7�	I컭Td���z�wʣ];PX0��J��w+C>�ָ�S��^OZ_*��]�
�ފv���%������V�ͮ�z���t�00�qB3�*3�a$$��	4���O�>��_�6:\}u��|&^y;����?����|�����9z\�Q^���9%&*�b8>��:��D�S�r�O��	ezԟ�QUs9�X��8�WwF�Y�A!""F�%hg�yVY�X�W�b
��)(�1緌��y��TҢ$Zs���\Ȑn�����{���m]YE��N0��b���td��	��8��m�$��	G�kP�/<[�9��d�(��x������}[�����j��1^/�i��|�ᑹ�n��/Jx�m@y=�k7��_�����E�dJf�����YDU �W�f������x���,�����,z��@���J�_dG9ȕ�AYZh�b���M��L��AL&�U����<��r(�A)þ�
F���5q����>��wE��m��l%���6)/�+Ѿ�g��0�iF۸_ȳx��:��Yd��u����A�owy>r���|$��;��!��c�����b��|��ᡙS����E�KB�w�PG�2�7;���+(2��@���I,���K��pTr�l"j�w�h�'�j�8�� �J=�g��&�RtL���|�x����EZ�/= ' s��-���BV��G�����C����~^cc=���v����� �*g��2��Ռ5z���x-%�����i5�V�!&�7KiA�����k���ӱ#�����S\/�g��9��/��>����>o��|*x�t.t6�h#2ѴaZqu��`"������L+�>��wY������y�@��8#.�[�	Ak�|�,Ax?d$L��)Kt��6	{�Fo�9�`�C��s��N������~@�و�e��pj����ʌ�d��I�	��,��`���������+�2=����	��?ص�F����Ȝm�%�&�<N�Șr��n�Ԕ��f�T2LQ@�DK�
���82�T���K�/9�����~�{H��@bl���ݹ�� �bB���9�KH/������ҩ�k�
G��;��A��G�޹���l�g����ϯ&� ��c��Q��f�My�e�b%����]�־o��|Vx�M<���\�]��.�S"֗<O���q�s(�	�K
��l�����W�w3�[_OO��)�W���r���v�f� ��-f��KD�2|4X>�!�e�c��*�V��p�`��9=�!#�o����~']��6U�k�� ��ĝ�ePF��J}����t���
���&⼄�VBN�^�+�:�]���o�G��u^�(���������#>��%G�Y�7����l����ԯ�&EYu�A�����T��	7�\+����ZG�l��,mFh�h��kқ7�V�F#\����Q�/��Wi���Y1�v�q�3(��"g�r��M��#�=����:�%�f�Q�.b� ��z�rtLLD%Aw��Θ���b�B��p\�@;���	�B�Q9��w�:\�
s/�����F9� ƈg��hfw�.���_�sG;�C`
���XM+���Y)�VT"�}G-�]JF�{����K=B��9yF"�������05��DT�,,��mӿFI��=�W�������G��w{L��oz��ϧ9ax�N�R�?�/�@���xY�༼��:pB̽X#��y��@#m�#BK�٠p+��H��6M6&�rHt�U��я��m��&c��k��>�����B���N�3���+����8ЗY�ʨ//���`�\�Vm�jmƺ�����c�U�!��wӓ�]�F��)Ͽ#�TuA����2�&7uR���C�fHp��/�^d�~> ��;hQ��`�|"��BQ����n[�Ō��m��_�01��BZ�ҁSp�	DQ� ��>�J�Z�w�QW��D�u��4�A>q��.	a3����e���o��}��-�%v[ ��}���F.�4�2ӑ=���1�'�ٸ� z!�ajer��ā����NHY<�rD�=�A|���]MXw ��r�}�w�C7����'�	7:p%{�*�K�1`���&�6�7�゜����	��l9�f�Z�J��|J�h�=�90X^+�U�F;y�>ѧ�ި/�SxEh
x��\�[PY����1_��#��)�^�:��n��Ϗ���Wu<��$IO�_j�!,i��v]������<�p��U/_h_�Ѭ\��7x:��3�m ���á�
'a���2�K����/
�m5'5�U���Z���p2�c6��D1����nz�{BU8w���M�gzm�Ky)�� �%�v���������w��vYC=�$ZJ[�t��\1��|���ɩ>$!{�4!��Y� < �Q0 1R0��P!��s�FG�`�äYD�8>w��i�����@Ǡh����]�G�j�G�~"�QT
��ZP'��������rZ��e����G�=o?��s/d^9z��\&�X��'�i=���$��|���y���^�ЪM���5-����描	E�p�V�G�cC��p~δ.��)#���Z�X�5vg �Q\�Ί4=\����V�LBN�ʫD�I�
�U� N�����*�ɿ���\�(]����|�x�X�ߛ��ݒ��_���G���P>��]�|\ǆ���]�]({)��JJ]��!('�I���}�O�����:��Yj0_N��`5���|��v�������R*V�4��]�]e�Y��!<��<q	K _���E��!]Ppn�^�2�"A�]���K:��q�
���ͯ2N��Bko�n<�jҢ?��Me����%���^�׷]��j��_4wT�U�i-^5�y�ia䡵���ң��JAWK��b���s�6�Җ��?{>������p	�MF�w� `�.��퀟P�st�x�)b��빋�oC
���S;�uZU�pv}�.:� }=�!\I Pۻ�$�1���41�~bK?a�	�Ѹ��D��1u(ۋ4�lih�}�ٿ5�� �=цPR��or����/��2�V����<Z�z��#+�U�C1�F��Mu��Pٹ��zP�����W����v�L�)�U��C}�?��:�X�����d-��e���d(�S�t�74�M�L\bo�k�D����m�Z^��.�H�,*�:���{��9+PT�;����l��������M�?T�E�)����������4rwCx�ݽbN��=n'A�Ҁ�&�0	�I���Ӛ��-rݯ�ӌ�aSY\$k[�~Kw����	�"}.T�sd��jJyS���L� ��^�����\�QM1�0a����N�h1��Ӄ=�����ow��ߝ�B~OL)e��`�,*�Dn p�c�C0����X����� ��2tFf������	b�����&�����}i}����y��u�H9���X��v����L���pV����3�,�O?dk:!Wik�3��ґܖ���p�p�v�g�{8NS��kg+����_����zLi�l��(�6$��$���%VP����4�H7M+=���l��'&W�ݣ������+��m��_[!@��w��6tv��0����0t%�n����B��Z.�l���F��3�(��#�'4�5���9��&,'� �̅��H*�Dn�%�ci��KH�]]y�9 ���S���Op��="~l#�� ���]v��'Q�X���)}�b�Sf�$D�g�Iw������2c�y�_N���u�R1���	�jT����`����e�� A
�;_�K�P�K���Շv?���f�=���<�:=HF?x�V�y�V`�Ä��mp�0u������v�9oO��Y��ʗ�����u�Mk��?���(ϟ�(�ƨ��]7B�3���~��A�V�5��� �� ��c,�C:�np�&qn�HM�����Ead>D��m���(�U��(�sAÞ[vj���k�Z�b*i����|�md�lGS����wG8�z�p�h���͖�N�2B�ſ��`k�� <�z�!��a��|�����t��U����
�/�	�!SJo>��zڍ����BZ �zO�-�˭�%��ܛD^O)N	+�i#���Rʾ�G��@ud�&\
x�c�xu�ΰ�:����<w��[vo��n;��<�G�f�YV��K���0��W�������^:�/-�LC�&j�	�@@aw[̓C�ҟ���r#­�l$������i�n��ƕ)7S��hT����� ���(d�f6��_ϛ7��c�є�W}��pT��fw?8z�<:^��h檵9��'d<�a�J�R��~�˪y���/�2����7�o
bB���<v]��e�R�w�5�g|?2w���P�8Hg8�pO���21�ufIw��	���Su> �B�쇤g��\g	��`#��&N=n�ii(Yވ#�������%lKXJW��f�2r�A��
,I�=��'����t��H�vx�X)�����G����٬AzU�G	��/��@B���R82yg��i���z�e.7�������W��'K2�潑�}
�F/}@�L�����/��uA#&�1��Qi]r��D�(��+u�}�.+/?�FB�o�}7�����ap���ylf�����#=x���R<���������a��,���UX���8EJ���y��٢5ګ�?��@���4蠅��ר�0�*��"j��<�a�^43�Fe�%JW����VS�FZּ[r�{H��!	�*9��X��y��i]�_�J���� J��K�mc�=[�"I ��eO���1y��{=�
��D�R�
_�OZ��]{Ugo�@��͂J�X�@���[�gI݅�6��t����C�^�`xU1\H��SY�>�ϔ�̛iF�Fz�p�@l�B��|D��b3��v�~�8<`����u����P4??��e��Kx×�����7�=��SdYqƿ/V��v�����{/�*��j����.���Š{T%i�2�Lx�k}��r�0@���I�$�k���1��Ux�c!y}<c�<�	���7:�Q.��H̖+�~��7*G�)؃�R���d��"D�@�b7��
5{�������k�Y�a��妫q��QMZ�X�5���5�fp5`>,���ؾ��'�d���1�2����}���A�A�b��W<���l�e���Fp�"7��O�fo���+ ]m�qr��jmM����0�^��BPDG����ط���~�?���{����a=*{�i�xP�:: �2H���1$9�阞3 kd�k���3�n�C�eْ,��&0"�]�U��t���$Ӌ>wew� �ݮ�5���Ʊ�5q���ݸ������1G����67?v/MIQa�������R6`���u�l97vGd�� 
�, "��	��`�*�2���*��lj�/���:Q��T��k�tUO)NV�Ĩ$K.�G����4� ��c"� 0�?^]?���?r�P��(�)�]��r<��~lv=rY<�q	H��s2�,h���c�*P�E��K�y&�&����5��q���t�?���>4���a�;�� q�}�YV��H��(.�B�(�F�9�liI�tE�B�ဌ�?<��Gb2����`)�~��w����J\�s|��޲�ь�	\������A�^��٪н�*�5X���X���M|�����փ'W=W������d[��諝ʕ<~�v�{}/p��s�)ۡ����= �M��m.}�69����>�1�l\2�Jv�����p�F9���VnQFE����E4
�1^4@����w�%u{��@�1�!�L��+;!h\���Њ�\����)��6�����	W���&�$�W�l���<Ҷ-0,a��Ն�{�I�Hv#��(h��-�(�
�m8qL����e�&�c�W�}ݗ�3��C�b���9<�����^�m(�%I����
���=K�ʳ�ym�qW*poff��e ��3l�L��*���W�-�C�D�8��$�	�Y��8U8e��ٻ(�MOAr���|�]烼��-1�X��(<�8�u��p�H� \,��w�(M�T�m(<m��&V�������Z��W	s�9�&��jbP_��,�k� �����PW%�]Hss'���CF�gŜF� e����65��8իs���K�����m��麚���1�z4�*��Mc��S�X�]�(�Lh��v�J��б�zA�"���������ٵ��n$p�@��|��Qt"��@C�������ϙ�?��&���f�f�����"�;M��f����ʁ��V�Zy��p�tH���G��&~G�7S�!��A�:�/�2�=���2�z��G�[g���EP�vf���%?���q��c���7h,�{�HQ��PZQ�x����^���?�?I�9�*�gZ��,��(&O�;��h��i1�J���`˹5��UG"X/�^��TU%fK'R��;��/Z�mI�&(�H�-�5��a��������rYV>j�|Ӗ�k�|`�Wc����p�
0��#y2�r4h���\Ĝ���*R^�U��������Cz�U)T��~ �W��*�����Ȝ����4���P����l�s��5lO�L+��Q��2�ĸMK����4S5���滘͑d��J��=�ײ��.�,���_�wu����3��L~���LT�+�a��"����J�T}յ`g66�R�!:
|v���O��٦�N����4OھGD��0|� t|�o��Z��(�3:{2u	x S/���z��B��e���(0�;��n![Uz�5��ӻQ~�c[��>x/�a�(#GB�:�(����7�,�/��f��F�aڣ��A�w��=��j�����%\k�<�w�)����^�3��:����&�7��r�^m �Q#���ϛ�-����,%6��?����b`���đ���������w��X���@g���[��gq�JB����b��ظ�[Hd#�@�ǣ��დ9�����*����Hxʙ���	h܁(�Nk����^ ��y��1�<Ly~���(ⱽ`���DG_�
!���g3�`@{��A���YJ����bb0���Q�57)(���Ԭt� LW��7:��HdѢ9�	��]~#?Z�p��`֎�a�)����q����hnf�4"��9�		�c�'��B�wٯ_+1pD\�9JY��;Yz��ge��Ilv�>iٿ�$Ӕ�P��9�CXbe�������,T(aĴI��|2B��Da�]�TYY9}�gG��^�Rb,ӣ�_m�S	��*��Ԑ�#���˚���Q�t�?~������:��Փ,�n0��\]^~�+���L4�������28YsK�F��ٚ��h���l(቉r� '�1>7kQG�g@c���q�91��ѓ>�w�{�s��i��h��9������V�T��/�e��kҪ��wg�kcuu������&�-��}C"��M�b�3[8�L�b���l��	���U��� !"���]��9mq��:��$�h��"[���3:��LM���,�~3XUE��Hl���	 ����Q-g�Z��s\��Ɩ��O_���|��"ݱK�(H
,K#HI
K+���R�"�twJ-�K+ҵ�����������;sΜ3s�>Ì^),�U�J�|�����0�7CN�o�UmS$�ɺ=�*����.;'JHƼ,�W9�7�_M'���D�I��C:^�^���8�jDj��:`���}Tg����c^��sț�3�l=�$�"�O�u	��ݬ�Y�G���.`d�܀c?z�.=#����X��d ��Lb+�D
kҲG�:�~}�&��',!q�<�wgG�'�l�������Di`|�����u��s�������i!���K����J�o�|n�mUC�u��gTg��x�_D4�����8qt���s�$ n
�{C�/$���	�ϖ�Zឡ���m�LiA�8�$$��H_n[K������mK߈?�� bŗ���s����8{���m8pՂT=��1]�1b&zV
���[~A!��PY���M���$9���#B�?z����Y
���@V��yr�|D��>u�����AW��/��z���.Z%�i�N�w�J6�4�b�����C��&$#���ˠ¯����_�/Z�]6��"?�Rm��>�
�P>	�z���E�d�m�� ?ϙ]츎����V�^��5h@���ͬ�������HN��R����e��J�E�缗FyN����d1�'�++X�|���E����^�߮�(D�^?�x�~��.�?0z܁�u���x%�ś����1��Br�*��	fbҷ�l�2svn����I�{q�J���g"7uv,�rq���짠u��эS�����4�`�
�o�WII!���p/u�h�ߍo�b0�W�Dq��iO��A�b�R~'��u����8l��3&ύo�U�������LHM��4ɱe�UT�nee�}�ܩ����N�Ŷ[W_�2Eu؛
��#�(N��z�I�^�b8Rt�zė�g���"9�5�����W�Uʢs6Ӛ���9�ݽi!�a���o���z������ߧ���H39|_R|�_7G� �!�����.?�/k�XP?;�	S)#|Ģ�)�V�;. "S�2�sn9��Ɋ>�B�$j�y	�'���vA83�?<����N��[VX��<��uB�_�v���O�Ru�Hym������&�dI^���gI�_��.�ե%�����������Ϳncc��,c�~p��4��6��2P
�,�9~6��l�̴�7U'.��%���<s#�\~:��X}@/J������ܫ�)�����T#<����Դ/$����ӑ���`ULʴ��6x$MN^�)]�|g���	�׿T��˝
���������Z�2�p���\���͕�/,V��* ��H�o �!�$��M���E��1��B�K���T�Ⱉ��ye���t%�LQ:��2�$�~Kop\=���1N��_x��R�A�V*Wq�V�������X֚�[Ϝ�6�qv˙&��ʝ6s�`jzh��r?K3�y�`˝�V�]��xHK��'a�̑09oi��~��q�XU�c[���%�-�9F}�J�A��]m�1��M��M�4����?�]/�w{0�ܷ~h�k�������$Nt�����I)��|�+�M�,*j��y��ŦG�p�&+1�����`�i�Ƽ��!Z�#�#v%�=��7Rj�'�w�F�����:	È�j��}��LE�h���"�`ps[L�
9��pQ���1&�FX�ar[�|��ha��<s�����ĉ��sV�{wnɎ*�q'�p���|�e3��@�$\�r�|��
�##���qZ����$Y�߶�n�r�����8���"5--c11�#M� ��1����sg�`��:s�޸�T2�+�ۈ�}��6�����MA��\�?A�8	���v_�"��'�p{2V(�Q6���@�y�*Ԧd���7��U&�{w�f�tSW1v5d�S�ԍ<Ǘ�·@��A�C�V��I�9�����w_d��ً���gb`�"4�g�#��
�(H�s��,]u���v����Ԍ��k(C�Ǯ��,������u"L@���*S�)g��V�D�P�Í�g�%�")
���_��MVI��B�x����?>+T���0�o��4R�Y���M�=�Yo?hp;��L����v�����'EDT���F��xP��U@ �n�O_���\8K��ϒZ;�;��ޑ�ޏS%����h:wD$)K�����5"�paa���x"e
>�n?�d~/��?>v~M���H���]g��%!e^���9�u���Y�*�b�^��O�tX��v|f��7SL_̣l���p�>�,�d\(�pay%�FsǤRM����^Ҽ>���ç�m��`��>G'k蒎�<)�^������n�gy<GE� �!BM�!��OW���m,pT��L�����-e�vy�����fEطϷ������� s7H����G��X�mI�"��5�r��ƺ�?U��s�wV��NٙoQiw'�)����*'��B&b+��8'��+B��^��]���=~���	zl�&s;Uq�Ф;�N��>D��pU�J۩�=�e�����u�K�%��j�3K/G;�����r�>��&KS��h�;u�?���D�/b��]�e��#�\P��d>r3l��i<��φǑ}I��vj���>�l�X�_��l3���VY�0�� �+1{�� �EV�tw�3e�-�Ga�;��-XN���-[�;�i7�	��A:���ϖf�*���c������~I?
�+�b[zz�q��D܎qb&0q6��������ɲ��#�4�TX��q�M�������8��� �;����)�%E}vr���ͱ��������%|y|��~:61aZrΩ	���L}9�~�~�(�]���Z�8](��im����@�����I%�%�s0�!�N˺���INR�	r"��ү�-�{��ݼL#ӑ�*|��?Δf�DH޺ ��/C��U^��r�$�
�>���Ma�%��0f�=<;�-&��ma���G�ৡ�K;�Wgiz�5��눡��Y��{��H����m~�4���JIh�O��g���|LТGA\����`~�DM� 	]ol���pLݷ;0,�'�2�KE�����)8�����Q�H3����\g�J�%���Aі�t�Jnm^�^�Y�fw^����T�fbN���x�n��8i5�x���\���e�@=v�TA�g�=�u2 /#lO�S���Z��.�jEDD�nc0��K���J��ZnU0n�b���~����A/����)����[Q=`߈J36�q���y�p�����}����]��7��Z�����þD\��o�$G���J�RO��<>aa@�&�8��)�����,,��@S�>Ca:�bG;���tx������"=��5.�\I�ook�_�#�2�мO�r�	e����>�L�~+�-��7R���g��z4q
�9�i
��w�� @�A8��5�����B �W-�I M��c��"9���ď�v�]��}в�@š��bQAA2�˚Y&}DWW׉��RQI�!u}ch�ȑ�3"�tk�v���+Β���>53�!��L��]�Och�Z�֦d]�2�`�a����S�1�	��e��>��gvF�etY?����J��7��Ū)�'�q��a�� �_�p	��s_�ʔ���3��|��[A�a暲���}�Ï�>�b'd�M�U�(�X�2��ޱ.1��Yo*;$�<C���ʪ/�*2.A��C� ��V%����<\���$n.��z9��w��!8��Jb�ssR�	r�K��@�;H̆uz�G~PY��ߢ�F[/�T~X������Z�z� �I�cê��)�F>NAad%M�M�8��a#�kE�2'�����}h �7l�C>�N*�1��w�@v��O����B���H�"-v��7!��<z�wo����j`S2�eh���3�]�r����~R�J����W����z��dS#z��z���T�v�ϱN��Egw��ُ�Y)~��ƬV�M�YvYR�T��<i��-~��}�߰ώOC�F��T�����CN�2��58�����|Dun2O��d�N-\���s�5󤍇�y�������p���?tZ��n���N�N]]�vw�ie,\���h��]F��7Jg7�� rv���}� ���3�82���(�4C8.�_D�>!�.j�<��h��ri�yQ1���{7F����K(�NN���еLP�l��s���Y�&��GA�F�)0x\*{:�'B���B��a���-�J��(�%
-d�� d*�CY�y}��C��־%���5ft�ft��[W�:ŐPI!�0�Zs�#Bo�D�=��`�{Jm��F١0�_yX����!Z�9}o��l��DK��_�N�q3e����b��+y<r�
�E�;;Ľ�ݢL�-��V�Ӆ�n��7�a;1�C��/ל�ĵ�[x�ì��'����["9��jc��99h�M�1=�	jQ\�z�^5��7g�Ϟ=[l��+M?�w,�1螖��v�_�4���a�#��r��b?��t�;�N��0S�&�6�	�C9*�Tқ��I�0�q!����[�z+w�^4w"�B�/�����lG���UB���Dt|�w�������tW�]BL��o��k�~��e:iCy`�g����<Y}8���r����/�%h484PVROߏ��Fu\	&���%AV�Ny/��C�C��Y����E�}3toߠRK�2T�c6�:��Y�~�����<QŴ�<W[�]̮�
�g�����"��g�1�ئV�D�#F�Xюsy����t03����{&P���=���y����"�%/�#6P�o��fVObL�Q�s�yIGI��3���}��e�o��R2`xAo2}X�)I,
���p��#�չ^�������?U�fkm����_�P���W���%_�9?�2�Tpyr^'~\�B�ʊ[�(ol��}��<�])Z��F��ʩ��X	��{��,;�ԙǘ��×t<�_�#`�z�w��(�6����( �|H�vw!`➤�j�/V�읮l1{Q,?�CI�թ�Q���&`)�Q E}��0������5����U��yQ9��K�I�KQӂ:x�{�Á�܅D��n��f��g��tR������Xh �S`ˌ7�zb��.F'I��%z��n���]⎷� x�z���� �#V����6>gՅ9"��ܳ�9�*+�?�VV�Ϟ��r�ejkI�
�=+�̻B!�& ��p!��/7��~뛘�O�r���x�F�?�S��W�X=�Ѫ�Tœm�����c��*rrr���	^���a��"|p�irc�^��)����HX�#�Pěܜ��Ɔ���rU��uf��k<�g�e�����%a�z9�'���P���KIU�V�?nfы*�,�]��"�ꐐ��QR*{����,O{�� ��N;F�sC�ǴO���f��m�*V�*�.n{��vƞ��UR�+|�upx/z�$e<��5u,��	�]#����;=ra��.�/��e@18Qu|�6�g�fj�8�ޑ>3c���U��cI�;Ŏ؛���A�{Q�X���>+��������ظ��֓����sU������i����T)`\w@���%T�瓂ZI�!�D�P��T��ˑ�@�l��
3ێ� ��� �.����t����=aέ���ˑ��Ѕ'��l�|��������d'%ѿ�a%�r�p��>�ޛ�V�h������e�t��%u�e��#�i�����ر�V�g%�m#c�i�6� �)*&�F����@ۋ i���fu��v����g����b)��I�:>k���3&߫I����j��i'UJY�65#M�S��A�)w�}���?6��w���Qv��>��)�*ZZ���6����������ޑ��5NZC����{evR�E���M;�3��Bk}�#b��0� ͕�B=y�\6g�p��I˼e�'�r�o%�ȲV$$R�9յ��h4�D?�8&;b'ѥ�~�Y�)���Or%ވ�b$5-��&'��HT�q�g��׶PѦ��X����GC Q�px�FϹb`cGI�	������'�&��i\��b���|%$3̊ A�٥\��r]��ق5��)XDN�5�2�m=w?Dn�sP�_��/$dffB���e�w�Z�3Y�]��0IY����x���Y�h�cǃ��%;`��-8���kl��4�p�%9��$�A�yݽ̙�\9�7����Ta�y���<Ԗ{G��`�@�����u(�y�0��YAJ�|0��T���8��O�5�xJ�uĹW��<���tpCz����`V}��)b��J��s
GZ~�8|M���S9t�dv�Mcb<u>>���P6=͐�0�1�aP�%𐐐�z2�5�8`�6"�π
o�	�j���A�U](����^��8��%��P���"l���X�Ia���!�*Z����mF��.����$�^���Qv~A�����ή]l1&w��I�b*��ϟ�;΁�b��������p{��k�e�q��[IGe�{�E�����o@W�uq��N�<[�\�\ �S�D�I����:��S�H���'�5�����7I҃���k�Ҫ��r�'m��"S�{��əA/�);&��9�ic��S�I�t��"�T�X�jggfJt~���c.���u����p�+���8Et)3:A "�%CT��Ɨ}�(���vw��OZ\�i����Xg�%�!�	&8��	a���ذ�������d*'S.\�qB���u\$@�4�߹`��W�7���+����S��8�n���] @���v��X�9U�$�B֋R~����k��l�H�����d�X�ԏ�a=��� �]CY�;X��wZ�	g��iZa�8����!�a@45�Iijl���O���ܙm�z�R`Ѧ)PF���^�>V��� }h�����V����ulf�Lpw�2�܍�f����-������}3p� ������n���'Oz΍3P����?�d���'pr�����b�L@%�5(���?������H�l���m��.�t86� -��ځ�	�A�q�nьS��K���,p~A�<��|�%�9uJ�`����l.���~�\,��,�~��P-|�R�K�ݲ�I0ԗ�5<������z���z'���gj@M��%�H8v���ȳǲ`���y�}��ﭏ�@��F��8*#0��"Z�-&�چ��Y���qk8�\"�C��s���4P�PEEN��$͂%b��EǩqIg0w-��
;t�dD>��|9�Z����l���%} %2ܴ����C�~!��/�8�:mN>W7ťt��M]
4ي�l&&?	�������X�ȁD��rs��hC��ל�\?~m�{+x|W|�������q�(r7C�[�_`rM��ǁ��#�7Wgة}V8�?�/"��54�@��`Fȥ�q��o,k�^�U	�0�5�P�%
zi����Nc����}9��C_��J�!�7�Z�u����i���F5_�f��7T��,7��V����Wbi�n�L�Ğs��~�O��:�e�yT�Y�[�`�~ �e�
#����dw����k�NH��2�l4�Lu>�9�"��ji���`D���%��&GQu:$��������O�1xa{�$ �^"�-8�j"�B���@�ݚ�,�ϔ�}]K{)q֪�
[mb�xss����fS�ː���)��Vu�3K�d�
�ŁoO	Ϋ�Q�H��;��E-��Γ�&���/'�}�>8Y��ON$�"4��[�P:+�6�.��=U�8��5���H\?;=�TV��_�����F1�_����_�U`̫W8��/��[�����]kk0!^8��T�;�h���^�bkd��<b��i����VK�S���$���0O�m��ҏ��S c�#�`H�փ�P�~"z�a��o�Z��4���t�ɾʖ#�V��UNNBv��	��j�[��>i���kfH(UWm��+��W�#z�v�1�w4���o��2O��ˠ~�g����;n�H��tvrr�#�e�'8�C;ِ��N �ceSa�տ��A�#ʢ��#�뜆P̱C�z��H���R$�:��w��ks��]o�-�r��3K��S:=��� A+)������ɠ���?<Vx�r�-��Z���\߻�{�_+b����Pe0��K�`?��3G�}Ѵ��ب ?�����e�W�^@O�xCʂ4�ȿۍ�[��M&g�*D��@�H�';� _�S���q'��)�����i�*g����O'��K�������.B���F�3bB��*Pk3K����F���s;Z@ӮH�N��DDO���g�N��Y�~����vt|16��05�x��f��ͬNI�I���`�l�EZ�b���<����~G߿�,�i(��k\0�������h؃Pji�G� �[��_���K�j�^�<�<Vr�Í�Ǹ��B ����52���*u�.[1R�h�i�o�E|��#Q��ȔXr��'K�����0����ϩ)>مE,�:�O�29���U�2��5�hk9�������,���oAi��$�~��i�'O���,���pqB�u���� �2\�dA��Lm���$���-6�*	���d����Xl�����l�h��dIS���=�<�'�~ �{�'Vݽr�4����QW��>Q�$�U�?UH8�#i,��p	� �O��ǳۺ靅gB"*1�[Q1��YR��i�$b�1�u]{�����j;�>�-������Ϸ5ш~����y{�f����X�'���.��z�ݐ���y��{VA'�Jx���:q����zl�@
z\��^�e��{���>�,� �87����P-�rV�� S�i�|��ӊ��[t�}Q_���\���4Y��O���,n]�)K�_C}��"{���������N��b*{�zaX��EĎ7��^}�D�hy�2f�$�"$�¿c԰q��eo��b>>������ƭ��7.�ݽݏo����JDl�P��xf�_SS���+�OѹKn]u�ހ�V#��e��A+3 �U���`�"mU�
�ju��aJ�в��_������;3�7����0�Oo�4 I�p� ;h��ۘ5���km�֙��=ӐފrsG�b��.���p�¡ ���g�;�]��(s,���i��G�gi�&��~�RX��ff�q���q#`�Z o�ӗ�/hW��+f7F@�=�K��%	��(\�Sj�Xr&��t�ҷ�����(���j]ֺ̏Ȼ���;H11�0J�`fZ5�M{�a\־�����1`�He��1zJ���K~��)dN��J�혏��>�Kof0�w��PNe`�L�@�wkFX[��M��AO���t�o:#Ȫ��M}�Z�6!�CxE�˳Fm��FG�a֦n����T�o��V77;�����?2��W
j? p��Q�%hW�� kb�DТi�ހs�%X�F�P1�>jZS�%ħ��$f�x:?���� �q���{2Q:d�������0�p���,����/bUG�a�x+���A0�s#��׃��5�rL=�Ұ�ҵ�'��m��r�&D���z&����~� 7<:ll-tx>n�Ү�M�H֎P��1��m����s���8����q{�7K__d�Z"�ǿ1����V���~�S�PZ_�3�۝�P=hܟ7!��Bg�G@h�;��"p0��wY���x]=�D�Pr,��ԣL��CSX�.��ކ��[:99a�'r(���23�|H��4(��L�`��1"I�o��a2��3�����"`*c���J�Hm!�P�<g��;`��~�r���� {O溭�5i�sb�K���ݜ�R�P�HC�8G�p��p��V��4Y���
Q �Nx�Ao�(�V��#��o�L�Ϝ���a���:!��5�ssm�bd`������{s���p�x�` D�:Wu�B��۔�"��m��VV4�H�ᦌX��mB�)E�·ʃ��n)Z��p��U�X[U=>q�Q�5 r��W~���ۛ�<�?Ԛ�W=�Bq��ެ����$~�����wL�#ݾU�"U"]���\�L�㢁�l�#ܱ騇o$���n��e��J�ާ��~~�̒���*����L�������q��D�<b2k�_�\5��7�-^��-d0�F��b�!s̨�H�88"4�I2�U�S����=�b`�'�]�vEU�j�#�E�Qr�f�hNa�Hq7a�e���)}%t�+/�B(<ñ2M�*0�;;s?�e�����	W�� '�6��iϽ�b���/q)�LIIl|��X
-fm0ף�y�P�5�"��%Xm�k{��8{i�q�[�W�[ c]^��zh,o�wk@I
00�ː`\Ca	�����3I���,�̔:̔�t�(����7�Њ����=�ߜ�E<�Z�;X
��X�D��
B�2��2���ڐ�����v�X|�aM&p����[ ����ײ�^����O�g=lU����30�[??�)�R/M~��?�Ѹ�zL��^@(�\�:r�4}�Q��	1Q5c/'���mt* ��űbr~W�u�������xS�4��l���z�ޝ�b����=y����[ <��*���ס���`#R�5�G9�D�D=�.��9���;� i�[q�@���=�w�A�69�#d�2��fc�a��<h����ћw���+��'�!7^T���m��z�����3g`k��=��1q��OfW["�* ���<��ά������K��x�oO�|��K��V
�͞�vH�N���ML���4��?�&+bi�~���ͬ�u��w%�i5^���:;c쥢�P h�͝_��ޓȗff�p��@���ׯ_��tvNJ%�k�M���n��SX/'v�3|�1��S�y�I��/t���z/!I������\do�o(+c�%x˟�D��V��yf ��]9��
�zj�����9R�p�I(�@��p6��1,����j��{!Y��ܸ�V��;�B1 '����ؕ���|sb)yȓ��f��u���ۖ亢$D�K��f�4TFS��fv�%c�e�r�	��$�^b��	ڨ�w<\�'�M�Z���F�� '�A���' GW�t�#�Qd���d��n�{j$�����֮�D�\��:��)>�\�g
^�؞s�8��e��ձ,��д���í[��gj\._�����H��P�������?u������W��?U*����}-�ԸƆ�@Oւ�^��-ۜ��/wXIM|�3k������Ίe5%��#���&�#R���uݯ`��W� D��b������$�@�����"��CA�!A�v��V�D�d��Q��f����G��cH�v�����9�}X+H��f�D�ǿ�E��:_�F��b4��q�!��;�M��h��}Dv���ySܤP�BFIS\�Gx�ɸ1�:���K�Ui�>b��kv_�Ukp���1兪:�d�y�ĳ�´�ɊyMi�����h�=y�< S��	r:69��3���sI''g���S"_��A�Q�<�'L�)`���-���r,�̄)y�[�"O��;��xjU~=[���s���qC�a����2mH��fz�{�d�� �b�^�Ó|��D�)����8x{���w�r�uӣaM���B/�cr��b�?�"��t�?!��Z����*W���eq�Lsa��>�-4P���%����ٙd���2
pFȘd�|���&��m�ΐy��/q��H���6�1�7$ϴ��&`m�9�G�A8D��涟J�<N�'`�������k�D-,=IW��aN$Z�
���ne��e;;;����2s�U����Y֞�慇T]�uua�,���<��K�z����wrG
��خmR=Cv��+�ʦ;��um/��;I���b۫j��''�������}�����k�W!p;w�8����P�&)�����-~�&4j�f�um�;O�����@��i�db�P`�e6�^pU�.M�b��R*��c�T�iK���K@�)*��&���F��xffXJ¹;�߇��4���kϽ�<��w���lUbaY� ��>�ob6����	}D�Ӊ���ϰ>p�Vj��������\E��pē^���RԦ�*s�+?�r��d.e�j&-����ѷ�*W��U6�6��R��~��l8V�������Sv~�&��-����6�3,��Z�U��������V�ֶ2�)��&�.�cXd��d���kk"fC�BN"��"#�����sV��Cuu�B�G�����܃Q-�87�H�yꤘK��F�y�կd�`�0�Y�Yku۹̵Z���䟧�~?��*L�:��Q��A�3S�M�JR��갫��TsR����G��˥(q�R3�%%a��T��4�B+r0[��$� ��gV�	�ߕ�;��zA,� �Y�J|#Mt���8:�N�;�-g'Vz$�[K�ֿO��Ya�ᑯ��=�)�!�r3���M��a���'���!h��X�h1�*>�ީKХ���{%���4���l:	h'<TOş�WѪ �h��;#م�8�XLe�YyJw
���/bIH�2�����~@i*�L�\=���陘\�2��7���|;O�&�#�>���Y9���������������c	I� c[����̑t5a|2��QLO蛊��R*�Dx-~��`���̓���K�Ix��קu�4��A����*��z�Mg��w2��!��ܩ#��±�W�����Z�૾dB�E�����cb�����Hm]���5�s�I�?��_o\S�3�(E����ݗ�{6��f�^�is������dH��]�á���a����s#?�����%8�]m�ݵ2����0�������&=eB�"9l����1r:+2�Ն�#HV�W���xE���^��@X��Ť�� ��s�����ҫ�.v�xt�s{s(����"Z�(3�3�$������v�YFu��)�[^}S^�>ѱU�4;"=�{08�k���Uko>����*-��:%�}�������|||VI��Α���n��t!-_��g{P˙Id�)��7��&_zȉ�!}]:Iz
�l��x�2�A3�����C�e��*�Z!l*l�������!aγ&8ծ�,�����I���i����C!d������^�2e��ni��
���MkC!�d���\��+�-�(y`��`f��2&�������5�i͗B���j�ϟ/_��%<7ص�,��2l8/2����N`�^[���W��z���8�Oz��N�M�����@��P����$cs��K��f���
.U�`���K�Cu;�����b�bK>sۏ�n�����S$]�0Y��/c�qpv֩_��2I�l���L>�yh�tK��m� ���GJ}�c$>X�&��ʧ�����ʷ�����YA� �H�ΨE�`N�j[ޑ�|"l�4��;�V�T�PoMl`�W���P��r��	T,䚬��]�?�\y
\�o�?�n�nLG�3/� ��Ù���";��}�CPJ�ٳ�t��_m�8�F�u��yC\���~�`a���ŕ���;yu�P�l[-3��<>:�WF�4 9n�2i��ח��8
�����i�ף���/�<��V��z}ܗ$c~I�_�%��Sqhn�e�ǯk�S������=�b�7G2i�?"&�X��m١�5M��nh��~�s��{<��?�&��{_/D��a�� !7��(�ܜ���=2�Q���)�[n���a�»�hn˯}�K ����L�+$�� u:�w�73�#By�9.�n��1�Kf��a�<C���?���݅Ȟ�В�VK19����-��6���Ȃ�v\�.G��[��B�{��\�V�n��
I �"x�wf�V��D�L�?U�D�m�n���r���&`m�abb���Zї���a����7�����wz�O�m�pIʖ����h��P8(D��reڎ�h#g��>��	?���;L�p����H]]������O
``�@��J	��?�
��$`8#����CD��џ=aL͍�t�րd���ol������s��f��`p){�+2\�Uc7���^h�����)�P+S1?��2�̱|�e�i�iL��O���fw�ɛ�Y�,eА��oU�x�UP^��y���>�<H�k%�z���2`������,)�xkK��%}?��r�~� &�h=�y��8�vD^5!���Ű�X.a��I�s%��ҍ*��X���];�"�j�Dh!7pF������.���
�L�r�����W/�F�>%`��S"��������B!{��E��ϒXIė����W��lj&(��/=�͖��!BT��5K�_�v��Dˇ/�gn�V��і��(D����Ⱥ��fhp�-�H������/݈��Q�?�;{#v�Ω�y˳Mڕ�e��4]'P{2�����E@;�G��Se�z�V����Qe�O ��$~��B�5��]Q�t�fT|���4%,*�i�>wj��	T��q��NH�8�` _Ah4E+c!>b,q��8՝B=a����O�ږ�7��Ǳ.ѣ2bc�M�'�~�`៫͂�z+G/��U�:Ǚ�ZFA����,�,ҿ֛�����˥�A�6ۡL��_����;�{6}Y�J����6Ie;�}����~ی��QlR�E��]��?�>��Te�q�;��3�"/^[J��E��X	����H`������`d�*�`{�2GI\��N���ٙHeU��*o�1{ 	����s �����_E�ݱi����9�Ы��*���� 6�U�X쐑\ÿ3���F����6!��o%$����Z�!�MȮ{Uc��s��|�)�`<.�8�&��hO�+��!�;xM��d�N�!�;�"1�	2�C�>��T�� 1w�\�yM6V��*�:h��e��ʔz����O~�hV������`j����0�D�k'���'I�Jmb6F�����=�!=�`f�����x�aZFs�CG;i�-@W�ʋ{|��S�ۻ��9փ�&�Jf����
�G��a0lOOMn��_h4�gN)85b�)�[9�9X�1��cd�ȉOa�;��O
Q��u�:�/:^O�T�.���9�����J�ɝ��,����:��E�������J�{����B4;ц����)Xl���I^8� �C� Q�֎�J;��/���F�����4L���ž�O~ɽ��33}i*�,���a3�䊌���r���z~?��#կC���Zܡ �'5�Z�����Q����`<k�A<�u�[*ޣ�ɩ�x�A���EN�a���	o��c��D����Ձ֧���$� � ق^����2�Wb�^Q��kfk�e}�W��f�e|�%��,��t�DDD��N�6�����x��3�'��ٱ�� ��)�קzd�.bC��I��3q-����)��ϟ0k�n6�CQ�ʑX1 =�����2�/�%��	z�gz����Jx�(�a=F$c��N�`_{�ϚI��K��~��U��W^n�����u���q��+�o^c|�1-GӺ �`�/G3�U�����*�F�E��� V�7�A� �M���m��{U�Z�y��L�.�jtjm�̰�qg#9:V�o���e�t���L��~����r���0��E���������#��
___�fd�a���-5+w֐h�}����'��>�����Өo����'�c��s�91YQ�����#~U�:���F�Ұ���چ��T>_|�s�£S�[J�]n酢*��u����Smr����� �0׵Vk4s6DJ�t�[r4����M(0��x'�?���9��R]���t��o�G���,�S ~�/��KЕ�$WHLR뢚D�kB�b��:8����P����I?�-}�7��T|��#�U��Z0i�#�@��`~v�H�{�9�TN����U�>���J�L�Q��Tڀ8i ���Na��_`��[����FN�K�ڊ�I��Ο� ��h�������y��ǉD΢"J=@�f���'J���
����^<�Ug�������<��9

#�a��~�3'�̚���J���" ��3,���Tkk�p�wyrLLL��r����:BDhO�@#��c��w����ǥF۵e# j�366�D.�M%ka��7��gq�<R05�J�Pu+��t���#{�R�o6W��8�]��x�#+����a����v�ϓ��:��o7�����wI�e��ݘ�~�7���dm�hŤѥU��v���3����W���	5����@ Jnb�K�������\�;\��/c_�=[C�����!!�f�kT����I!�3T��h�o�mlc_�Y�bʒ�f��/��O�ι��<������\��r�'����?��tI;ߵXc�˗���B{���Kk��G����	ë��ݜ�l�ן;�Զ��X_pDtd$�L����r�����dW+�=��X�l���B(Z��P$YZ������NJ#�/:N���%E	��a_' S"؆�+{��S���8�!�Đ���7��Qh�ۙ��fEg��}�~n��Lx�G,�Wt}AӒ�{�dV��LLNF
j
��sfl0KQ=���g�D?B���yq�����ͭ�@�'4/9��5��ը�m���d[������+R*ߗ�Lr�G��ڪe.��+�$MNVMLL\�q��0��&�8<��J�ѩ�p�*n�ų��r�)��������
=�u��|6)�Ssc��8�~q��|_~��w-
��ER�r-�)|�g%�������_�I�v��r"������$\�ִ�5�I�y�1����a��M�H�ZZ��������k-�nf}�����%u؈�S��$z����0z�Mq��18K?��
R��UL�@ϴn���2�����t�#�c!����J���v�2^��3�W]�S���U�ƌ�<'�"R��u�$�`�����RY�GPݿS�CxS.�|�<�/�+xpsc#D7��dl��rJ��(
���g'W��@�ԩSm8��\g@�+k(���������2\H�]Z�������	x��92;��dd��*M]�t*��ܴP1��O��$Yi_�|ߕ�<�ȡ��=���>@b�H_QG���da7S���H/�'��JZ��KB��o2�� ���7?�����`KP֬�P�
�9�Y/77���!&���:�2b1����}ݣ��1T	3������a}�Kv�RF� 0��0p�RYi���6�{y��{��a��hǀ�uFg^	�,`��Ā��C�/Rh�{��r�� $-� J��&�y��,���w�'	W�w���E�ٚ�����[>[Ö�ꎞO����F��2�ooG���<Z��9k[u��_�`w��C�yP�i�b�˵Bo�1�EN#4��4*++����!�N'N���;5V�ߧT�z��o�G���~��A��T��*3o�B�č�ì`��ƻ"��vHm]�������j�ӜI���b�7Ό��`a��\� 8��^�?N߾��(��燰٬Ma������bu�~�ן+�f~��z�9݁;$��}�]3.�DE��P(�s����7�P�20d�#�4�r��xѼ�������l>=��Z�n�	*�P!Z��N���C��y$�:����kn��%,��ZZ�t�iB�)���V��(��򝕺���,��	���_6�e�F&4nU���d�J�h�MW&��Yh?�n�۠9��_���E5��H�� ��ZDt��ŖiGM���Sٿ�c��l2o��|Ҭ���(67�{�xNp��Jբ�Sj�x%�H���*�,���bUY�}���ɼc�j&�i�K���duU(�犁ڮ�V��?���xD���`�W�z��+��UJ�5���E\\|e��<�[3d6}%N2��d��Ze�w�����۵��O�k�>���ц�"�?�ʈ�w+5p�����P�Xl�9;�(1�����e�`R?�7+a+�5����8^�Ul?����ɧ�l��ה h��?�$s���;~��&q��M\TR��1�j��&���xݿ�����o�:
��AQ�ݙ��[
�C	���+�)MA =wk7w�$/��~� a�ؗM�~%�5���]],=
-�Kr6��.�Z�J�����X�ϮPD�G�y��Yg�`O�_(*�Y{��g�"�X}.@� ��p� ����C^y��LD��|�hm��'��*�ڣ��"3^�չ�#��0�H�P�`04�Bi�Z/��.FEF��>��eQ
�?lkk;�5w��ܧV�6��z�^��a��ҥWR]J'���)�@Ӂ��un�B�uN[��:,ɑx4���~���a��mR���^��D؛��,�1�?-~�R���1�7yȓ�wh�����r��>	�>;5���)WM*v�?!��l\��y������) �T��`;Y ��Ӂm�����y]�z\���7���X��
R����݈��П�rj!&��z����+�{�:3g �c
K�����������E�"'y��Gl���/o&�3d�R!��yq����F��C?&_բP��r76�X�r?E3ف������ˑ�̥n��bi"�+�?B�8x�:�BE����I/�� =ƭ��?ܼ����r;RzAZ�^/��?�'z�KJ�U.��Z�N�P;��d�q
�3i��ف�Z�k��W,{���HCͤ̾5��Қ<��%�������(=� ��7h�<%�Vu6��l�cl�r2���')<�|Ea��4��=kN(�J�Q��p.A�i R�St�j2��%Gg�m=)*}-�ޒ������w(x�`q��ux�=�~��Z�9::Z�$�F�lGD�b't��-�)��@9tM~9���z��8�$9k� j�U	x��N�l�r>~��?~D�t��w*�7���^r!�2PCz诨&SlԈ���꥘���(�&�*�"��{EǦ�B���͒������Й�A���#�.�~�����4��O"k��������Лt2�A��ŉ�W����U׾��R�d/��gv �T����^|�ɲe��@����hRͶ;z��%O�"�;������A�@dt] Q؈:Fo{ܷ&WAA��f&H��ѣ�aҫ{r����Xm*�,����b��"��	�^堔��囻�J�?3����/�6q�E?׌�幹���s�]�F��j�V�!5�un�&u8��m�o��%-��zR%!ﺭm?��c�p�BC#E�^��m���Z�LC�������]0�λn)�\�TC�N_�`��_F�9�r�7�� 匣(�tR�@�u3@)��[=ĵ�7�����T��ݪ����wh�w$L-�� d�7�ZSC�<Pf+da垢��۞'���h�zrB�r��dİm�#o����|��!H���i�~���"ɪT���/��q���5�����K��6��`�2��1�	B��k�A2�����p�pc�X�>��%��(���+�l�#U�$'!@�8�0�B����Cs=

�|x_��^޵��/%���  �-v*��f����p�f�^ղ�ݟ��������F13�<����w�gpBx�9��ȕ+��L7��\����*�EE___
��V��iB�^L�6����#$(��-�l�h%���t+  �u�C��!Gor6�44�h���Y�@ ZX#�ȟ�_F\1gx�"X��(`@m_󟠀��q=Y���FY��e� J��з[����"��2=�#1.J��8����<eL�y����*�����؁({��3�=�nnVa�=�&�+8#��v�`�-�kd���Hc�TCT�U������؆�����!k��hE'��#�0��:ݧYx�Q�N��t�9n.U3��踫U�b��]�:��8�L̕���������_��2��R�^CL  ��7�1Úx&�PK   �i;Yp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   �i;Y�ɯP� ȉ /   images/d509810e-83a7-410e-8a4f-883955ebe6e7.png�US]��q����a��n�!��Ƃ������F����;ܜ[����x�jUW�5�Vw�9�Z�(/���� �,%)�~���_e|q+���, ��$<#�Vu�?�M�]Hbn�/��8U?�=�g*K����FJֲR��Eus=u�:o2���"m�~�r�N�/�I�
 ͛�i�-]��RYm?���j�q��R^�[d��$\�!�����jZ�^#����������.���>���M��
f	XJ�I�ߊ���=#���?��+���'�����	�'��*pN^o�3�^:cB�bj&'�=h���?�ؑ�q"��D�{t�[~ON6M#��b��ؽ�Tg�H>���7��@�Y"x���,(�?_���_�g|�pO�����頦����T����ٿS�_�&v`�N9�'~��ҫ�:}�(����i���:�����t�߈8֤pQ�l茷�A��{8���r��::@����=����� ^a~�9�|[��$!3������R �������W�	�$g
'N3O��}����`x}%�]0�C����Ae��Ķ?õl���+*J��B7Ý���.����$���ǀ��k��K�Ǟ�[�웹f�f-cN;�y�wlr���jP+��SX�В)��p����MX��E�gϝǩ����e��+мvs~�!�Ű�3�}:���(%yEM���۫�"��ȓ���76޻V,�{T�[F�Q�8����W���8
���;aɾ��؇���}"�@DI�i����ft�<���L��կ����3_F����}�߱C��P��y�`XH�Y��H{��k�_�K���Gi��wI�O�Doku��cf5�=�i>QF��e����̭���<�9";-�2�ϡV2x��'0]u�lB�Ͽ���3:�6s{w��I{2�s���]0/������o�\��a<�bpXR���a/�����0�XG��7X��#�CǸG߬߻L�����W'����M�Ψ�l|gd9"�h	�<��(.Ż�N>��9��7t&\�T
x�����=��1�ЮS�Q잝��E�P�M����7��2�<��k:҉�b}��JL`P��,Pz���85Y'����c��(��x�D�[�T��ؘ@���k<oyJ�*+�:�$�����Ӻ�S7"�d��0p�읱9��%�1.�����I���kdd7�R��L'�͙j-
�,�J�[��4y2)�*������Y�03_�UYG|~�K���Ekj�8[��uQW�a��>a!4^�Хo���κ��N0�����V��h��o�2������g������m��}��:�Wɝ���Z�,es2��i�|f�GҔ�ny��w�bvÈ��^���ex�܃�M�0�4��h��|�����#�s(�~{s�A2���;{�y�b�h����#���jص�zz�du��,�2��|�]�J���Ȼ�^L~�[�zDr�=�8���9��E�6|.��T3]��zq�!��zrh6x0+@�%��_�maG�20�S�eXIF�k` �o�7]888�:Y��J�ϯ����E8�;��1���)}z'�Ү:g��x��*s���!�Vf#q � `B�����N��-�4���ю
g�U� ��2-�! 	��B���6ޡ�}�����'��Ǐꥬ�\� ��������@�kN�^ϑPU��[ٝ/�=>�(�󕑋_M��1�6\>^�(����R?a=|0zo�}�-K����{�D���S����W��i�C���c��6�|�$O���u�j���]�dwaF(b�m}�%��m�=yK��P?ł��'O�t������'���C���6����ӏ�$�Ւ�{��|��]wK���t^}��Ε�E'�oq77�g77Jt�(a?_�=sZ�pxض�PaaW���>9ҵ4���'�������X:���֡�U��Ezf.�����E�����FEi�G��4=qa[|����~�(��D�M�6B�^�����\Ɉ�ʹK�F:!	�C����=�X$e~ejk�Ũ�wC;~��P9%����eX�%��\7��:�j5�.��.��23�F�拴�QC�K�N�g3����D��QzrP8::���М>�U�״̐�(�F�à.�{YJ�\h�]wQ�WWC����_��\�^^V�fee9_o�:���V~�C�y�ڱO�׋oVy����l!z���{ʒ���'�=eH'���֏.sDM)ď�c�b(u��ŏm�ʟD�^ZD��%<�ֳ�w /D�q�PM��c�ϭqM�y6���3�/e�k/٭ L�`�}���ѣ.��ڧ*�w|�;�P:.J̮g/��m
�[ �וJT���bY�7+�������ofy�m���[�"YG�ՠe�]y���4���踸~BCC��yA��33~��"��X��=\\n�m}0�O=��\n���Ց�d��<\q�ZuXߜ]]��/�����1aue�`��w~�i6[ XZU���^�Օ���k�̅]Dp�j�'�t�s�gN~= N���G��V����x#F��&�O6h;��= ?����&��������o���'�&�s$>��ZJR�^��9ZfBn��%ޣ�&���<x�dr�t�Z��ɡ������%���2��3��������m�GB���.Ѳ�f�-U*�F2�j1�gՏ�+G
],�#O���8T�t��{r�f!����`ސ]���Y[WE��^�LL_�/n�^��(GG7W�!���GGnȸ�u>�~�S�G���Z<���'��P�\������a.o�_W�����O8�KU:.��ӽ&(Qċ<��^�����8E��j���O���z���FE�]��ҥBi|rZCX�\��	1�k��m�M��s��q%�h��w��K�!h���F�}S���j�y���/n.���[mM6�Fr%�e��9�$�@5G�}w��}���tj���E٥���6<%Ү	ss��O��mk��@OQP��I��v��Sve��b9#��I����r��!�I�+/�O��P]�m|<��Z���R����4���b���?qQ?���b�x4�������W7�/��th�����@^��>*�#(#�t����s���Ӕ����J���fg�b��B�b���0y��Z5kA�z��8ɔ�Z̟֨娎��E�������N�uc����$�*�9i���8S)tk��6c�#g���Yqc�M�v�UHl�0���3va^ݵ�b&=�2� �4e:k�ޢq<���>M��0v�?W�>+�h�����@��:�O�h�ժn�l6�a�f������:�7���G�*�]@L/�oa��z���� �l�n
�D`'��)�O��>?[�5O��H"��6�<_��_J؎|w���u8�٫[#������RP�2n9i�<B=����kߥ���x�	��n�w(Z)�M��:�kպ^���9_Ҙ��tE�0��fmmm��ߊ�� _��/��~�x�%�����~�0>؀��T�8��Kg��3�XW~��s�����*���b��R�-��6<#�ٌ���b���n��L��+5����>o�O��7��>�Ϲ�pV���H�x�uD�m	���F�m�$-Xh�'��L�4[�2��e��

�/�L1{ۋ�.S�j�]?1}1Z�	�d>?�{�P �2�1��S/*�D
-Oe���5n�Bx3��;|I�	��RT���K[G=ƦR�7p�07fOM��[�w�E���.b���A:VY��yHf�Z�a�]�������Z*zܙԒ�2���y�Db$5A;7��l��T4j��ĩ��k^i�}�O.��Y�R�-���v����*����~�;-!|.[ݩVNU�ϻ�=u���"w�)���h#�W����������څ��K��uɦ�&�㉉	�&��.�I�	
��e⊬/Beں]����N��LfՇ�P�"�����5�iW����V�.T�U�9�L%�̝�B�)�t��к��n6-8����'gƥK�q"�-՝4�m������K�{h�����ܻK|L��	-^���k��5KD;�}lJ6�~4�4SRd~��a���He�v���v�r��?�RZ����8�� ������Vp9I��\�e���λ��O�sN�|�#.&}N��XR"�7�.�!�]QzzzvF���������o���F�w�m���U�oK�W5��΋��'�.OΫ����NEY�֜���g�4��/�3�d���A��}�鶃�g�u�v�b���2&��ݡ�,DA�6>����<�����al���-��8�aAZ�l�Le�؉��eS��W����s��܃Uw�/;^-��YWk�ԉ�r��yk6j�U�<�`����F���8�d��S��Xh�Y�� m���~	#O5��\	�*���R�>���*eL��w�W��Fǲ-񊏅}ؐ$h2B�#���Hx�~J!�K�~��,"��u+�[ͪ�;�tω=�/@"l<:Ҙ �����C���b:�Š;��b�Z&=X;�Q�^�p~���[?.U�����L#(S�~;�vu�_+�y�d'�*SJs쑄���Ԙ�_f�He(4 �_���|��B���/6���7�K>Ĕw�|�h_}���T�o�(� I�9�֢��9"A�����W�9���>��>3��;�K��7�I*���0&C���]Vz�;|k}���rA��T�F7��R���Exbӯ|Z�8:==--(�{��С�K�}n�Q��2��+vX�"��f�mn��Z\^���\o;˴Yk�3�~�*)��7�eL�F�7A��U�(�٦_���o5�@���g�ҀT���M/%�\�bR�f#;Q���>���)�Y���VI�tօk3$���BA"�v?[j����0�Ӊ���/=�lx���l�ºa�J(ۏ?i�����R�8O�R�?J�Q����s�~$��˻%���{Me��S��w)«Vrt���h�%�mظ�P��*
����xzzzn�ꦦ$�Վ�m��ԗY܆���j�ew�@���� -�c�mm���]_�NG�x?�s9��3�)87ݕ�(D�"�p���g-�@�M��A@ޝ)D�l�Bx�<{����t8�4�Ԅ�=7��y�^���f�$@�)q��|%)=LW�T܌�r/�ٌ��K8�}��)π�-Ch|�L39.�Y��vǢB2'�Ǘ4,;%�X*�Q}ks����\��!/6eSU�����A7*-�~���U��.�|��ɂ)��\�s�0�ӿ5�B�<�����1^Z^.EM����F�h{0�R��g3k)�^��=t#J� Gd�s���<88�w���������p�~�,���<6�2�)��{�ww��mtCY��WEkHyd�q�͞����mo�/�2A�U��p��ɑP{5!*k.�����P�<ɯ_�'�����Ӳ�j�x�[�p�L�HD��6�19���Ԭ:Ś0\�Y�cR�˳r%KL��""5��,�-���jSՉk���e�P�ԛ�ƅ>�^��@7�ɉ��^bk%�o*���/�c��p�P��+�,����;66�R,����0ҷ�X�J���Ӟ���܌	��Z��mt�ZZX��Q�|X2p�& ���+�ˢiǫA�R��	��x��#�ٰ,�uC��vQ���h'xk�8h,�Tȸ�f8��ɛ˗�)�/hGܨ>��[��B��;uu������R1`Y�T��kG&�o �T�qq<$Ñ�;��H��sh�yA�\�%�1]��*��5�6q{�O�Y���S<f'�[$5,��f���]y��>�Vw9�r�^�iP*�j1��i�W�r�4�	��l-bv\d�����I��񑘩�) ����
鳹m��\���>��ZTrr\͍���H�u��hA^FD�5��qb;8#�����=��ɾ�}ER�<~� �	�O��ގ,	�A9.���K�}���X&<j�X�P*-i	t��5�!<bG���G����t�gS�*����k�׫�o͚¹��6�η��T:�Ȓ�?��hZH��5��ɸ!���8���T44X�z�Ke+Q�w��8�&&�!���-��EJ8���h�'-0��F2Ioa�A���ޟ�tϝ|��~}���x�6��u뒎qOYYY�� �N9OO�]�r"$��옅�F7"��?��2����9s��3[�ң��ᤇ}�ȴ�z�C8R ��N�ث�(#+�[�2��cL mQ^��uP�u�YƱ��1b[��%
g���ާ?�Y؝N�@��q���?����ƮUlOM�`���lؗ��oK���!��u�C����H�R�',�Ht�A"��$?�����PU֭�\9�2��Ω�5K�ѕQ�Z~��'!~��j2<�p�O�[�O��4��a�HA��l�&�;��R������+���HˍS��p_&�")�H���F{�/A��EX"E�|�J�J�H:�N]O3feeG�)o�o����h��l���5�Ru+�m[w�=0<K\+������'N�0��򩴼u`c��-� ��]�e�l�����~�B1�l��4~/I*S)���Sx�zk�5zE=1�B~
�VY`M��*���ߢ��;mu��p���Z.��+
q���[���Eso�_,�8�r{=�9^��M����ҫ�5����������P\���q t]�i��Of�HtځH}���&7!�K����N �;:Cj/�0��>��)ٸ��E/�hǸ��2�/��_}����W*��+d�
����-�*��ƴ9��Ա2O�BPY@B�b��A�8j'%���������湆0n��"�[�K$<|���[��~AQuI���]H�*�q?1�6�W��k�g1�$Sne�3��E������Q�J�O<%b+�!�����ꭍn�oZ��F���Y�������8\u�$����8�2~\�,��@��;��.�Ut3@���_L�]q9�Y][��������\m:�\(Wkt��vm��0h�U�k��[�A���r��r=$�M�'��d����%��;#��<o����N��(�-D'��oW^T����DM��M�P����E�sN�����I<!����\���?�5hU�F�$@��҈�D��<O�D�Fy�<��
k2�R/I[I��9dܓe�܈��Ŭ�݌nZ�^�P�}��&j&��'�³�7�ƽg�Ῡ���V�ɍ�,�?O1�k�V��g�ٝS7����&g�#��t��JL�mw�\�Y�����d�p�B�Û�t�$u8Ol ���i��>����I�Yuכ��g���ی��q���v^�WAW��������/��o�����ȕڦe덬�MLw&�n�ǒ�&7���b�|^�֑{RZ�D�Ē��A�ǥ|�8uP����Ju��v����M���Q�6u}����qWV}�f�����Q�Xc��Ri`�d���d��vN ��'?/@A0�F�}uT���AqN`A3i�ڑ@��@mH����O �j��.�S�N�t[(6#AC��7=���z��xh�V�<�Vl ��'獫��Q�Y�w��D������I����K���90F�������yr�-���}�d��vdФ�E���Z���r����JZ[���6�I��~�4'P�T$�0�8ٓg�b4t���&��[�Wss�c U���v���jk�j^]9P��ۨZy���I
��nX��������]we��߂d"��]
��y:��bō�ƍ*X�;łh�GK6���'�u�� S�� �~3O�rA�CG��F�Lխ%@��zǧt�ɿ���9ӑ�i.�v��x��� 2[�Ȗ�
��۝�}�(I��Z:a
��V����_�z��,OZ��?[[[m��/���xxx���).�oB�xgT2������sxk���:g;��9�>^^j1�ő�΀}4I��a�������QH n�������B@?�n���qN��WE` 8������5cj�No�c�/\�u`t�߳������G�����mF������*�fH�����*�-���2��Vgl/u��C	n��u6k���R~�"�������ުK�~9$�Ή�SƱe�&����a j��QL}�ꚥ���݉��j{Ni�/s��&�8���������������J�C�Kl8,f�_Uڟ�~3���!9o��2Z�}���W�$�Բll���q������-S���txJ��k�5sE&�MoR�Y	��������b����������M���tfp�4��z�3?�K�./�����z�����Iq�1h��ƸLA
-e�ѝ���c7x�纗"1��}5Cfߏ�il��/ t�Y]�EN��=���A�g�ǒ�jp�����ǒJ;rM���P�/�aض�2�b� R�u#,.2��|T!9�n�ڑ�f4���t�v�O��2<����sS��χ��V��3���	��+s�)=&��
��ΠXn%#�H5
���A�-,�����=J[�o�3rznfu9� y���w��9�m,����
 ��w.(��>K֢�j�Rz�]�K�����ѡl�D����4#n=t�G}�
ê��z�ټ�ң濘�Ҏ��t�?�_��4����m-{�HP� �_<<�PHxw�T�_Z��oyeѼ/���n@$G�7�IMMMM--1*�rs�7ϝ��HZ��K�X�Nt�P����n������vySG�0����QNW��x�f�f����eeR��7��>�l4�y5o����_3���g�&����W� ec�#C�{���v-�ގ���%��y�U`!���eVd�K�������ܕ)dr��<�y~�_� BVy�#X�s�p|{�����%8��U:IѢ�������KW�_;d<��m������%M�����2$��M�y;���g�8��E��3s%�R��j��-���*]��]��0�����x��&"�S������U���ȣ��F�6�vU���*�p!�����//Q˥�..�?�:�Rm�l��C#"l��]X���}Y�����]"Hm�w���R��ŀS�S�c�_��a��:�*%��g�����:>.�e%?H6��H� h8�6�-�^a�.�:�L�94I��Q���;b!R厷q?;�t�hė�$�	%�ka���>�f�Bp���S�(`%'f3��x�|;�WQ(�|�w5�v����*�ʙΰ�#XPn�������iF �����vLΎ�w�y2�#'�-x�K&��*jڈt�D'��C��ɭ��6N�5�r
�Yi*@t����Ԡ��UL:��3��<Pc�*M	QU�f�>q@ĺ���$��T�iZ���v
��w UY�b#����?�W'E-%����/�1��z;_�anۏo6�~��]��|�5O���6���ӣ��7��Pi��Z�����Z��g�l|F��h�[(��/E5��Կ��,e��L�si�ˢq��wٟ-NL]nt��^؋o�����6�I�*�#��l)��� 
��1
x�h(o�����d[G��^��&w���JÈ��֍l�w�?��=A�9@p���mO��h7�x��Д���������}�"̽΀g�)�&*U��z�����"�<؆ �%<�D'�&�O���jq�t`l]x�b�S�6��d�������N쓗��?ܣR����!Y���ٜ���v�ϣ��Z�b��Fֲ�nэ�9S=]���EsS<��|�8l�O����^;g5[�.g�/�>���Ɔ>*� ۮ~<�oBܾT�F�1�Q8;�I4_vJJ�Lև��2}��~�݁��D���]��S����Go��f��B����%��.�����!I۷ğ�c+��|a�.ŎCe��_���
�a�
�l�-�X�$u� �f��Σǣ�%-)�,�a<�$��V��̔If�q�����~�i�/���&���۬��;��~aH:�BΔ�4�?׎^i�s� ����퍀H�C�lj���v�cd�&J2�ǟ6�U�tY_�}oTx���S�x�6k�V��P�EfT��э�P 	����P��XEp��j��o�G��4��Wp�z��a�z�-9���zޘ:��s���zcr7���s=o���<�-����$sR=IJ��g�sK�1��I���'$�}E��ڂ==����g4"K��G��WO͕п-�7�`7����`B�T	b�j�ab/�1�ĊБ�d�Z��WJVO,df��1dC�]��j-��yu�`�>���1�oQ��H��n�E��w���U�
�!�h8`�}=�p?dnp�ys��v18*�r����wA�U�>5���Tʿ�i�-!~�Y�+H��d�VH��r9H�w2GԄݺ���I�"#u�%{\m�L������p�ˍ*�y���,�`g��0�����
\��xX�e����:���-mr�<n����q�9���9��	�I��E300�l����� ������f{��Ũ���M�N/@ɻj����UT��$�tڝ�0x'��P
\�:�y�)�F�W3�U��j�-�.އ�L�%�j������>^�T]�d��<����DI�:25�1@&����s4�r��0�L1 �3ݗ����<o^R,Ɠm��E��Y��c��}����=�v��
4�����Kog��c\��N�7�2��'I}���)CT�[y�9-�̸�m`��m���=����GM�؊��p[l�q�*�x�٠Սh�Q7���u��G�;;;A̭�.I(�R��v�p�q|�w��Z.ӣ��
�U�~����]�5$]R�MM�wqجr��8�����+Ȧs��Dp]�,n+�z��<�ov�8uK��P�+��~��X?�+�ZlC穆���Tj��u�G�"ulk˧{T�6ڌ��]<��J�x�׽4K���i�֒��c�@�(L9��o%|^��z��o�e����h�����99�-��!�y���ܒ���7(�btb3�Q/@Dk��U�@�e4��F?����0�Qp�]��k�;��Y	`�(�����wS��_ȩ��e�9HE���΂�����`Õ�V���j6�Bk���8��0��yF�y��.k�����B��q������C��\��8�&{���~f�6��К�- ��pW�@-�+�@�djz�f<��ڨ�����!��Hs����Bh����&�畮ʠ'�ɹL����M�j9��=��:^ry�ˊ�Ju��+ȅ��6�_�D�h`A��3������n���ŻF�t����{��C!��$��cHd�'
��fz��/��ONڮvUDg��ji�QM��gꞞ^�ꮟ��N
��/c��'��U�C��� �mD%f)�1i��)f>']V�H��7�d*��n��2�)��m�/(Y�������ZG�G���?�ű�j�.��c����9�6�Ì�4����s~y<�:}�YpS�
���{��Wr��K������n��{<�'�"W��<U��P��e9�u��F��;!�i����)]A�A	t:����u�;!����*�E�dG≨��D�����~�@��cxn5Yi0���x��z��S���MY�Y�ۓ�gx����j���G�w�N����Ĉ*��ڮ�c
ݞ�9r}y6��r���1!5כθ���X�Yz��=����Rb5K��`�o�;�&�<wBT�I�ۉ.�=�>�:s���:6wn�
�o[���ZP�'������S���򐘧d�x��x1��ћ�XWs��J�ؕ#���C�ehF�����
��ai'2����h��u7=l4w]�(F�!t0LO4t/ ��p ��@���<�c���yq�J��%�uۏ�����W�����9��8�)���Nd4�#��z���f��fz�1&�ѷ���K�Z��\��[N�}�������hH(�J^Mٺ5˼�A��j��.�P�kR��ݻ�
�*w�B�z�̗a�|�&�}s*-z@-� ��M	�eO�ٿ� m��@��x���� ��<C���
@�}�� =�ݏ�#����_{�)��F��lP1c���4�]|����8�g�t5���7뱾��V�W��C����)D ҏQ�j�cU�
Sp�=�����gOq1���X�v�-٭�1zOkk�r��-T�Kg�R^Kn�'&&VX��7>mn��nQ��#��Ĵ���C� ��h��f�͛e��M���8%Wf6O�\����z����C���̝�T��ـMN����ͺS���hHO��щ��r&��^s�>O��ey��[7�����Abt�L��(S�'�	�䦇�6H����b��ieq�Mf��|�a�:���-�Kq�2�<�Vi뉣C Ѳ�J��8�B���!��!�h�����v�vȧ�##rܕF�E��bn�;����3���C,�K� ZI`Z���ҩ]�ylk�R��e�U.z�8�|%�-�~����|��;4��}S�|����I@��G���������4P��_ý�u0������+���� &��Y������%lGGIII3�R��W���R�=��"9��.���0��"��JϞ��8������.�� L��dHN()�J���qy�
L�/��M�Ç[�tڣS�n�[�����ʆ���N��	��b��Ǔ`.N6��*�M~�h@�j�dc�������x$yKJ��,���x�tEM�4������+EK|��s����t�Բ�fE��)��{�(�c[a˴bN�Ν�x���W�28�p���D��A��V��Fi���Nج�o��ڃ���榞��U��۲g��_�u�Q�ʍ���b��bTcUz���2B��8��@SS����2��Ώǎ�G���vX��{���">WY?���b�|]dT��P:�2��o@SY�R,�Og��/*uXmv��e�z
6���yj�̛=='��-�-�+���tV�kԩ3gLy�m"��V�D����t�u�R��(����~K4�ǨϮ�'%sI�R�9#��9Q?��Y:��sC���%�2h�,�>)��c��k;���fG�4V"4���zkZ�����kEMk3�@���9�I��������@o��ɼm�Q�D�}��ǊB{no�.id[2�ux�l1�-2��7B�[��&3��NFڴ���8h  ����R�#A�a��e��aݻ�KY^����;[�gO�:��N٫j0.ޖ|�o`I���EQQQ��GE�Y�����w��:�� v�?���':nL=��Â�����9 �5�#��M#���� ��ڔ�;^��uPB���
��N�p�QikΆ�@x�̯�LRN{A��ojN�+���@j?L�Zf
:#�|�x5[��|9а|	��E���C`������:\9���0�����[��B��=��u��a���;�����{p����Q�}���YU�6p6���&����*�E�q� ��q���k�)��,���2(bڴ��	��dv�9^��;�
U��Wր�4|�}IrP��!�4 ��LB�xY$e0�t!�B�9��紥a��͍&�C/������������`���fM}�����Y�CD���'&�~u6<�����c$v���a�.�+�`Y���~0>���o��j�{���E��NI}3�ߴ�\��Zp7u��H^{!�3ٟi�K>�Ɍ�7��T�t~^1��*.�Z��.�e)}�d�Q���[������x�cu��I�[��
�]OS��m?��t��"��l�K&R��_�����������OL�`Z���VKs����^�$P�~����Z��r�~������{��D��Iܥ�^~-u�,��@���dH���K�:��GS@�v�S5MbH+�%�{�@!2A��Rs,P�8v%�39jCΪ2�O�F;u?%���k�:��B�A��y�#�r�8\��yY�,Jo���\r�1�U��ce������pU{�ȭ7���bb�^�W+��Ol����6s�Tp*E�����T�g����s��F��s��v��PǗ�$��xÓQn�Up�lQ�	9�bc��߂�n�K��.-�.��N�Q�l_
��A�:o�""H��[�_���(�2xv�䳜Y��눁TQ�Qn��)|���<	��'f�\��I��(�':W�C�����(�x��?n"�Jf�R�ǚ�ޞ.@��Ҧ�*=�; O�����<�TGH����ӆ"��9�Rs�Y�8�����e������S�Ԍd������
Hy��T��{:T(9��'x��&�MGSYrl|EfƳ4K[Gl���v��#&�z4~W���MQ��M���/�	��ڒ��5$a�_oW��o�t�]�������=<tƈ ��}�kY	�`��B�V��Nl�e��=�&�w��Qp;%��t�lNtA0��7�'g�Ol3�a9��
:��h'�l-n�4�X��>�wX��>��4�&2�"1��+@ �25/6��;b)�f7U~�5�TO� ���MV+G�P0X������Vr*NJ����ض`�߂k��`�2]=�K߁%�5Rs�۾�
Zgyf1m���_�$�Aw20L\�`M�����1��:ҩ%q�}��I���!�5�2�b���@tW���i�Y��;V����c�Q��M�����0�?8<-/ש�z6��?�]j>���jx��-f�(�%�1ьp�B��Hb�B��Uw=�>�,�~M�ާè��^���g�u��=����m4����)����U��d��sx5��L������n�_qB��1��(���{Zw:�^w��r����]��ʰ8�e�(�|�^�P�o�N���O3�?�7{��V	$/�J��?�|3]�� ��A�/���.�o�#�C��e���F ��I�fn��v/T�^���{~�5#F����a��"z;1�g(RQ������=��������J��Ի,�A�f�3I�Z_N�B4�Y �^X��{�8g鬆�������,́�>U��`y�|1��BlWb�2����_�JO�ppp�I�{}�O0?�^eCYkk��Q��I$�ȹ�uq���ؖW����mO�B0��+_)��� ���kn��(I���\��u5�z��������)��߲K�����29e�7�ƒ�������IVh�9��D��CVj��t�yWR)s���B��x�h���+a�'CM�(3y��-n�|I_�D��h��2aD��1�}��\B�_~�JR�H�	��o;�@��)ՓI��zv֞��D�	h�\�Ş����	��7B{�eXo�"e�-~���1���2Q����+����r��Q`�rb�����~�R��n�61���o(@l�X��$+]UYY6�Z!�fD���|�[S�}k/'5�p�Jf����.�W[N	�ͤ )����h�%��źB��?&�,���!ɦ��_�G�۲��� �էOث����~\uX���
b�Z]��ӭ!J���jR;:������ٿ��VPO�؇si��g��ÑĠ+� Y�)�����"���:h��F8�aT<�8�,Ty�t�[	�"��af4&��Nt������h�'���Ӏ�'�k�L�>y���<���'n���K�����Otk%��H�����*=ߏ3ˉ�&�ѣg��)���` �z�}����Fq��2>�oʏg�Pq�y6Y0f��+����
��U�����V}CvQ��P?��a�B��g�<IA��S��u�P׈��Ѥ�sv
.cq��9�~6�1!�Jh"�T��[�`C!�~���MUzep#m�N�$@RR/�o{~�R2-��$䘈R��8SO��=�%������+"8;�PGG���ZL�� �^Jq�sx*H,���O��4h�E8.��z|���ɇ���]4�6�T}��F�M�!�1�Q6�rl��j�Aj4�gVJ&i}c}��{��Í&�?K�v��;�|�ʕ��9���(8���~7Ő�����Д�/�ǡ4G&%��+RΡ�7N{���c�$���o�& ����|�9�w������G���ٚ�.5\�\����On+L��Ч��0geM�A~2��s��ΌZ��f�x0tS�V�Ǡ%%-V�J ��M?"��&�d&Ӑd �@�V,�ȱD�g,���f{�Im��߆�9X�NݨbR(TB��E;SD�BȔ�?���},7�3������ ��OOi�o��;N )����ZM��:�s.�?�Gۻ�5�5�����@k���^za�ٳ���$�IÇ����w/�<�&S((흝TXXs����̀H��=ݴc�Nz��g�=[��0{"� �/K�ʱ�{ֈ�W��Ռ�{�֌g<A����C��X� [ �Ɔ�v�jzw�bڼu�{�X*p���=��+,5X&1%���E!�
Q�mb�qT(4~ �����V1p���u�n����{��H��z��<Y}/H���E~Vp`�Fy�׆Ba������͖1�7��r���f��x�|Ya�����p�|�������!��e���9V�!3Q�w�� ��!�D����JK������0���h7�k�q1�S��TiPu��"[&�w�U�TH�x� �lnn���'N�H}JJ�W��ܹs7G9}L_�|��/���kjk�[�z���@s�HTI�P`�b�� /�B7�(�>c�Vu2�͘q��1B�q�?���Ћ��־���8G%t,t)xU���#�H��uja���!�ص�}%{O.t��aC�K.�9Φ~��?G��aqbo�'��/?�¶���\w�5��^گ�]�����w�G�>�4�a��+K�b����/��r����t���w�#�<Bm�-��C@BЋ���n�z�Ap��6a���v!��:|͞=�f�s6�))�6}�����whú�l��=<ƎK���'4mک�͡�M��z�ム��RY�R�=7/������{��A��~/��]�R�C%��S�e%�XA���G5�jX�ڻo�_xT����!A�,�������w8���a��'8bO.��@?u�1Ʋ�ߞ� [��}?\�xF8���\V��K^��eF�f4~�@_l�=Z�з:;����~�����s4�C���x��
��چ�Lʵ?<؇�{A��<(��!R"!�}��R�|�(���q�5/E�&��sٵ���K��\�W��< 	 65����:@@z[ EC�xN�hh�(lb�'GjE�|�>�������g[$Nt�ӭD���_��[]M��UT���r��q���.��k����O~�aӆ�W�Z�k����)ד�Zr���NB�SZ,	�sРA�1kօ�>dȐ�#}� p�z��uk_nll�Aq�б��F�IVz�ҏ��pNk�r �}&0~ʣKA�9�94x��ߞ1�4��Y� ����k���� ,\y����1Ut�7��X�\jnn��+VғO>IpI��A@"����6vՇC"?����X�ApJK���~������b��^�_�%��/��u����C�����_R{�!��v��N�:�c
&M���s�nz��7h�ǟ��6HD:q����� ��k6��~�;Z���|\�S</�#�R��UW�$t'�p�N���?��S'�q����o����YK�؇3�<�+[u���g���ǞbϏ��D�ȑ<.h3:� o��o޶�:��Gޓ\x�u9���?�������5�ˡ��a�kii�m[6Qg�!�:`0��XT\��U���F�?(]A�۶m;�ܱ��Q��G`����*4������ ���Z�����g����]�|TRڇT�SgG���i���nQg�w;+�1�QÆ�"�2h�uL���t�����\���dJ���[#�[����{i������.b(B}�ӰaC�����_��y2j�(�� �%��}{���[��1{��8�`�[�,��:��ɖ{���w�w������ѣG���Ǎ�墋._ݛ���׀�?���7o�r��5k���1�w���BW�%f����jY&��q�Zu��Ί���<���]��~�G��'�ڵ/665]*	�W�V\*9;-t|��cws����]�BeA�/���c���++��;�SN9%f��:����:���b����4 �K/��~p�,0��Rظi=���d�G���hm�Z���w�u|X@�׬^M��_�v�A��>��Ӵ#���r�F�0���G*�}k�Q��^p�t���u}�P+=�������xO���FS�N�{&O��GÂ|P���(��!�*��p�i�Q�>e�q�V����o�Yn8+�k��eT�#�w-�>�e��5����2m*�����W8&����g��_x�4�|�,��pԤ���C?B�KqC1�����1������s�.�r��˥��Y�008Frƌ�ŀtC���1w�(��������O>�E�ɞ���nVzN�>�.�{M�0�	���q�nGGծ[O���v5�8@��@7�rM�9���
�+������p�"�����8�Q�y�<.+|�M�i�zZ��G�zU�����(�P��JKKhƌ�4w�����I�?�$�޳��

8��z<�w��4}��+'1EM��]���~�-Z�ruutPaa�:��zޕ��,�z)oO���aCG�س�e�z��iٗK�w�睘�����3w��Ti��n�!��UP4��ԧ�x���o���+1aO��ƍ+/~��;w\�
�NBg�jǌ�u����-�ٱL*-+���UY9�7�s�iB?���D'�5��/455^BG�8,tI�2�K%�آ�p��޹�CpH�U�Z�~Xq�p�(�(���s/������� @@�ٗ��c�њU�E4��`]�A5'���od�5�����?���h@����;���!�KX0C�?������؂�sY�F@6:��8���{��%�u���JT���;�+��r����;�Ĭf�{�3O?�~�Є	�8���{뭷biq���������߱��ݹc/=�ȣ���E*WDX
�V,�xl�蟴Х<�;�~�ӟҴSO�]{���O>��b� tx0F?�я� /�k�Y��}�q� ǌ��믽�&L��J�^�5�����u����-z�v3�g�>�n��z�J���k((,fE>�H�I��<
ôt�Rz��h��|�9�EW\q9��0.[���>X�H�BjW�6m�Jo����܊�i��_�K'��� ��{� ��3�P��䆘��dL������z�1��΢酿,�]����j	w�E�Ǐ�q�>m:�^���z�i�f�2NC6|]q�U��#fB�l�(��\jGu" 
��멬���]u�z�ͼG�w�Z�~UT��"��e%
�������`H(��
C��x����t�*WI��OA�r�
^}x���_��}wN�0��s�\������6����K��c�N���K��Z�B���%Y����R&������������&�c3^���ЋV�^�L���y�֭cBߺuk̥--e���{�v�v�+މ�]�ʍ̝�y��K�x�h���t�7�9��D�okmg��g�cA��0�6������ү��Z2x�AAp?������`�݋�<�k�g�����&�b��nˢ�Bq�1R~��yA�)��
�<vҔ��a1��a���{���
S��Ό�3�{���'p���靷�ee������>�{?}�i,��m�D?�0�\�B���J"�⓼�)�J>'a7:�$c����y?=��S<_��`��4�bF`!H��w�W��'�~���ur�i39J��sѡ(�wl� e�F��{�]z����VP���2�2m���3������"�t��|���x����̈́��;�ؓs��gӍ7��$	m�(E�P9��d�P��TP\L��]M//x�>|1�=�.��\�y��V ZV��.��x�Aڹs� ��kJxb�/�����~���������?>�-z�}2�hc�
�r覛n�
�Ņ%Ը��~���W˾$3�K/��~|���XC=<���'�ߞ
r�(�a%V���^�`��n��z�+�0��C�V@EE`���X��[���g���ϓ%���rj���+~�鎒���$���ϐ����LįTW�ab�(�h6l��7�gN�Jh��Q�ҥ�<�m��Sq��}u�#�9@N������T	=��,�[���3�����g�����ɝ�CF�ڣG�D'��UkV=��NB.7A<�]j�ia:��7B���`+���\s-��A"L&^֥�ȟ�;vp��ώ����4m��t�o�	5S�±<����#x%��3��{�WqzVyy��37�^=�z\�	e���"t�#�E�����q��X�]p�\���ۙ(���C��?b��-eG��e �WU��vvtw1� /�R�-ǎ��}H�7���������jŷl-�����O�4k��J��Q�E�/��GTܧ�q�h�'���o�[{��WVF\p!�����\Z��z��4r�(����h��������a:t�������VT0�����ܹ�����i��m��9sfsu@����[�/>���z;L��t�G{��i�6j��Oe���M7�Hg�6�(��1ٽwmݺ��z`E%��;s������k��o~G]]4lT�vک��5�������t�����;���&�z���P��~4����o�A�è�ˤ>\B���QZ�n���Q�tǝ�����|Z��[z�����iP�@��O~�!���<���y^�?�����N�5�~�	��x�uWӼyWR~>���-��x�f�*ڲi+��"�@̓&Mb;�	�����g"t'�'G�ۄnW,ɡh
�a�Ge�����⹳��jD�I�y뭷�����O��W7�]��'RL�P`9%	���4t��C�b.wzyy���̙�kM��b�脞�jͪ���o�q���	:[=2�CIEcw�m�����-�A&�^~�'}�J���I��X�nc�Z=	�A0�=�g�F�8\Y���a�4u
��'�Ӵ�3Dz[��Js�=����"�f@�(ʁ�̙-,�C�+:b�y�'Xq�BcR�#�Y�*��R��AC�0��^W!,-�h�%L� +�ݟ�?dK*^��hƌ�SU-�� ނKD����D�J-�/���\���(lh7,<��S�p��P������(�����е�^�A�9yܟ斃���oy߹���
li�+�Ϥ����;�O?�O>��.�}!�!�2��y8�{�{v����T�_��xGa���Ǔ�?E�v��8�q�y?����-z��4h��O���yL��::�����f����U���-�3���Ѧ�8���5d�p��Ɏ �6�o����n}-�s-�0q,4�̳�(�%F�>��߇�q($�_O�=�n�+�qֹ��Ӈ���O=I/����+������K��Cݴ���������M�@?��}���sE���������>}��b��0�766�SO?A+V,�\w]~�e���܈����"Z�~#����D0N�3Ȓ����G���X�I�n��ʢ����@rȱFl���
���Eg�:㾉g6�}to�,���K/�Z[[������U}Sc�lt�E�E��j<Ū8&��`EE��g�>�_4��X��'<��^������oi��+��2�X��\ƪ�nŋT�������y��1�������^��i��@����,�?��O���QX�\�2J���q.���S����^�i�~�iz��wغE4�Q����.3����۷s��u{�E�2�]���{ǖ:���	�$�����E]Įl�Ѯ�{�����;c'��e:}�it�]wq�3d$�AJ�xW��"4!��pT��o��[v���=t�\��5~TcL���Ns���C��yt�y��M��BÇ��w��=�{����^~?�������/?���E4�+�	��^x�	���ĶQ0n��r����������C����GƋӳ����s�LQ�q3��2¿��/�>A0$<w(�p��gqqv�#M���5��ѿ��oh���dy�TQٗ��Ẉ����٧K��a/:L�@���0?���r��Կ�`����]���~�i2|Q��'?�x �]�^��^x�/��ە`_�:m"�~�m\=}F��N1_�1��@�X��Zx��gi��tۏn�K.�����
��/$j���-8��y�챑%G-�%�$t<�i�;׿��݃Z�1��.��3�`ɱ�T��i�ߜz�[f�:��+.�k׮ҏ?��nٲ厺�}y���[lE:�}��A��w���򧚶&-tl��3�����/<��`	��(�����r������{= t�KBwZ�	.�^z|�8
5��m���p����X�����^K]r19��M�����gײ( ��cG�w�M'Nf+�k��P��߷��0��+�f�D���8B�]c� �!��h�%ށ��n���#YF������!���r�\��~�q��E�V������Ϡ���g�+��?�g!����Bɀ�="��~�Mn?��+���sV�@�7����"Q���'�3�8���n�8a2���#*��L8�=�˹��AxA.|��_�.\����x|��{[1b�$QQ�_��"}�����=��C��`���GK���ʅ��ۈ�bo{�1�^M?�4���{�i^�!����TD~����|��������Z���-��������*2(��]����+�>�
a��� ����q�    IDAT�(�:e�T�馛i�����p���K?��N:��3���H(�O>G��!u��q��ɓ��m����N;�1����� \k�/�M �p�sJ�5t���'ik����/�������X�{|pVA4J9^��emm�S���U�wn��i�	�nң%���WUј1c���a{jj&�{�%�N�3��-[6b��ݽ{���;wp���.��)�z;��ۙ��J�n�>i�$T�멨(�����'�ĉB�GҎ��sW�]����w�-]j��֯���7qO8��԰(��E �u����VX�N[{��9�	���cy=f$����Ѵi3���D�d�z�V^`��:��@��{>��Q__O,`�Ζ��S���[ �&V��(�鵭uI\�^v{ʂ����̄�VJo���͜��>j4�Cͱ��~uN����=��E���˖s{e�-W-C�DX���4�	�S��u��t�E��{�a쾅������bj=�®~xP�u����ʼ�[8`U��m�Ex|���/^c�/��A����/��Ё�C���e����s���� 9`o��H� ���_����zޮ��V�p� �r�<C<�?xo	�e����c\4�b
v��ƻL�P^���{�Py�B	�����2:�s�ko���)/��ZZ��5����Z��
z�?юm;�k��M�4���4z�81C]�����v�}n3���?�A��x�����X�)�(Z��6(��H}��j=tH(T(�k��y��<>�yL&t��S�9�Ϝ$��e�
R�)��(�9�F��qd�m#F�|��.�����*���W_��u��?��Ս޲m+�#x�d�*띈���S��2�:�L��8�r=zd����AM�GB�G�	O�׮�����?ss�+=�.�l%�߳ಋ2��;��o��fv��Ls|�;�8p��&*�!��,�^v�=��9��AiFW�C�sk�|�LfTز,���
d�e���/ҢE�8�I�1b��s�a�˚�L(�i����\s�8o{`� ����?>B�/f�����{h�i3�PG���ع{�z,�U�f�=j̣��g�}����	X��K9�Kq�:	]�(%
y�PX\A��*"�D����ǌe뻸���W^~�-���-4n\��G�r)^_N��$�BF~8W:�#t���P2?�����������]��^x�Z�ruu���"{���~{�A0����2����\�&�<�J	����I/q���\��覞�N
[]4�j$�v����3Φ���V,_Cx����B.z edQ�%`E�%v�++���n�3g�GyE|��/�K흭p�ׅ�_�`Wy�З0M������n��<�<~5�o�6�߸��en^��6X>.������`AT	D�����w@�U]i����m7��ݦ����@%�NȄ�g&�af���2�3)�R�CB	��C�]�m�]�dY�����>���K�XK��K�{��{���o�o/8w>'�Vo����OxM�����\펵�_Е���=������:�-t}9}�3���c5t�;v����d�}^�2崯͜9=�?/��_}���ٳ�����^7obe�.vy+�I���'�%^2�oB
����e.��cG����� �?hEtw@��._�?{���������rW����lX�Tύ�~ܮLy=��u'�E�K u?����� ��=w�dd� A����e�mjn�H ±w����^C�g�FR�~~��7��瞦}������Ĕ�i_r�%�xB���@`@�+em瀎��l�[��c	8�.���LQ��i������W��*� �q��X,�Ly��ǎ�� �l�@�2e2�XQˋ��Wǖ>,Hd�s�?�g�/���9�+-vE�*�sBb*F3g�f��Q���ڵk9����܆�&
	L2I�U��'��%{��.���!�0	�6l�Dm�M�^/���F� I��&�ؔ��ҷ���8i�4i���O�ъ��s�.��Dۥ���&4�]�w��]�4q���Ⱦ��D��@nD�f��ۣ���w��Lr(�! %+������S��.���F�PUU�W_}�>��n��H��N��Ip)�A���/�����:�_\��c�ax>Zi��5������`�؟:�qcG�5�]Kg�=��@�m������?����+������޿_��o�^E�h�����'�a�KwB��A{�н�AD�A���Ve6P�-x{?�������[�/�_4�?��7�=G>j�ر�|�E_��?Hv�e?����}��_l�?��
���i���_�+^R`��f=n�����Y�ʊ�7o�{\�������C��W�����]�fM.�M�*���ݸ�:��E,c���=�t5�j&���U  K��J�vN��}�t�71��T���s̻��`��28���7���7�SO-b@d�C?�8!�

Ӥ�b�_��;����Ӏ�y��a*[���KIt`�!k���� 9.�ki���71�+8�2�$h�8� �Cye'4��_��F�18x"|��(An���i)���2�n�\�zyX�(O{��؅�Tigq���ӌ3��`ţ��fϞ͞p�����v�"�޸�f@-��/��υ�I���@��t2-8o!�6��˾�u����Ŀu�Ai��������8�ܹs����J�8����PS�4�"nxT2@q�6�.����� I3��h��'}��ETQQA����\�����&L�/\~%�]x�Zښ�Á5����1�4O�S=@����Ρ�_|1��Ş���F: k��Y�u)�gX�8��R6����/��	|
+V����G�,E[ۜ0�I�S�.�뼫��k(��2��24���!i���*�����O�5��Sc�>��;w�OF�-q�n�ڽ{w᫯���}o�Ν%+W�⪃�f��B&��JΆ�Ǥ���\۰9}ѓL��5m��ƶ�����=��X��+W��c����Z�fM�X :�ܦ��77���qd�����\2��%Ap�`��/��E�&{�������K�]9 ��G������odv2�,A�����?�%��U���4����F"�r^Õh?k��m2�q/���.J�a��;�5^�7 =2 �"=���3ġ1&(pY�P�`�δ����P � �?�����z�g��5���U�b��P��\��s�0wlQ�|la�K0g�.A�E����c�g#3U�Ta�Ox��e�����(HѠ~����3�Єɓx��[۸�-I'xa< |dߗ�^I�w�ٵ��KK9�|�YsEP;�AA⸦�Ǚ��Ơ~�兂����=�ILxF�ϔ�I���j���N��O@[T�[�	噳gs]9�A	�s�='�B7�.5Y��7���̳΢&���?<P:���<
�X�0�p���up�W����ߏ�#�_��_$O�<
N�2�j��\����Mva��_&�����V�
�% :<:��^:r�/_0��UG2�O�;o����7��P�\�{�]���e�ۀ���r�R3\�F��= =Z\2�@�4�n�Z��}+W�����u?\�fM }��͎�.�d� �nsc����4}��6�������eM�1nwd��y5��p�?}I�t�PPGX�z�,�P��K�p��d�#���.X�
(�e����x5@	�k��p}�5U�N�:�!��y�� ��J]����f
�>@�X���1��>P^ԋ��C(�J/=<��1�+\̸��ĳ! o��)�� �������O �	po��ŜB9���͛�
<XS8qu 2��<p�P�T�Q���PT�hB�'�&����|�Il�>;�����"�9����&Z�b=��"�x2�c��̍f�Ë�{�90�P@ �%{?FcG��xt-��ڄ^ �/��
-[��i�UH|�	I2�������SOa�?�,��`z �Y���TPTH%eCh��i�PX؛3��9�üc��l`m��f'M�H&M����s��w�3]��o\��8{��:�4 !z�v���;B8X���M�OL�6�G3g��mc�[�l)~�՗����rS]ݾ�P��@�y�2�i�ޒDC �V��<�d�Ht�sY�ђ�A�/��:�=�Oq�5�cV�Z����~����aХ>U���3�BLq��Ͱ���(��Z�8�@�
W56>b���ڰ�X8#;<���A�l_q��
� 	+��Q_�~!t���	T E����˾�ۀ��X�Y�{5�u�Pআ{	�+ƅ�@@� X#�O���z|�.-��B�C0B �s���Q�0P���0�������N�,U��[��s �5�
P����T�q�s �`V0�3�s�?C(3 rX��x'P�%D1I�]<`�7�\Y�8�X��O��� �n���4�ωxn��2l(� �l�qC�Aڲ������2�WT2�Ǎ;�����g>����Ř� �� ��'�/{��|}����*u-����:�����|n<x�Ӝ%�ʪ�mqm ��c���x��B���~jm���?�ɲv<G@��宆���E��rĈ���sYXP���w�=��zƯǏ��S��9]*�J-����;��8�=�������Y]-t'G�X��~�t��%-�{��d��-���@��Ӄ�?��^������ڵkЅ���ݶнf����2>73��T9�u#Ħ��$!�7:��f�7�8怇��1G$v�]j������7��Α����!�%d�� �,@}�w][��w\�dbȘw%�����%���x)���U�U��������ۊ���V��zYl}ڟ^spq�ep����z�=6 ���s�3�"����5�����[;���p5�f���8.���,��ωqI�9#N�s%��♀wG�/ȰW���Q#��b�����/�Ic�G@��y����9OJm<�����ϐϏ���4�	����?Id뇸�	�*�U�$3�b���3�sP�8y=�}��Q�Q�bh�(���{��=j�~�V�q��v�� ������q�6���I�ϖP8�Y3�z����/~uw��Y^$|nCCCy ��$[����7�>EȆe�O���v���<�?tނ9�����s:Y��e+�}������֭+�{t�Rc�Y3)N�7kb
bz����g�Y������8A	�^��1VXP;vl�{ݻ�Q� ��1����F�x57�x�ui����lhn�4�`I�������K���'�@d�i��H��(�( hl۱���ZB�)�nv��Up�J�(���ʀf$��[��t��4��CQ�8�Z���5��c�q�;]j�UQ�w���	
��g
�Pvt����oV��2G�C~��5���:n�
� RThlY�Q�]�����z?�g�uU��1P
�! ���s��(��?������_���"P` �I����cz��s-S��kH�?x�:
���U�	�'�����%���ʌ�kU,t��հaC�%\�}1�5�%%?�6��?�;�1'��w>��w��|�'��t���MMM}�@�� )
��Ho�#&�� ���Yn�b�
�Pn�N�/Y��d�C�-8�?z ����=N��}Ŋe_?�P�ׯ__�88�ٲ�Eī�s��
d�6U �
�iMޛIV�� �WI� .�BI��xV.H5��>���K;��9�� �*q=$�!Kntv����X����P�6v������d5n1i��@d~��v�����Aь�8)K�������g�nX2�U��@��ƉM��X�zd�1�{
b�L���8}�
v��ajkcU�C�����sS����)��;��'��!��������qi�j���-Д���K��Y��?���f�+և�)�(�p��=�x;���u�c�.��;�����kZǮ���{8OJ�T�SB",�|��C�	�,�V.t.xm�7URv�©�C=8�zQ
�l��h��y3�܃��P����JJ������߿�d��������f�:��a�&
!�?�dɒa7n���}��I&��{ �`�߱�}�æ��(��g��u�
D��%��>���1`@�Pl�A��r�n��W.�����'�ׯ/R@g���Q-�1cswR�f[�*<l�p�n�m�y�Y \�&cƌ��|�;4c�i��S/�g�Hac��� Q7&6$�A��3Ğ��k^��agq �Q�0e^C&��~�N>���a�s���ȸ��_�e�)�)����@˂�$j��r�g�?[P; � '���	#\����Sω��e@�\)���

:��ir!�#(.d�{W ���{�]�<�P�L�0���nY �ư5,��pu�C�G���!�R��P���Q��9�f۫�s�y����J���b~�JV��#a q~�C�\嬘$$	����J��^P@b�@�@�]-o�nJ�[�!\Cs28K?fګe����޵ב���B�'���k�B�F�����6x��!<'؛�@xk0xbڴ���<��ퟶTO�R��?�ۘ��˿���|I4�VG%��t���$��J��kt^���\��Q�6f̘xi��_��p�=��i?}�^�֯e�>������nٲ��p#�����������6����2���:�LAd�Zo�0��>LY�ޱ��=�.A4H��A��i�y�9n%�4�� �[�%�(����C�!�
��ȨVkY]�p��q������n1�Gy���ժC�
0��lKW��\��ɊO�\��i�^0
*G���	d���A�3�+��g�}o�
Z_��!���v7֑d���x�P"	E�oU@�͟�]��3_T*ϗ̀�y����n|���6�l��#}�Ho�Z�^�=^@��wf|z��~��"�+m\����(���
iܸ1TZV�I�ȁ�x���w��>l�Ї'O>uͧE[QQ1hÆ�'WWW�S�Cs����jl�U������ �z�8v�A�떯���a�ɓ�X&^6����N����%�p�k���n�K�/������[�l�d�*/_+�\�w�K0Xu�j��b�=I�����u�,b~ ����'L8��������?���cOp=�v�R7\��Fu�#b����{^5gu�B�������$��T��22��J�j��������{Y�^���{ �=�R�����	h��C�;*�N8����^g:.�Ivu]w�<=������!�q���zW{ٙwcqvTH3\V��k��A��p8D����!�\����I0�����%e�2b����jG�)��񫲲�����F�����x�qN*E�Z[[� �[*��U��&��ð]��Kq�{^���'��J~5��������w��u{@_�rٗ��yEEE �5�%'J�3%W��fU/@�jk�^���h'l�qp�#�7%�{޼�t�u�Qoi��mBQ����?=�'�T(c��d_p�yt��7;$1��Q�������	e �����79�� ��'�|��(��,fp��}��1��`5��	�=^n���^ё��lp�k{�O��u��v�����R+��z�Ƒ�od��B�v�s�#}:�}/��]9��� �~71����*wX���gN%����X��p<;p�؟9��Ե���P8\ޫ���eee9r`ͱH۾}{~����V5z��=��ع��榦q�P�d�pޫؼ��vL�c�3İ1�$&C��?MJ�b��o�������ſ�q�9�����̱<� �7�8pwEEE_t�De�4HNZ�[ݙw�U��.�0�DN�4o�}N�ݝ���!� 1�ƍ7^ϵБ��α!��}��R��rZܴg7��h
��u���$� W ԥp�C�h����    IDAT5~G'7( ZR@Ǽ��L���vJ�*�dx�}�Yؙ�Y6@�Zd^�x,�  �(Y�z��]��+�g@G��|�]�cG���!��� =c̪�}F�l7 �����پ�ʼ����Y#U�R0g�X��b^}�U�C�>�<(�G�<�q��bEk�M�i]~adc�~���ۿ������ׯ���,���un�#.NT�w萯`߾�����+�S�k΁���b����DbH<�����#���=��ꝰ���ꔳ�EQ����z鐒��<u�w{ �pV�9���ʕˮ�__��͛���rgm���5�BW��f0��8�Zժu[� �d E���f��+���
���jh��Ķ��z�ꥒ%Ey���}N��e������H^AkO$�	�R3&Y@�=JV*�dF9��Q�� u�A�'��+A�H =�u�G�L���$G
�6H���9�5��Re�#(ME��.�s�l1�N&.��Ժ�.'��'�˯�p���;0�B��Ѐ~��B������({X6�x6%�~>�1��1 �k���h%�4� Bmm�� Q��=m��QR�U(�~7$����o��ho^^��w�>5y����������`^�%�i�I���K%S�{��i��Jۚ��665�hin���\���V���T⃌�LD��]��:�7?�G��sh�:��Qo��M.��S#r��B�o=Y:��׳O����#G6䰄z9�3��}��Wؿ��������DR�P :�`*��.M��7��bq��.J/��v��1vi63b��4��Y��cĈ�ԧwo����m�2�+���vd�G)��ޢ��잿��K9�@���h�
3%l���F��}�wW�b��l̓�@�T�x�l}��;͵h�.�����t���	y[X�ʙ���ޱt=��� j�& ���d��1�{n[Vcv��.-������pNut���^�$؉��q	���RK5��5���:�	�OR�zYY�O�y ��"TP��Bj�H$��Dk8n��í�P(�c�`0�L&}�x<��Қ�����D�ѼT*����E�����J� ��;���	}���}���x�lv�VФ]�'M��o�
��������5��� ��c�u~��%���p�e+�]�P_߶m��W�\�,T�m�QL�L�Dٮs��e���m�*�ҲPr7f]y�4k�,�ڹG��h{u󉃾�oo�������i���o�	�O766%8��lH-!���gΜ�����/]�1�Y��eR|�������P�e��fX~������û�M���r�-5�3�u eZXut�v�3��K,n�Z;�tc�;֏�T��#_��}ϲ�c��J�@�[��2ϒCх���K���j�g��gf�K�N�н�_W�zg��.u{}��,�K�b�:b�����<z�� ��~D�"������zu�R�D��ÑH��e�V��'J���a}ӨF��4\(��ѡFX��9��2D��942�t;i��ퟐI��nX�~�����X��>}޿� �Q��> �@{�A����?�����{*++��8��r�"׆��N���f��u���vm�&�hb�{5��k-*�K��O}��[��N�M˖y���q�9�?���ZQg[H�V)o���k�K/�֙����Ƶ��R�zru�㚨-�����&.�� ��g�x��V��B�d�;�k>x�� нV\�G��$ȳY��@����q�+cR��5X=�����i��mQ���	Φ!wh�㙺t����^YD6H6�f6U���乧=���3)���6("I5@Ǹ���^�
��0�#B�HC$�W�~�ۯ7[� (��HءVR*N�F8d��
!M{�/ ��.�Sݾڹs7g�#YcYgH�bz��7�A�sf�3DJ��:
v:bϏ��l�p)��&OS�����%�͞5���;���Vv�Q�j�=�/]�����wWWW3��cTӑ���\ƙ�2=}��rq6�TY�tcC˾��K��L�����>��k�qs �����C��QC�v��&M�Lx�������NZи�`�ܫW!7d�袋xS��y��,Z�8=�̓, �z0��!XŊ��tҖI�c��N}�2��;Gr�l��l���s��5��BJ�V�:�@�0��Ze\��5��6`��M�V�?�,)��Ù�7OH\�2�����A�}i�.��!��ȓ����^�!�O�ӽϺZv�CO������MA��x��޸�Iqb8�e�m@7�r�@A]*�J�I&��QV�p�����
X��B�����` D�p9�L�
`�
�8�(�P��\5������
��ErNI�B#�l��xp1���3��d��}���)S&��Q�%���y��ΰa���ly�
$?K��, ���� A���n��Gg����5nP��4�,�R]s�5t��\r���ڝ�Î�64M���+4�QN����O�^�-��Eh�
�����R��kI2��ө��̜�'�x
��=��{�QZ���L��øæ-�I�u��u�
[�G3��|� =0�6[@�pdXXl�&3��
j�����e<����D�H/��t��'���˘�f`S�L�	R����gNt/@�+t tGv@g����H_@�������e�^�a��mP�dU�O��r&�c�{�p&�p�Ė;�:U-E��>aY C�eF<f,�˃�6sX��?�.�qpQȝ�����H$�rG\�J����fϦ$��r� ��ԩS�q�,.��ܹg|g����}�H��g�{G�?�;T���Ʊ�a�����zgV�*ꢃ���@E�υ,��9( ��mڴ��������͇�vh�h}�d8�%�K�y�SIZ�����g����\��s'<��Дe��b��p�B���{�YN�mV �����Ҳ5�P��c���z=��@@�cT�s*#^6���q��wX����ZRO����� `��:�}���E"] %� ���3�K��T�m�gn������:0ޙ���4k?�vϞ���.�;�q�>� �+Y׾��>]6��>�ך�סZ�
�@����9�CiI-�WJ߄B�oZB��RX�v-8�� &o�*8>��/��gn�r|��B���U!�<쀹΋ې�L�qֽ]���/|�
�cƌI��xb��9�<���O	&z.cf�3 �K�:��x_MM�@X�p��u�ڋ����ن��6�j�ڬD�c�qC�������r<Lv�1'�����Ud��t�It�W��'��
 �����/���=x�����n���鋷�D��z*������ <����a���p]x �����Z��2�%�n�ҕr������� �o���v�[`w�n���̅R�����g<�i�q��ʛ���k�1�#ϸw'y1�M�Q�H[�6���'ۖ�B-渔/�xd{n]3�ez.��}�ñн<1J��u{N��٠̠k=?���3ʂ[���`�u}�Z�Ա��9�k߸�U!`���?#��(���B��?ݛJB����~���X������ͲL׽�c�ӦM���F�_c�9���@�
����@_��Ɔk�k��A��i�Z��	�q�?�g��~��ERj�q,6~�2���Qچ^��=�&A���^~�%t��S)�ۘ�����.�?<�iJ�uk%=���r�2>�M�->/f@w�r,�,C����psu���|g�[I��z��u8
�s��s�'�՚����aՂKոV�`a+j�g�99��X�f@k{�[��=U�g1����9skb��n$w�@.���P;[� �{���9�&�f{^m0�����ٚT��p��$�ʣ�2E���	�t�c���z�vi��^g}��>r�y͚*��Ks�GM�S�W7�gSxm%���Q�PѹB��#�g��i����OΝ{�7{ ��vWg����r�ʋ�6�����Dc超�֜;��\�[���i�6Kʟr�����p4l��a��{��p�Ý��X�j9���k�|�Jjm�Z�d���w�N�5z�tKq���Ï9���j+NL�q���Z�ߍ��tg�:Y]	8{��i�vR�[IP�ө��,$�xpMt7N�~�U��>��}�~��#yk�.u:6G@�K@���C���y1��
D7@0s;�T�����s0C��H�������Ӑ����`�0�v�� j����Ε�3��uދ�Nz���X^���^�f,�\� @�\��j���]��#S�S`��𵗼Al���_����<z���8cX�J�����@^c�^���~i���y��|��l쾮 ���c;�@�����jjjʼ =W��msz.^�X,d����o[��Z�K�mH��馛��`��xЄ�?>O�ׯ���=@�zr?M�6����jvѣ�����o�ZE�<���[�[�Z�`����mM�S��\@ݭ��s�t����h3���\crW����h����'r$�_o�t$���!�� ���� t������um�V���ɓ�}!	MǨ<w���=
5߰�8yR������tP��fu���`�������<2�Ė��f�\-W����������Z����'�ˢ�0t��@��%���4ֻ��1�E����3�+J��Z�u2�8/wxҙ�j�����.6rtwv�k?�)4f�(4�������Fi阽�sݞc�~�=�����w����555��p�D0��Enw$�6-�Y�n���]��d/��	��jt��{�/2g���j�:u��	t`w���i�^��%��23ɢ��V��>w>؏Z[��y{{�V�\I=�+n�
Y h����$��Ր���ɝ��ԣ�,�\�~��}.�Ұ������$����>ر���\ �Z��)�L���b��q!�ϗ�4���P��Zz\�es[X���@�s���-Q9F�xG�D�iPX�.��X�6���=�	S//c��cr�O��d~�ٔ����ኤ�q���v��+6���%'��a)����l���Y�xN����a?b���=���_�Z�[<!�i0�T&U��ȷ���+2 k$�IR]f�M�NWk䮞�=W�En��l]I~(�C���1#i��A�.X0��=���L�ϻ=��Z�f~��������N�s�H���`�F/�q����۸=��e��T�W^u�w�y��f��C)Hg���c��� ر�fϞ�}�ъd--�,6n���3˖��!%�lE�~NN	�P<jl�Y7�v��lI��f�y)^�zY�:&�g �)���w$B0 �|.�ArQ0� 5؋��P$�?���k�k;�"'�އ�P��5���/N�R��rݿ�L�ӂA��1��okk��#��|\�`�a�����'|ܱ��u1N�Y�>is�s���W!�[�=�0��D�ЎR"�k,e�<�D�#�T���� �/�3e@)J8���fJ%�V�(_ϣ=���$s��0��~͒��՞յ�uy�������n_�5fٓYJD�A!JM���=���gN��$��Ԇ��ً��������L(M���L�riB>��7ػ�ξ4S`��q,r�p�`Ń�}�qh#;���X����<c������������j���Y�]����x�&v�p �;6,l��������/�u0)��׭[�� X�2ǵ�D��ʗ^z1'��*�M]XX���=Ɋ (�Y0��VtcW.�\���㵚�}߱�]�l�>mɦ�ڳK�\�D���@_���GQ8���'���>�|q,~�x��F�?������  �� �
�9"|�c�@����D���1N~�9W�XN�����33X�i7}	���(�s&R����w�	'���E������B�E+N�Sk{���;
��ǹq��H���&V. �L��1���wO+B�h��k�2̆E��Ѷ` �AI�m���'��+�k��2�m���s3��:�E��y����*��,;t �'Y��o{�ҟ��������wu�%/Ͼ#�g��zX�ş���cƞ����ʢ4���iӧ�������?��=1�.�����}�ڵg�������� t��i��.��E�ζ1����v�����j�8��v��&hȐ!t�wp,<����q�=���f�P��zK��;��|�TVVB��QS�!�o��=�ȯ����"�B����͜U�, ��m!��{%���<�s쾆�
5��B�!��%9�|������b%|��e[�I}?�b���SC��.�c>�X�����C���k�ѳO?M5UլD����u�$��X��n��:�������E����sm2�R��%�
(`�ji����6�1��Մ�F�JF_�p���.\��x���裏?���f*ȋP*��{������
g H��=Z���u���J1��������j��m%X�z�:*����$��K��
o���-N�A< ��9�t��.�:��Ӏ^RR���z��9\w}�n������w౪ʪ�>��C�u�y��rݨ�j���P��e�������/��N9�*�Ջ�f7�裏X0K��l@��������3g��@G��s����ÏآL%���)ٞf��Ǳx�Fv��t�n�&ےq+��;�o#�y;S��fE���l�s�9����/Ҙ1c�-�@P,i���(J)�_���&���$� �x�d&�`�$�\���%�X�uu���矧���'�ۻ�]��ΣmҨC��b�g�}6}��`+�-��	�)0���>X�胦�ƣD" hY'�,�Bɣ*.�4̀k��J�?H!�V	̀ CE�%o/�G}�6�_O��$�Q �$eBs�'M�Z�M�c+j]�����{]t:6�uu��x����]+��m@w[�����al�#����Wϣ\���Tx�u+2�yO�$��u���6'�f :\�O͟?�=z.;����}���g�޻籪�� BX�p[�����i�ڠ٬�6(ڀ�ĭ}>v����r�9�"��C�g�'�䣱��[.^��,��f�,�����_��_{�
[]L�1���u�����s�ȹ(D^s���kv�@�;OŤ
.k@A���[��/���I"�1����o���#vxO�Nt�*����5�P"cP�e��~)��&�{�	�+����L}q�P��C<@�5�9f�	u��X�&Y	! $9�p����� k9�O$hS�F��V��v�a�Rr#~.I���++H�K$8w�]�m�o�q���7�F�M}� 0�ߑj?��XK>� ��^-9%(�.Vd�[4����I�� �Ն��r��lx�k5����C�����[�q�`������ՖW��Lxֲ�5o�3V��|W�G���]�Е��.O-iY�=�~8k�X��}��ug��������`R[�|��YL���&�>ƽx�Z�]�׭4���Nb������r�&A�5_�,�AP3��͛G.d��� ���U+�g��{,j�._�y���G�&����s�7��l�!|�(��e�uc�=���s��_��_i���Η�q�]�ⰰ��\A��jh<H���^}zS��"N����Iq�����G�z$��)� µ�����s�o.Jg�}:����	jhl�ŋ�o~�+)!��:��HX����e�K_�"��.����R<����v�ko�F�7ld%��$���4�w@���@����@�^n����ް�qm���Vo��i�t�YgS<�b=���)�@=�0�^�R2�y]&�Ǆ7b��kG�"����)}�k�{�Y.��uLgc��`�PN�f;����wTpӍ`�����m����ʅ=.���)���¦�8����#X���+��W�[7�n���+���W�XqX��m��@�usd���5��vM/g�70�1ܞ���=%�U@b��y�TZ:��|Μ9�"��5��Ҵ7�x�>��=Љ���~�vG\��    IDAT��MM�Z��	;��3m�K�x	s���%lܫ4k�t>�&��D��~�k4y�d��a�"+��k�������;�.���+(��p�b�����Ps3���2��#S�^}�\��(az[ǩ�������2���4��9t�s�;��D�g_����E��-	�9�"�cs�\"�Xԟ��"�喛�s�R:���֮_G�>YJ��w�b:�c�5��f��.�vh�z<�Q�x. �������ׄ�9������o��>}�͔G�aڰ��x�AZ��Ǽ��r���]��Ҡ�н$R.
�������"n����>EW
HW�t�$	�e	����nѹ�w%�^�*;޲����<�3�uzͅ�l����Z�T���Ї�JKK�r�V�����t�'����r��Y�v�z���j�'�|rT�~8z6����D���B�$7��.U� � MV�2%,���R��zkk3����_^�3���;�g�n�hTjP��Qj���pҖ�E�i�))ݏ[�sg���~?��u�nW��
����U`��m�i�vM �4i]s�ul����;\<��i �P�0�`׻��k�����o�AMMMn�?$�I=����ӻ�_ӡ��B~*,�g�� 	Лo�I��!�r�it��W�7��n8B�����Gz������V���&�,���nΟ?����op�C-�liWWm�_~��,y�Kg�:����
�ݫ��3P�����56����0��ð{�>ji�����`��B#F���-��ŗ^���C��+���&S^^�����Ѫ���h�b�R��P.�mxc�N{P�0�E)���\�?]C)���Zsـ���θ<�p�qo�'�����r�X	� L�M�R�3�������LR ��Ї�JK��Z���o�ԡ�����n�ׯ>}���O�TW���ʕ�Y8'�ݍ������^^������\��)*Ԫ��vO�o�CE[Աc�r���	$[�+�����$�T�Ii&��hΎrJ��\$]������B��~f� ݜDځJ�m� �4��%(��l��.q�L_��P�0Ǩ�f�,�	���$�w�ܹt�7��]���o��֮]�Jт���9si��ZZ��[�h[��x���uC�9�Rp����*/����4j�h�9s&{��y�BB��n�����z�oj����=��I�Ǣ����W�
����;w.}���ٍ� QU�z�_���o�?���s�bue�x��h��QTPPHԳ0b�VB���i����~�f�^UKm��5�6t0M?i*�/N�=�(��ۇn���4��12N�L���|�Z����i[���'	Ғd�c�v� �!�^��v${P׍}�l�`����F�h���^Ӷ��cSW�g���=��IGEm����-9�j��5'�����Eq�z>�P`�g���<���#P�&bT\<��L�@O���==��=�~$�(���}�ڵ��ܽcQUU�X�oڀ�5�^��Y�I����q8���P
��n��������$��`s�T߼y��<\��(�wHd�gФ�8����-foH���%�:�LA���z$��K��s�o��f�fED��k(ٙ:��,��`�C�q#��q�P���}�ݜ_ѷO/���?Og̜� ��%K�������_N�Ǐ"�:a	!�&(�C�+��Jo,~�sp-� ��?��!���v�4ׁ��PS[��|�9zz�m�K�8�4��(a�+�}���rg0��iǞ:��#�П_}�"� �=�l�1�4Z���[��?�����L&L�>E�8�nxt�
E򩡡��W�Һu�h��-�{�n*)H�f�Fu{�g�����r������ӲU�����-N<&�I {�P���cY���Lr�,7c�te���
����s��Sg2�����%8��v.��LA�AY�a�=���鞰���팽�����#te+d�����L�b�@?�p������nݺ�;w�>����x ��U�l�#�P�{[����JX9�����;����#���ϣ믿�F����۷�Ig�9�Zuԙ3"�f�Y���f�J��촏
��]ݓ֞*(��{$IX*����l��ʊ��0I�^���� �,x��_��W������]w�����}�O��}鑽 ��+غ�U�G��h�8�x1�&�z��v;��x1����v���j�*z�տ����o}�-�D4A�H�œ�آ'��I��l�Fh0"��|X�=<���;���%{��a?M�8��;n'@"k��i'11ь�f1����H�cw+�;Hp��no#ڶu;��={w��'ӡ���oI�y�<myl�S D+���=��G�*6S�y�����͎i�k�+@�j-���Z�� L�'��m1�*�ʮ ]���˝y���V@���e/�-����޼滫{̐]�������%���J�Y�4��(++{��s��N��=�Uy�����v�ک;jj����}��+�m�fz�4G�Ԇj3�B7d0Ǎ:�fΞIӦM��`U�"D��`&�A-(I,9�%`���b�r�k���67[����(Y������id׽q��u��nj�m닁�($ t�3 ���t+�����7��ng�-[���~�3.i����KJ	9��g�9 ���
g� �ľĘ�1��#�`�̳���}{���_��܏�߾�=�e��`^>hl��=���yr��b�ƹ�-�L�w���!�}���sR���v���;铥�ϗ�ѣ��ݟ��/<�B�,)�ӑ��&�H�b����煨�1A/���^��&MO�`�|�^*--�����hܸ���P(�Oɔ�>^��-���6��+X�)I�E+��T���R�e�!�������7�W�K��c���{%���d�`u�amy�O{?tf��ߵ�����{-�/����<]����,� ��,S }��I���Լyg�K�;���L��7n�8�f{�S[�n� ��|-���~8B������ �9�Ů$*p4F��1��/I�
(	Ѡ�QI�ǤRƵn�m/-�v
��&6��n
��;18��&��w3C�FFÇ���#
�j�kl\ϧ|�:gna����x��b� t�X��SN9�n��v�/�:*~�0�N�<��y��QN�kok���:�.����kz�؃� �{���+�Q"�`@�^�AQ�~�I�����_���,�J$��!�k8HO=�=��S�C���xw$b�+_�
��Q��Z �C?L��z����I'N�cׯ]�
��W]�I��PE�Q�C�z
��1��1f&�a�!�ݻ�O������#������_^�p8D��k4}��\!w?�����rz�ᇨz��%b�>U@�3��4g8æ��s2��P.B�+��>�Z6���yg�߶���,��,h�e�9Â5<�ů�ۙ\�q���"����8 w��r�P~��p�՜E�>� �ؐ!C͝{�w���zڧ�	��1��7l�0�zk�S[�n�@_�f�Q��y.�$5{3�+��e�}�����T�]'(�����88�!�ؕm��8��G�n�%�5�v��Tz�۝� ������X7wv�˱�]�I4�c�ʡn+
��t�*P�;� �� .t �9g2S��iK�.r����IeN?��lG�v���t���駟�o^�@�P����A$����&' @�����Qc�p|p��\7~�.c����RD�$���K����S[{+[�<g	�;ԡ��Ib�H��;{[R>ڽ� =��?��x�f�<��M�B��[�n�^���\��@�~�1O7�ATބK@��"�����_~�**6��'�fN��մq�f��1g�}aj��(�WHKW��Gy�j�+)��G�a�Z���7��q��x��� f�t?s���.u/�s�����wfa��d�y��+@WP�b��X7P�QmasQx�"�z^
��v.���#@����i΂<X�#F�:䱳�:�����"C{�9v3��}˖���l�zj˖�����΀��XT��Dۛz<%�;ؽi � �(~.]rXԸ�d��b� r�LW���Ń�nT�K�A�mU�5�xg���$��c�8!k^;^a|OW�����Q+���Z�����c�u $.q� ��u�]������-���?�)�y�8�T���>�����Ǝg��nVD `~:����Υb @$��9��l�ƍ,�/��Rt�o������ͯ���g΢oo����x��-�c`��k�s�Ա��PK+������sOӴi�h���f�jj>t���������OcF���������9 hߊRFP��R�ݾ�k�Q�����Y�x���9`ƬY�L��B#������SU�V�c.0~t���z����6�[ڶB�H[�n�N��"���*���v�{Y�]y�WT��g��G��lvY�}M|����̵�P(�e����f���ýߣt�rW�; }ذa��3g�� ��>��?��zEE�ĭ۶<Y��b
 }�����B��g���V��a��  k���H"aJ���3 M6�D�@�<����R�h��ݭ�M1���W2U�Ѵ��$5�jq'�qc����ٺV_��,�� W�h*�rx�1Lh���t���Q��W]u::N��|���t�?g���SN�x���l��/��R<x�S.�4�+Xz$��-*]��[Y���u��<��5�������������S4��W�x�y�!ڻw/��O��iij����]�����oI��X��goW3�ڷ_�^���ښ�qCGp� {Qa���Q�'�*��<[��E�#���� �����5k��/�)S�3H��M�m1q�?� mٸ��vt$
*�+5�V��������K��sU^ʁ�v��;��Uj�&i�c���� �����լi��#��^/[A�=�����{n;�_/����U�R@W}��ڇ��ٳ���СC����{�;63�Y �	[+�<YYY9��wߥ��7��3/�,��;,�NhI�f*m����4�& �3��/�X�(9b��R�����]6�qA4p�j�qIc����=��.@ J X�Ѐ��pw����!��pi��԰�i�Z'�_�F���#�V,ƣ�:q.x�����g-��$s�s֠̏yN
�z\,c����nb����h��J��޻i͚5t�YgrM��];9����-K����[ρۚr2\��b���߳o�|L�J\.��AIZD�S~�#�OЛ�C��}[�!�隆9����7;��-��ϗ��p��UV���>C��|�ƏK'�t"%�Qni
��I�=jg�k�4<3V � �DKs+3��>�n�GꙔf˶m4�t(�1��飥�����ʊ���9}����*�E^�Z�`Y袈�<A�|�����i%2�3�E�dF^�n�_���m����� ��2���xZd�nPvָQ~�M[q�s�l�s�U������e�LW���f���=��@��8)6��C:lH��ѣ~;{����X�G�,G����WUUM�+Q����͑X�Kpٔe~�t{�+���%�X8�9j��ʀeW-j���ֺ�[)!��a(�gQ�_��a�A(k�R;�B����,U��9�����+%5�c��T˜i}>vS���2B#��bQ��.�l�L����1r�yJ<�ه�r :�����G��e^��q۾={iƌ���lpO�^�@E�
�uzW�L�9�/,�lx�4AY�|%���W_�1ud��~Jô��w螻��C@,�'ƕ��� �]v}��[�э��!ڵ{/=���/���Iq�L�N����u z������?�G����0�pDڢ">��o��¿c��z�GTUUE�**�s���&L�,nt��B��G��B���r.r:L�<%k ���!�"ə*��HW�K׏Ug{�>Wg.w���{6�uf�}/+���q��z~1�)��^��{3����4]͟�y6e�k��θL��s�����&�),��Ҁ>l��( }֬y=.�c0�y���o��
b�iK�,a@�š�?еy���,+�7�N��!La��Ÿ�(&
�NV�`"�<>��&����h�-t�@2�@�@�(nj��a��84�&��h�oX�L
+����}S	>��W7�S�펧A �YQ���՝�4b�de�B���I����y$V�; ��e�x���.�a�V��Y��J�{0�7��cO;�4�~�[ 7��q��p� @��`�ԥW/�,��H>�I�:�u~����O�P�9���.��s7���ً�C<2!�V���F7X���'џ_y���)����Sq�@n*kk�H(�=�yE�Y�<`��)�-!���Y� t��6���ġ���ߵg/{�O�ĭz�YA�O����|���TP*#�֤X�Iz��37,@��m�t?o/��R�87H������}])�,r=�~�Ɂ餤�L�����b���Y�6�b�R�@پ�=~]{�|�o{�99W�̞So"��n��j�B@�	�#G�~�3����0���� ���m��[���Z�6�q�Z�1�7�
�I0��gS�ܽ�9�#�ϵX��9^6�����6%��+,�%��K����s�sD��@�s�0��d#�
���a

�>��U�eu�Pp-�ҥQ��c�'�(	�Ϗ�&��u�dLyj<V��}~еn�kÙXF�&�� ����^C���w:�A�Ú��/~�LoȺ<x0�3��k�r�,V���5�����N�XxMU%[�p���*v��p�pׯ�&�w?���hɻ�ӽw��T�ܘ%�c�;z�� ��_t�Ŝ��!�Lp<��~��G�w���ae4|�B� 0��"o>�����B��!�A�~�y�H��X�JK�`xN�` ���n��ٷ�hނ�4e�4v��#��ӊ��}�-��k��u��gr;ܠn[�6����^�z����c�J���~w�н���m_�sUƳ��*#�Oԫe�|f3�y)��ݞ[�Y���I���Θ+ps�j�СWr����h���Q�F=z���gO�ڱD����� ����OVUUN�+�i�]�.E'k�r�g��݋3����(wR�|Z��!��Z]�c��	20Ú�U�N���z�>}�2COk|�{�+�����`�!V �⎍p�,tXg 4n�1�8� ��Qڻg�ܵ��By�z>�������� �����s (`aT�Om��T�7g�s}����#ݶ~�d*Ka�8<�/E�S�[� �H�ǎ�$9�9�V vb�����Ā��8�.�c���&�sd���O���Y�w�J��	���� ~��7΁�\z�e|^�@H�����t��w�sAH1y$Ǳ�6���٣b��E�l%Xќ��{+���C�(?����I�@�F�E%�Je����CQث���#V^���Z[�ػ��s�����AMu-{bI&Rt��4s�lS5���!��z�!�ܺ�B�C�:�bc�\�n]�_� 붬� ��+�%�{(W����^�,u��-h{o�{
¶B�KI���<�w'��(��X�c�}��Ǌk�Lzzu��BᄿL>�#��ߔ��&f~�!ۼ,t�raڴ��G�������G��
��q�	@߾�zQUU�4dۀ�ؕ�ԻG:�vܘ7��1����p���7⮩�D��4q"@ �2,vo�b�� �6�: �����rbS�~}(��5j��ɾ$57�R8�.bx�"mjif��ǹ0�6�~�G0hH�µ1t�B���C�Rss+�~�ӧw#c`lm�-[7ѻ�.����E�cБ<����c�l��+� :ƃ���RG�7��A�s�K�e~�u�`�E�	�Ʋe[<^	Q ʸ��O���}�0��*�c�9.�de����a��p�M�,X��[� t�',s&�1.k�Dp�#�K.��n��-FQJ��������.Z��8���Ӈ¡ +r��7�xi����Ќ��%�iTV    IDAT0��UۡV�X���������^(8�M�e��_x>�=�P^>���R��/E۫�(��辀̝ㆵ�e�z4
�>;�lo�4�@���}ܙ��ws���۔M���:W�t�3W �A־֖Z�jxؠ���=�9͖Yo+�<�c�g�	q|^(� �cf�x_ॹ;�oȣ��xn��r��5�ЏP��{�Ы+&�Vmg�; u�j�w@gNmĬc�����{�8o�J�xK{'d�c؅}��dښ4ʰX��88��4-�� ��%Dwjoo�'�Mp� Γ!�`�ŢB����Baǻ%D�
���%� ��/1t�q�s��㏳' �%�C���k*Wr�#�M�C�j��h��&��c��)@G�J��O��?��P�}�I'r��mq���}�p`.}�� �U��s�����yKmذ��XA!{�Woe���t��0������;D�<;�N��s#̂��q�XBxV�^G��/-[�1�*ʣ�S���gҸ�c��������*�dB(�}�~%ڄ� ��E�|5<� ���ߖ|�c��/b.w :�C�?a@��o��k�B���)kG��$zd��.�l2��g��Z�-�l1l=�hsv�
�L9���^@��w�����fυ����DR��wC��4����y)I�}_*Lh�0H�B\ފ��5ʖ�1T4�]A�#�5
��;z,��D�#�z�����㫪w<YU]5M'й�7;����������p֢ۅٍ�ŝ�.�w��K��1:~�8���.�9�'��U�f�'�LlH�k������q�?7ԸHQ�L2�`��7�
)�p�2� ����f&Y�n!f��1V��޳g������K�R���]�
��.����ρ���9��N�B�m��k�R�F�ôa�&��C�@:��'O79΄PF�>}�� ��a)�
����1>($��غ��Р��n��m&[>J(=�z㭷��_�I���*L!����q���������[��A��M+����w�[��߳f�J]�y1t�p�G"�U�ݻ���}`�u��p�8$0Fc��{�N�za^�Mz���W���<K�B$H���>�x��w��];j������6s��Xm��n���T1��������k[���]7����
��$��L֮(��t֝ȏl���}����vy��煇�KF�x�,w�W�XI��{T�UDH;caUDB��-�'B��7��v�z�V�8[��оq�Y�8��EY��"�b*%���a�/z?�6}
�3��qƌ���r?D>ʯ| �j|Uu��55'B`�ZY�nd�������ok���wm�^i�$ŉ]68��x"E'�����Є���9��lk����X��%�ɂ8�g�-k�p���%e�ODc�A�������R�ܧO/v��ǹZ�Na��ybå�'.s;Fh ������ku�vN�B�W(6�H��Q��(��_i��w�S;�NL�/�Ii�_=�p�\8L+V�`.wX�Æ�6�S�N�{���{)87Cqx�A�h�j5�������o��!� �~���t뭷J�Z��| U	G�wޥ{ﺛ����
:��K�@�&d� l@���^�n,]���/�zw�y'+#`����/\B�J�52���^�_���U���l���>����X��~�/^L�-m��/}�.��
È�F�H-]^N�>����<��V4��І���-HSm^^�j�ָ�V:�ַ�^�u�t�X3��HI&�?6E1�R�#%�� �����/���t �W4���c�VO���񧩝���X��9 ��IA׋ǣ|�'|��4;�xQ�[E9��\�Ov�ǥ���	_�F�%�����G~�p[�b��(s�W ��k��i��&�V���jv���]�{�^**ȧT����'��S@:th|̘��9s�eec{�܏���{��+++O��^@?	Bo����ϑX�k~rt[۷�tg��f����J�j�"x�4q�D��~@�&M"H�����ò�L�f.qlqta�b�H)_��Ș6��M �l���*=+~"|��,8�7�u�,,��u��8��]�h��Ǹ����c׮����Q]�u���Pu{�3�U@��q;,t�׬z�}��P( �p��p��p@�ý�;�	���k�Bڣ.w���w����֯_�qzt^�#)�k�AjO�h�_��}w��:[2g�
�S~Q>���z�W���x���9)mͪ�<�9g�f���%��X�W/ɭ(�˷&�:&^�F�*8��%	��l~�l)����E���9j�a���^[S-%J��J2ǽX�DqS��t-7���ۂu[�{�q�i�6M��.��N|�CW���\P�<�����;�%��b�ki#���]X[�e�}*�b�"�{PCp�V@�DI(������-��5���e����(;"Gd/车�����Ro���F�P��T�P�Qy�"0L	_�44Se�Z�|5-��{�ذ��	(�(�lg��'�#�d��4t����1c�9����#D���g�kk߾���w�y��6\������xY��NW��)C���3`n3a��R�m���������谪qLyy9�}���K�1׀ =��5��
�8��YY��<(0��^K�p��8E7�� � B �o��UP��e�6�ӧ/��ҥ˹9��j�Z�H�_6դ�i!dϱ����=g`��+��8��=���.��qvx�~}�0ܷ�d�/��a	 ��j��|�lp)��!? ��Qvł��I�{��ձŉ"t<G(���C���e�9�{�|�jQ�V��=M�4�Y�
�"���|���d��|Č� �5���~�2����ϰ�����"��܋�p��C>?-y�#z�_SMU5`us:B7��t��Fq��s2H�̇�Rk?o�ݠ���e+�����v!�[\�J�����FǕn���k�׮��q3Λ>�|3sJM���l��{eo�y6�e@�*<HV�����p���K)��/�.�MԄr�\(��ׅY8y.�3�u\���G# IoZ���Z�kB(���"�����Q��V�^G|�%ڸ~�[)LP0��_���Y�ӧ ��G��ݬY3��q�w�J���n�UUU�k���v�vt�W�P�� ~����[�q#N�U�	��a�#ɪ5��������TYY� :6�$�IV��0���f����z]uUۛ����9gӛ�&���u���d���A
ܷ��%�1�㏗rD.p���p���Iq.#"M(��r��Z� Y�H����R������X �����\n�j����<>F=.�]-,x4F���@� ��μ &�;���[o����N�rG����c xY1�%Y���_�l��V��ae:�=h���s !��<3n]g ��s!!
���b`5���s��,{]�i�֩�������ÏPնJ
�(� ~n�<~�/�.lzr,�d�)w�-��B6�C
�
��@ma����	=��8��a�KNCqi. 9�ɽ�rp�ɴb�
FG���e{����ʠH�Xq�΁�p}��_gO]��(0^"$%b�aޠ\C.���P,uIb�u�|]���VL찇�93��P�K�Qii��҆��ʧV�F��v�^��_����Z�%Z(��R8�f�0��Z�1cF=6s����c�]���z����o������ ��j6����6ÒΡ��)��
 ��72Ώ.j�i�X2��z��H�x�?��?�s�Nas3�
��Nh���S�=�؅A�Ꝭ�(�X9:F��
vz=�I���Zڈ��@���s{[�>��c�
�:Ѳ5�{��;#a��1^�����[�_l�e�����?�23��i�X��ŮB$>�P(�i0����U�1�:�pI�r�p�B���������`j!F��&�V7�<�P$�ec t&JƸD񝿽��My�y&��=�0m]u�s8���a�u�r5�����$r&��<q�}$L7�x#]tɥ2v(;����O����[�P���LF��~����O�?�FHxd���]��=�9�O�Nn��z���]��@�lBZ���Ӏ��i�vç]�ztz����r��U"PP5 ����w�yC�r����w�K��L%d8��89��ۣ|���-0�1����Q���;I��=�*/�K�T)�Qq�@�m3f>����Oy}(�B�d���?H/��2����k=D�T;��m\A�*��G���Y�f�[�w����n�[kk��|��vǩ��/��_^ a��,t��.����r+�J�e�b��	5����ﳅNI~A��O�S�Q��ٔ�	9z���x݉��B�SυZ�|㢷�t��;B3 .U��q.�^�d< �W���Uԇ8ӑ�]��pħ��-r���zg�W��1a��m�Lq(R��7�x�~���p��wo���ؑo A���!''��	�i�~��X`��3��5荇�g�k_��<��h�[ﰅ�ms��^\����A:�����o���+y�~���2�c��y�ZW
ټ����t�ʀ���˛*`��A�o�2�1o�^v��h�����t�=�Q��M�E���)�%�e2�յ�Icګ �����{�YU�Y��͡2PPPE*f�mn�����lwOw���|�?3��t�m@1�m$F��AI*QPTN7��[k���S�"t��c��}��n�{�9���ֻ޾^������\���&)���x��g=O#c���5��ס6��|_��50zW�����]oݐ�2d>�g�z���ZC��#F�?��72~�$U`�c.�Q��@��[֭[C�'"Cx?7mx���9��=��������p��Л���F���Qc���A���� ��%��Jsk��{i�,Z�P�NqCb�Ϯ$#,0��&�>49rd�ӦM����� ��������[jj����>��駟�u��+��;�w���%���qZ�X�Μ�nrװ��@70t��y4����۩�EҲ������P-t�߹a*��y����Q��Ci�By�ن28���MO�d�$HYu#�l�D�y���V�)���FR��v~Rqx�����#��K/��yr�z���p�By��)�������p�0D�WH$dÆ�" �ؿ��c�46PxE���gM�O>�d���k)j��QM��ko,yS�x��R��~,���<nT7Ld�b��}%I[k��0o�<���Pg* �x��x�,)��Q����;%�|�=F
���q{��|P�ȃk�;���}�<����#����y�,Y��Z���6�NC�mđ�J�P5��LY��^T��>�^��cR
�P��А8s�V͌&^��<�l�ޜMס�ؕܖ�a�<R�_��ϙG���rY�Ʉc�a�l�@�k��������[n�Eƌ/yE��1B@���L���s 5<F�l��m���RK'��6�z#��O����)*�gn進�R:�B
�K%!>i�쑗.��/� �.z �~IH2��X�+**�v�?�P��"�^����GU��Ч(���@�7�*�����ӻvnΐ����Zr������,��/K��(����z��?�zp���
{�e8�d]�z��ըX�M���b,�m�V�������YԲS����A~�'f<U��3�w�=$_��ҷ�i����u9�c:���>��ǨUi�2����gȐ!�77�2B��K�>� hlv�xD`x�3�6m4� D(�ʣ�6�g�}V,X��E�q�0 aL���",$����!��q��t�6���Ɵ�oZ�� 9�Ѓ��?���*������cJգ����@��w�� H���7��)��Њ
�h���+�0JA�0�$:��g�9�<Kv�������r�=�r�V�n#�ԣ]��P�'�f�/D po��mkbn�%�ʲ���Y#��j�7 ���C��!���Ӎ����rڒ��X�x�l� ���.
'�D T I�1<��.�n�9���t� �s��({�կ~%�~�$]n:r� u��@��x��Rhň�T}�ץ9u��f'��>|2�a�_���d�ȑR>t�TT������?T(M-����I���F(0L�H����3H�V�9��B�{����a�{@�����z��uuu�������z)�J�$���w�sst;�š��awG]x��]иhlS��S�����& :������[o��72���1�& ���R�zQ���O �`aVTT0�;~�x�� ����� `�@�B����Cy������\�Zo����
� ���l�!�f��9k������֣�s}�ϴwTcʈ�ذ4��|A��p�|@S0�=`����'�F8'Hvځ�����k��n~Љp��<�&��G�Zxx��K��*/�8O�y{)��x�&�n���8WRF���<�L�e{S3�|Sq�ϙr1�; lex�{�
q���3��0<P��'�~$/����[�֔@����׉v�0&.��RӤ��C�;�e��E��+��3�@p���;� ��C�*������=��P��I�s���L��6�ɔe�q��b+_�����u�Y
R�����)DN��1�~�Ō�q4#����x&�p%MjA-?�Ղ���\��pFG!i��`�B���	�<'��-�#S�r&��x�2u�xB!��ʪ/�d�� st	�i�NCX�e_}T��;�v��0a[P����"U#GK��J�7��L��_~Y��9�hi������q:G���3IF��>|��Ӧ��<�=������^�in]m�xa�t5�n&�_��!��9�m�[�DC�X����\0 s�w��i(��
��o~#|�x�D��N�J�56e^���T`�f�|��xv`v���Ëh�s����k� R�  �����3F4B!����������?�+���Mf>B�x>=�YP��9mw�-F���X}&�"(H�O���6���pk ���Ѝ��i��J/��������q^l������x ��|���q�	��o֬���ˎm�3dB�t�ox��m˳l�+�Qk�LQ��ꌘHZ�!�}x��A�aY��{G�J�q�u�5��t��돚脎�.g�����H&��� �TW׊;��,.IC�mo�F�P=t ��L��g�B��K�=R&���Z���m�Ӭm��5��X��)*�|fN�Za(���2��C�������g �%��H�3��O��C p��E�
�4���.��Qw�����Q�'3�F��
�P3�����XBh��k��}�?@R����-+���� �ّ7��0i��%�� ��X��;�ܵE��k�h>��#E�ŌdU�#��O���&J$������/HOG������H��4=t �����Ç{|ڴ��@��{Og��zMMͨ-5����:� �;�l��/�k��w���Z�;���F�}���ys\��ӃW@א�nl8y*x�S�LɄ���C��׭�`=,�(+��>tq����
������O�ux��p�ǩ־zK� U��m�έ,�gX�q�T�3nO$B� �!t{�E�S%2ڗ���̥cs6�B2t~aL-��*.��q�4yD-������FM�w�?<2xhC��FUXX`����b����
#��a;����z����c��oD\�'=�@����Q�$�e�9��Z�I�a��hi����h:�v�(��g�^Gj �� N!��	���j�������\�1�0$@ZC܇��N^?�|�$W ����s��d�����/G;_��z9�==~�ݥh\u�w���5�e�/*'S��D(�icl��b �&�U��ƌ�Zww'K����H�� ��@¾R�    IDAT\h�Pg�#<��qeRO�|�*���{x-��t����a-8SbI	��A'BS9A]
�B��H�~��G���ʪ�r��kd��}�;����n��O���na�,����%d�
��e�[�����7��C������T�k��e���#���3�<#^�G�1�qK)8�g�^��q��#F��{�a����'��/��������2���>��̀��j��� ��(�'�gq�z��+�����a#��� ��+ :<��S���(�C�{����H�rS5u���:�� ?L�-3��
~�3��!�y3�:n�?D�A�s�w
��r��%h����ƈ�\�s.~ �ʕ�(��z�iJ�L�!��ߑ:p>��B�6ٗ������q���L�8�u�d��C���5
�x��}G�Q����#�`�g�� ��r0�n9���Fm=��1�p�jl8�;�8i���L0�n�)	K$�N"α�iض����d����ܑ��61LpC���t��q�F���!����V��+�<-,��M�W�0�7��;�pY�_綂��@]�M=Fɂ�|!jB�)0�F><7�Ģ)�k�jJ���<u�&�qc�`��Oƍ���qh�z��3OnB�P6씢�|��0k��P
�)"�OG�Y�7��F	����G{`��)C
3�V���.���6���#�悁��+-#+Gȍ�_+cƏ��hTZ�:���1����Τ� lUuo��Lk��[*��45���tn`�!��9��c��~�eܤ}���N��J�瞓���K��G�.�����=t��O��w7~L�����Oeee��0�S�f� }Tu��[C䱿�s�= t���醬�u�����u��qJ��ԣ���*�J.��kfΔ8 �}��O�o�o$)��̿%�$8Z�V����?=��A v����O?�t���/���A#ύ�,@
�!<��~�'
�Qe5sT�����Ob��^����0:^4�����8�8q�)�����j`�x+Xf69[���3�U�t�ǆ{�e3"��G�y\Aa������g�q�3g�ƙ6�EE9\�����{�^��Ru4��{��*�i5�z\h~���@$�~��Y.��b]���7I��y���Ӡ�iJ*����q�' ��)T _9����֭�*�lŮl�I�s���~r����7���'@{ܸ	����h���ʅik풕��bY'�h�L�	�t78�*�R ��C����e��ZY��+��m����a@4'%_JJJ
d��qR1�B��k���kEI"�/6&퉱������A�ƺ�큚R:��1,�ۼ�Z��o��l�h��J�dD�P���kd�ر4ZZ�)�=��C�;�)C�C���^��^�<v�&�`�p~�p���o��-�+��ɧ�.��@i(��=]�Z� ���T���G ����G��z|ڴc��@����{@���YW_;wkC�4t��R\6��p�Z��aV��n���Q����Ӆ�����ud����S7�f��>�����O(0�aQ -�ɵ4�Z	O�h4�ae :��4Z)�@Ȅ�q^mVr�9�P'��Ə��}"_o^:� �WPB/�ދD���Z���f�M�Q��@����7��&�%gr��c���3�ʞ�Z۸G��������}e����u�QR5r���4�쬤�]�{L� ������M�ER`9�HF�E=��.#�P�1 �����svn��<D\?�ό��6�G��F���Q#�]x��o
elJ*C��(�PP2���;��C�0��C���E�d�\De�0�'	/`�����s��5h^}��_�o3\;�^x�p�!��Hg��>��J}�v��Ԃ����x}�Jǌ�����r�����''#�W�ƍ�����d���$m>��1�/�ŗ�L~t��ҿ�DҪ� 2�9�U�P����u��+�OO=�\7"*I��s�&L�SN=C��4Y<���]�A�x}��Y�Z��)�
�(�;��\f^}��7Z���4���`�裏��bs#kjd�<5�u����59��h�</I��`�����A� 2�_\$�~�L�4���o,���NF-��s!>���H�Ǐ�W���ԩ���@��w����k��Pw8&=��:��\�F�ѹ���_��\���[�OmA77���τ���հPF�~�֣:�:�^��5cs�X ܥo��E��iz��VEJ��]=P�Ƕ��f^/�˒8l�==k��)Pa#Z���I^A>3E+z�  �g8�� ?#�~�9g��{".�a�f��!���r9x}�,b�9���+�Ӄ!���Ӛ��1�!�2:OY��O��"��2=��T,ec�¢|�ҏ$��#���4�&��D|���j(����CRȂ$��o��ٷ��f��4��&E��9,m�?��饆LG5\;X���z����`��S���zX�r%;��(3�2����G�O����xn�=�(A�8���+��>�����c-Kە����%٨�ɇ�a������d`Y�Y�ְ#���c��@Jmkk���W_�'�|Rv47J�o�|?FN;F�4V"����K��fY��g�ګK�]c��n�Y!���,8i�
�O#`�SŎ9���<ǣ?&˖-c{c�>JF�)��x�y�q
���|������weŊϥ�v�x�i�`Z1X��y��;Z"�457�������h�ۆK�D8�Gnٜ3⓻�������yN�.H�y�J����ȱcd���4&?x�D:�$���Z�(bb���� �U� ��=�����{��k��U�ܺ������G(�c�RPS@wNz�G��>'��D7!�,�Z=@����o_^>�S�L�ϼJ��@�F��x����ci��䍷�!�4�^��L�>�{�a�Ax�@��W�DPn�%3ب�*O��+��'�eH�>��5�iT�3�k���>/�5��y����$�ټ�Fz�!� Z϶$<lL:>�MYt(�����2^/�����e��1R>t�չ�c�@9
�^�#6�+(ȓ��*y�7~�1����$��/L�>��!�~�xblI޲el0���� �O?]�Iw�:QE��h��k�} �EX� �<����Y֭���i�$T�����D@����A<a�I����b^�QD q��#�<�(��9��n�F�'S��� E���_H{k����d������0$@��ٞ�N/<���wJ���*u"� ]~ :��q�,22&�̵��I0\ ɔK>��s����M��hٮ�����g��J ��vSI���.io�/��J}d.��--MR6d��q��r�	�HQa�!��l�*�!B~�}�/#�H0,��O1�䑷0e�Ar�g�رk)*�d�#������>~_�1�R1�:X���*������:$^I���v%�f�9�i�kR�:-�q��F�S�:vl�O	ZÀ��ɐ�är�H�/p4`�Щg�� }��xUU��)S��!���(����t(����<���| ail��Ek_ce��΍(�	��q����`P1�M�޽B�V�9��"Q�)[?M�֥�F ֜�[o�%�/΀ B��Ե	B�Z��Ҫ��T�RhyiK�)|�ٔm���u�n�?C�#�����̤�J�"������b��A�%/�DR�5�< ���-�qK�_2��Cc����u�R���˧���3N�=�l�w��:��������?Y�;��(C???�^�'N`��ӹ?�	����3RS]''�x<�	x :\;��ߏ{X��de��!���.�o�R���<slʴ�D��;Z�9���&��3����Zy������ˍ��dT
��
Y�'~�a��E�^f��{"��_~!�/��ɹ?9O��x+>[aBS����9d^����\x�%�Ͼ�3w�n�Fy���� MD"�d/(�������͹��`������Q*3ۓy��W��c(�H4����fY��g�s�X���i�w�
���$�ΓM���Yw�'�|,������3O��Qi�
�Fc��=q��n	��Mt��K/͓U_~#��O�U������j����2����8I\^i��&_|�%�0�=��n�iij�m�%�ϓiG!�w�L�4��
  ��s\����D�5k䭷�Ȣ�$��&�O�G.��"�QtEc�u�vy睥�w۶6d9�6w��	�)[%��3wo���x�}ʐiu�R�XSV�B�<K��q�H��h9�.cƍ�с����6�&��`�Ƹ/��"w�����qc=�����ek�P�홾����n��m�[jnn9�/@W�on�;c��Q'�W^��t��޾ӃG�*Dl�G������i4�T�8�j�S�3���K���ŋXǍ��D4���~^�D'A��c�s������HPo����k:jg�p l��Khh�]K�]{k��<˿lC����ހ�ijm���� ��@��b9�jz� �s����Ֆ�r��C���ٻb0�5�&��g��l�i�z�i��ʸ�q'0�P����BIq!��/���*���!�û�ڰ��7��Zn� L�-mfyb��</R$x�0�gksԸ����r�e��Q���y�ݏ(ʳ��ՒHF%/�4����k���N��}�n=Y�H ,���R۰U?����B^��rFIP������Įk3������IQq���,�z��7��'������J�$	9�cv�Ε~Ռ�zZ�n3޵>�,����y���gq�e�H �7 �|�V��ٲi�x�I)�d��J����d��	K�%��ɛo�%>x�$�m�M�駝 ���K$��$]1��Bk_8�y����o/{_^|auҽ��x\	��C�4�8Of�8SN:�T�y�RS�]���s4�YAD�'�a9>9��e���#��Տy�����3t"t�@KS��̓��Y&�J��̫���!�� �˖��t�/�A���V/��L�z[������`�`nH���sf�Ӻ�8��'�0:l�>��P���4$R��d\\)D�Ҍ<�X:jTUl���s���]X8�io��㾛���g��{����sg�]s�j��~2�lK�<���:���Y�VX��, �f�)�N&O�LP�Fd��K��^���v����Q��P͡c=��z� �y?E��\�	��e��=�NF U�L�A�]���<޺�Z�� ����E�p���H����Kz`�[$d�'����ю��u�������M(/��z7�B���~��-(�!�a$s��B�C�7a|F=^ǰ�J�����Qb��*U��qG3C�������1�'Ms��og� �Z�cIӇω�U��H/��"�(���0�v��)ϻo�%�Jʀ������0=�ɓ�7�xC��r	eG1MJ���|FjP� i��M�&d���pP��
��̔3��-.7�y"��_����S֮�Zܐq���@:��8���.,#ÂR�l�r����J7��1�L ���G���%�v˒���m�ϒ�d@I��y�8�쟊'�_�����=�<��p��2x@!k��Q�ȃR�u��^�J��Jd��,k����Η�h��!O?�'��[/^oJ�n���i�+
��W_)��1]�)���5�w�b(��,p��I>W(1^|��r�i?&�œ�� ��~k�t�D䰩�K�H�D��u�꫕��SOJ��K�̼�>L"�pmod�eC}��?�ᡓ3b#!���k�˔c��m��L�m��[�NS�*���@om�$� Q#<?�<&��sc�	����?��踱��;�ȃ���x��w��n���Y������[k���KB�Μ����s�������g<_�h�J��d�ɝ�w�ѢF�H!� � ��T��^��+���O�����<;�O�Y��ɘ�Y�tuf$Vy6���j��� `)�U�#��e������e�����߬aJ���En��4�h���O�T�yP-Z$�m��LI���΍ކ�s�}Nݹ3�h�D����g���a�P;������N����f��M��ۅ���9a(q�wv��!d���WR�wȭc��;���{��o��m`������Q����6D��$ =\�O��.���C��K ��ٳ��^�T2&�%�tDP�,.7���b8uܷ7l�燔�ɠ�eR�
�H���Ь!������U�\+�{���N�W>Z��̞5K6m\/~�Z"�4�8���yF�=	���t'��ר�9]C§�r�\|٥|�._P�^�Y��A���U���ĕ씠Wd���o��������K6l�,�^|V����~�q������Ҷ��V�ԚR��!��m{R�����՛���o��?]&Ņy��tK��ҁ��+��c�9�a��;�λf����i�KDQ�>��r�u72<����J����o��o��2j�Xqy�,X	�g�|���K.��x�۷��<V@׍9c���������� ����Ym��)��:1��Q�$��(�c���������y����W<�.��̐{UUUt���M=�_�����?a���t��j���~�� �Cj'��Љ�,�\��Y�Ko��jyn��<tq�F��$G~@z�����G!% �����CZl�D g�;*��],G��X��T2�c�E" Ԁo�Y��R�s��/�?,PS��} ,� u�Ft&g�R��ap#����}�[�������f݀,�r׀nB�����'g�6jK����Zp�%x�AY��J����w�r�Jn� ���NS(3J�Y��`0cc����)�� f�H$���#�3���JO���/���^(�y����q����2�H�ϔ�a|] ���腯�-�[�9�+�J:����rgM:�Q�2��;�6\Rho*��m�Ŧ���ж���˿�a��� Gqb5t�o��L��w�lټI|��j��?R&%����[�Cw�f�^�D]�\�y��(�����У������$!_B�~��]y�u2|�$I���j�72����㏔iS�0��(��ӨJ4����A�
"1I�x�y�n]��~���g�ϓ��V��Z&\|�{����I���g�}��i��#��� ���_��K0����l<��nS�Ҧ1��H"�5�� �y�?'���J~z�9�#,�u[�aC�V��vYT �3�1��vw�qh��Z�rf�(��gD(˨�9#��_`��YfUû�j#BM--���D\����XgnF��WUU�Ǐ��ԩG�S������x�?���. }{mÜ���#w�CW �t�:�>7���e�N��C'�s���	氌I&A}���`���2�A�B�}���#�2��H��բ�=Q�ҝ��q�FJ�z��4^�sõ%S��]��@ǢO����> l�aiY$D�[Z-8$zG8�z�0@*�#���]m�]�ȃ1��Zq�m�}W�VJ��F�|�8*  \��O�>��5�\\Ê_���;����䇂#QP�V֣��Y����5�m @�;�`��9���U�|��r���k��"d����~[n���O�'7!h4�I�����_p>u�Y���q���
/�/��O(f[J�,c(#C���;���Ź���D����g�	��n8���Ɏ�RTR"�����!Sq�������]� �^���x�H�c�?�&5�k�~��K�~�"� ��G���"�x��	�E;�a�����ʱ���7k���G��=B�>r���	���F((o��;)?�9!B��(�|��Ȋ��Y�d��/%�$�G�کo���O�~�iS��{��t�B\����r�����7`J�P˭�1�!�DI���x$*��͓�W��g�A�_��f�    IDAT���:{Է+�gᬰԮ �������e`l���2�3�\4��.�)"u��	������t\K[��l�c�a~x]�ek	�F�JL�8�)�����B�c�{赵ߎ���6�����ݑ✠�^��=g�]\7H�\@�0�pZ�,J��24���f۹���,xd��8�t`\^.���� ��b������U|^;�����6%��>p����vs*V;�c � �P{�PtOW7���65�q"�)���]��E�����Co�ꦇ��N0�nTR\�ܦ�es�;u�� Ǝ��B�R�B+�0�?��3����xO �����S\P�����8C�1VL\��\%�K�����v4�A$W\y%������ҥr�m��P�&:7J{^b��<�p���!��(n��n`�ߢ���Ņa	����=���F�T#������$H�\�!�ڻCJ� �������I�?�`��Bt�������z������ :��N@W�+�^u���:�16�;�Q�;�ᥗ_I�|��eS�6�g���޻�ߛ�2�=2u�����e����d������Q��~t�����D#�+�f�aj�jF�:_X|�B�⋵���(�n\MB�ߕ�d�[��`� =*���������C�܈��n�QFTUr]G�*�)XR� 2�����yLm$�)F��z�IY��7r�Y����²���@�}k]�Y&�u.���eg
�0�(+h�#�\��G��͗::8�U[�[ɴNG(Ӷ��� S��p������ɘ��@G�]Iq����d��>ߟ߈��zc�l"�:��T*�H���T*�,(��z��w��z��'��>p������
�v�w�w�O�~�_��z?���j���.��va(�%�7�5�סl�vk͜���R@Ǆt�:����ߙk׍Håz�s�`çl�����Cr��M������IK�4K��.t3 ��U@�E�J��)ET|F��W!_Y�>��� 1� ������L�Qc�p�A`Jh�Ul��J��ׯ]�@�2Z"�VQo �]�#�8�lq{}ѐ;Hq]�fO����T�w�D�+�;Is���ϸf��7�h��Qs@ �G�|,������_J��cy�~'��w�@����j �AÊ�is�Q�z���W��I���@G��.�x!�N������c9�Pؔ&l.��NK(/Lu��_x�X�������SO=%���W:!���d��Q���I$�!t���g�U����`
�!w��^�Bg4�u.-zu�r���Q���h�-^_P�xse{Сh��CR��g�i:B�)��5`+Al:E��+��!C*�+�?�B�{��Y���ē�,�g}�UW�77��U��CʱGM�SN:Q����t��q[����K,�)��ɘ�c����Db.Y��Fn��vY�n��|iqǐ���=��䔓��?P �n����W>�x99 ��DX����e�U����̑���Iӎ���] 4�	JOO��f�e��26�޼YfϺ��^~�E2j�h���N-�� ������ �[�F��t��iA�p+L4�3���������&v�S�R`J��{�G�K///o���z��r�z\�~.�k���
�\^���I��r�bX�"��l�ad�+�r��D����'�N�bn�;	# ��?�*a�)�Ѧ�m X@���v����֧ˤ���\Vf����|⳸~*�����V�eܺ����{�q�J&a���E�﴾o�;�J���t�g�ϛ��=���o��/�"yM.�f�^�>��������cUU='�A[VyN�M"gW/[��aog�]C��T(*Mϧ^:7+�@n7����Dx����m��3��A;��а�	YgY����!~�ӄ �^��ca{&����D S� �n,T��AO�;˖�􂜳��X�d��d�8?��Y�9�\ӍJ<���#�=��#]��0u����I쨟5����,���u�+2�Ύ��� �A�6�Ϻ�������EaB�y�2��+��T�yWg'�S7\|7H��#����_Ia=pͧ��Ν+-�t��!P
��n�;�clChZ�0lhzj��!�إ����5�w���RW�H�����N���Er֙�ɹg�#��y�meg#Q-'�D?�7����&�M�S�'xL,{�����䜳ϓ)S�1�&"n�W^ye`J}]IqhO��`��r�[}������ek�\�2��)#T �����H���z)++���+�~�	��]�(E*�E�s4Թ���dPy�~!
��s��=�)�@�P"�����#yy�<i��&>?������F�I'�B�d�-��V�u�|�z�i� ���G��Ȍ�~*.wP֭�$�f�Gc(�H:��aY߸�c��n��'I4��?�@����44�Ka^����`H�8�h��a"ͅ�F0/>��2~�$q�CҸ�I>�Ш`:s�ܣ��j�ԇC��I�E(��~�`���W����cO@?�[�'��u�9m��L�'����\ӈ �J��w�>��b��n�]^�7�ЅH��r����~���x<����3�2�&~�#*�m���NN�?n*v�5�4��E�=E�=w.+��td %�v�L�~����@z�{j�!���S�A�.y:�N�yq=n�����~����%%%%�{��{@��{m]��-��9�aM+����. =7��޹Z����4e`J�2-����LiP�nej,:=t� M�$�6�i�(@H���X�5�U�?�KW0t��8U@X�D%�f�� X�X��^M*�������z,j��я������������=�8�O�Ȋ˜Ob&���m8�>��^�.8G͡�k���s�E��g_|.���{$�`@;t�\z�E�QbC$�:��膈V�X�=����b�˂!�^�tAT�7o�44� )��n�w��A���e��[o%�:�6bk�`���1A:
����&O?�������&Ç���~r�L?�t	�C�!�j�\1/�aYrT�*�A�l�����f}��I��Ah�}0��)7��/!��To� :T�Tb�����z��6�`|�yϜy��#1��/Vʜ�"���JI�㒲A�r�YgɑG%�������CsdҸ�r��J\�v��s�Γ?=��$R]�JvK*2d@*�W�\$���dI�<��'k�?�)�׬��?-޴�),)d�e}��je�����?�7%�B�u�R��~���^9r�x|E�̳��SO<.�-;$�3�tt-�<���Η�O<�skǎ�2�ŗd��o����D&M�W\���hj��@I�\@��V7"i��3�Gv�C��pDX���u����LE�@xq~׆LJb�=	
~�f%�߭��4Շ�	�\�_��d	��1aܬÓ�����!��;�n�Ѿ�VO�t�rA��8���r���H����x�:��5�?^�~���әJ�V���VYY���\�����-[�T�m�y����G��/aH�G�/�K@wz��@��t͟s3�ޯ�ߋ��6�)�9�����}��ٗʲ:�T@��.zJƤ��KVCh0,t���=��<, r�c'��E��K/������G�Y�~�C�u��{.4���Kx�>��U�u������l/7Ε��s�c@��qɥ����g�#����7:�������O:�Q	�����<t*E/��=��t��9��Xnf7�9�!=�w��}����u`�Cy!<���-ez~^Ȕ�С.�����C�����8�;��6y��e��Ik�S5\N:�X9|�a�v�#C9�ea�>m~O��u�>7�����=oܱM>��}ٸq#K��#�0q?�A#���Ȓ�A#.��&���d�f���<����u.;�@��k%����pc]�,y{)��g���JU�p֫��Ѣp���`�;R���j��Kgw\z�1y��Ǎ��K����2��J.��J9�)�J��/�yϒo֬���ߓ�T""Ⴐ\y��t�#k�m�;︋�K �K"�J#��C9Dn��&�6Jbɠ���[2��Gd��zI�{�]�G���\p��\+�i���+�q����e��I�J�dGS+�㰿m��8���@~��-:���Q�j��x����_ UBlA��ˈ�a̱#�`�m�Z�����3J����Y�F���r�>u%���G�E��Y 4�z��h��Yҭ��2un��x�C2�`�t�v���(�g�}�OrM���	x��:V:��@�/���\RR����e��7U�{@߼yse����[[ZN@��7ߴZ���G�;@w� =���J��,��4��9A\����ai�����I����V����F���,d+�j'M.�eC&�5 ��k��@�I��FH�c��q+�Z%/��"7Sd���[ax����=�hB�]��s��k�ל�7��E���ޮ��M������+�#�@��Dc�Ŋ/�C�b�g����~%%�����an$̱�Dx�y���.x�f�����e5�Hy�0YՀ�3�W�X��q�y\^���s�]f�A���Rr���[ں�OO�Y����tw�Iq~H�-��U#�_�	�2�+���p�:��v�1)�d�$�;Z��y5P�?|D�m��R4�,{�C���d��o��2UxN@�Qk]Ӎ{K����k2�w�[ @G�� ��t�tK#$����K�P,�?@P&ٍ0��%E���[o�SO̕�?JN�~�J�ISK�<9�Yy��$k�`���.jÑv�醛	�ȵ��j���;d���$���ϕ����\z�e2}���ò~m��9���\��xܐ����[�M�&7̼QʇVIO�+_~Uf�}�Dc��c0K 1��zƙӥ~�V���"���
���^*��Gb1�45��1 ����Nfg���c���W�c�2�/$J�BlLr��7v�hF��k70 �!w�ߐEs=I����5�������mt=Q;��!��AF�׫7��y�8�Ο�Juz_��b�s���>���
��{Ů�[ϗk�8 ME��_+L���"��?3hА[��j�{�6m����斖���;����:�ܔ,�c��}�����UZ�=��:�p6��|����-A���ht]������ɘ�
�Ze2NX���VgA�	)�k����6�����
+C��i�u�`�k�u����KF�5�r�G�M��z�}���Y�^�P{0?��-߃��0,���~hɃ�����=��I�I&e��2q�x\V��a��c�&H�s$j�O�Q ���~Y��G<mm� �{�5W3���0^�,z�H�vC%�7�)��ȑ�3m�:�̳g��B��S�:���OɳO?%q��MD%�ʸ�c���+#1�3�~�>�G"�����iˏ|���f�VkG+��[�7�~O:�F

��?��W�z[�������GC�N$�R$y�RR�z �n06��%X���4�N��D/FE��G����>�46��{����O��L?s���ij���@�4O�۶I8ֻ!}�'r��Wˁ,�����~&��e��a�/db��ӟ�\�8c�����Z'��0s�x��S�4�Ia~�u�W^~�:Z��Y��}��[��u��<i�E1��2`� !?r#DHi����4� ��ۏ����ζ��E���Lr�~c�=�Ls?��W�A����t�(b���0�$ё#�8o�kJ���N��VL�u
�N'��h����1^����9��H���ԝ�`� g�u:2;��p^����kC�G�w��}E��w,N�ޕa����x����c�������񲲡�ٛ<�����VW��ަ��Sn���v�2�{��aNْ�t�hH���Y����e���t�#�JK֡�	�6;Dx,{_g=g%ǹ�4�XÎ�*\����F2&�̥g"	6�ߏ�� .�}�%��/�!�Pm,�M!w :Y0N؀8&>l##���ǐ;<t�Ҽ�z_����d��͆��t���t�a��C��g�ʿ������]�K���d�VJ�ƀ��75�.#�:k�;t�$Z�0B����'�1Mq��W�b�MT�G����s��4��pg�Y�%�ǆ<��W\*�g�e�E�u�-�Qy�g��g�$��.���WH��@~��B�l�^. ��W)��֍��e�늕��1�%��3b��3����%6���na����'#��9��#KS${�;7e]C�D%=z��R�q1��M6�"�c����P#�̔�Ӝx��2s�L),-����Ȝ��T��wJ^�QZĸM=t���ӟ��*�G-~Kf�w�l޲V����=�i�!��s�9�ܟȀ���>���+�V}-�8��Mn��z�T����2i���3!��X)ιO6lX#���ƀ�x�)'�	'�H�%��'��˹p������%�pKKk[Ы�&9��'� :*'��Ã1�3W@���6|(SOcƌfd)�o�*�۪��RJcݓ�8а�|���
�oҰu89
��OI4Es��y�m03�]��d/x�9W�� �^�XQ�^Hd뜯�������h���:Q�G����m)**�=h��?���v���0��t���ﵵ�C�n�����|:�s���>��!����5,�A�<�z��\�{R�S�E-݀/� �"��0��!�xm�1H��FU���5[if�\ljx!tۗ�w����f�	qA��WԖ;InGu���|��]�����E=nI0,�3�r�~�)./LO���#�!����ss�*���nk��%�eC����t��}))N=t>Ӵ�1���~���R\TD/ =a�xv��:����� _TR��P%�¶	�沰�=��3�d���*/��JB tj�\2�B���i  �!���E����<tԎ�4%ii�ˋ/Γ'Lbݝ�/?,�K
d���ȱ�#y�̨��l
�xn)K���87Y�ɍ�&ʌ�^����	�ɯ�k:t�C��ko/�9s�H͖j:����O�v�K@l�6����s�v�pQی��}��_�
B�X�W�!	��&�����_|"o���Q�^�;v"�`i�@Y�n��{�U΃T�S�!c|b��1BN<��r�T����h�,xy��ul���-ބ1��>��s��'KI� �����w?���^-ItK#�cG��#Gˌ���>�$MQy��7e႗ؼ�(��V�C~
��^6xC��,]&�GT��7�T7ZbqW�����1T �HX��M�iгg�-�Uc�����-RFa�!C�m��))	·��J���F�{M�c�nG+]�.�
���m��(l��	�r�v�Ԣ��wz��cr
���B9���]y�zM���s�]Y �Fh�(��k�ʲ�S���l���ksqq���0aҳ(���=����!�f755�@���3��M8'�}M�`�\�X�q
�wt�i��0�q�P��^�̝,�ﵤ���k ZI&�bۄ���&i��B�JnSOݹ0p�~͂��ԅﱊQh��
9R���-����ԓI�׊1A����à�+a	bd�v�k�ؗ_&?=�<#����еl��-[����f�ֲ�Հ`v�H3�ދ�"n7�����ʀ�bR^.�-�d�x��j�� �&�x���<�5R�����^zi>+f^� �,w��ˋ�]w�%��U3}C��F7y�¢|F6�:g��N Rz|����ɣ�<$�d\�����-�Ǎ��r�C�I��c+&����A��0gA�[�x!��%���g��������\*�ϙ#��[�ݍ��L�>8P�� ��D�-ks)��3c�FP������й����e`u	diŐ��8������|�VV�_(���$T��-�Ұ��Q���,3���{p>|G���$!n�l�yhW�c�����$�C�R�u��:�D%��CY`�46� 4
|=r���?H��;e3�ښ��G���aTc@�[    IDAT���/�@���QJc��f���%MKk[;� Z�nٴ�s��1H֢������:�tI�����3貇{�� с�B�ύ�t)#ќ�1�)�6f�}Έ2�ɤ� [=��g��y���;��2b���=�/ ��=z�,��O3D��`g������1���#�pHlD�ߑג���x��o�w��z�^lϧ�����
�!�D�"�d�5��w��/�ǉ'�'0羰7�wS�X]��z���֖�`��ё	�k���䲷������CW������w*�8����lo'X�G���1��� �h�.F|��Wq^�֧e���7�Ζ��h�zX|7�Q�-�~�t�֎!��>�@^x�%
� ��)Y�{�F�9c ���_&?9�<�n��uv��ͥ�����)GS	�eg�k�ϐ��g�`Z���.���ȵ�r��V-��o��l���%�H�:`h����GE�S���<�b�/�#�h����P��^�y���8q��/�ǐ��w���1�L�;n¶9<��g^Cz�⛓.��t$����O=Ab^yY�T��Ɂ��+cƎ��J3s�~c��#�=l7.��҇���� �����}�p��lq	#�i�W^[�<p����L�ԍy���̬'�I-).#���	7O�}��s�	���F�U�C�4][��t|�)��bz$��MM?��n�s���~?T��V�Ѿ�zq���TQ�5��cF�y�%�+m��/s~���覛n��#�sk{�|��'�[��-�'ĺ L�s8�IƠw�^�T��]�&x�U�k�FN���j��i����=�[x)�s��X�xA�=�,�������'�O������4���L!fO���A�ݿ2=k�p⧫�Owʅ��
�;�4�/f����f�9���;�sw��.�[���k�t�ʃ�i�t� JC�O'��)a�p[�"������ۅqM&��D"ѝH$���ԗ^����7nܸ=��9��0p���o�n�����L�� �r9�꽡�&�f;P��ŎcVz��I�9*]����?�sC2��Ԝ��K7]0N�aO@��q��3�t[�2��4K��<�,z�&߅Li�|Fp :u/@�
��G����ݴ�w���ح/g��tLw<���j@]�H��� �	�>� ��r՗����Xv�T1cHjC������͏M
�iJu|,9��c��媶�K�[8.K�_��#s��e#'�9#��ΗE��=��2/������}��:`�ǧ�f�wJ�i�D>�?�<��Ò�F��ɓ��'���J)., k޹Q��� ���������yP��cO<Ξ���/e�~��J�tZ����%��Ï�v�~Ŗ��|�G!"�*)�6gq:�QNTǮ�y�\;�w����i8^׍�k}_�w�kέL����w�~e���q���l����zC���������ץ�讪�"�Q��O>2��-�7rnAB��y2!�l[Z�/O�)`H\5�m�0���H�U@�Ա>�0"���<㵻��֛���yy4�����h�7�!~��=ww0�������<.W(���].W^:�����+�AH�.u:������wR��<FBw��/����0�"Io:킢�7�D�]�9��K]�k�2���R3�mL�t:�I���d�ek�R`�x<����tʡf��8���3�B�>U��*�I0>�;�M&S�D"�����t����ʷ"�-��ō����{����������.oؾ�����3᡿��+t<I�ݚ�'�bv^+&��Nv�h���	��sjN*����ݹ����x�y�a��AO���n��ƅz3���!� �� &�F�I*T!,�m�6~�ш��s �@�� ���s'��1:�ny� *��f�g�n�}�]Ҳv�:���F�_Q1Y�`��9`�����j�q}��yʐ��F��B:��<�ϟO�D6 �P�⼂s�	��E�؂��%U!σq�R�үA����YW�W"��K�b"�/���="�xL~t�r�qGKQA÷�EV2�K�\/Z�����+��ڵ4�?`YHu��կd�����q�[��L|�!�Z�E���	I�bt��|���;�%3StOz���HO���Z����ah�qNP�յd6@��S�=s��}A	}�{	L:t Lݸ��΀����i^ ��x��h,E��O>� :N@�}j9+�Hf}�&���(��	��T˹��2�v�(�Ĝ�QK�8����5��¢"��B�`���B��	�I��EZ��l��1c��ؿ��C�td���O'����;<ֿ��T	7�ľ�3�:���^nPF��kύ
hܞE��D�钒��g"	�Y���Ds�;{z=.rm۶��"��JKK�Ȭ����_5x{{���8'��Cw���V��N�\OY�^]�ȫ!���[��*&����q��������{v��s�zz�6F��~�}���}mNY����#�n7,b��БG�=bQwvF�Qj��̳sv�l3��=:BRPZS@G����U��mQN6#����,[���_B���,�|�v��}�]�j�*n���C9���zn�M�e61�!M�yJ'�8s���O�C�_�4�5x|y$�ͺ�.�����2z�`�"�SB�cF��w�Ͽ$�=���bQ9������N��%%R���y����d+.�(��Ի{��!��zf`�{�|�̙#�p�\����T�x�<住��{�-�7��;%>l�P�c��C�����(�8�̸���ܵi�k��߹kE?���it9>���~_��Q�:oё��]{�����Zɢ���Q���曥��J��c��_� in�o3:�(ڵP�z'A�mRu�8��Y�v5C 3�[��� �XxLA�L|83Æ�ҲA�A�I��&��f������*���L��F�u��]ܿ����~8�ޏ���o�����z�3�����t�.d����ML �ٮ� H���uc��P�w���P������hL��yNpvޓ~�/@WK\�Q=CJ�!w�/�QΚ1�r��  ح����x�˴����C�cO�y�ь@8��Б�5����O���37m�~{
��
Н:�n<�	��%��^�
������;I�����t!� ��[������%}	!�Nc0�~���*��X��>����'<t�� �^~&��ȑ�@�KC����������N���/�Ѵ�����s�Qrތ�2��T��!��P:��/J5G��2N���y�����c������+����1���ݏd�l �����:����z�N@��8���n���}��i,;��]mi;g�����_�aZ��OP	�9�����9�N���1��[n!X�wG��e�W_3��a�z�?x�؋2M�,�67R��M�J��Qf��;�s�3}�%m^�͔0Gp�	'ʀA��o7��M�Ic�m�v���P�>x� ���x�	WXٰ�#�Ñ��|�����a���Pucp��uR�3?��*��p)<,l�*��;��cq点s3��6z ��b�̵�N�}w:׋p��	 V��y����)���R<��2�%��ˋ�`�-�[]�PVX���N{ح��'�d^��=�Н�n�S91^��>�� ��C��&<T}���2-���3�<+�qVh`c<��9J�x��4��N��([�[�x��'I�C�3��`p ��r�}�)[�!w�͡�y����0ec�&�
f�O:{�2o�|��Gc���<\.:��2b�[W����FJ�t�2u��	��P#*��Q	\��>���I��5�tcs{Y��`���Ѓ��֚j�  )���ȴQ�\=۠j�Iq}������\�`W޻3䮟����3e���{.���:ס���o�����п]���k׬!S?���ת*M*w�Vgdӄ��o�0ciS$�5ʒ��Au�'��{c1��C�Ȕi�р}���g��O�kbFӠD7a�82dpzРA��8���? �f��u��� �m��ZZZ�Bٚ�ⲡ��IqN0�0�2��y(&��=��S�x��[_����;�s��ר9)�lY.���ǔI�ou�zr'�=wss~_n*`W���ԟ}�1d���<z�#��֧T೒�*�]��J��� �y��-=�(�����mx/g~��`�C��K�������8�[=�,���� БCG�Z~(L��駟A��c�1F����gH��D�yt�2��e�E�:_]�.}��!�h�J@ ���-�����z. t���Q�@E��0R"n됟}�����Q�0~��;�,�<i"��F*�4`�m��m��^�]�z������9�����oP��t�`~���L�9q���S~�Q�����v% :���͝k�@���H��Q��W$)lw7����7�ܭ�o�j fg�#�n/�b<���q�4{)��[�b�0:��� /}��_KSS��z",���}njA��kJ��17�mj`�a�qR�Ǯ1԰������(�'N �]	�?�Qth��c�9�$+h 3[Q1$5`���'�t����<�����O}���q�������@w��NpL:� :�Lφ�mr�����H��A����������Z����P��g�F8��6�7u�Y����2�﹀�*^ #(�M�:�ߥ@����Ŋ�,'��Z�<cd�u���C�ܟ��@g�u�.�U#�@��,��動+�g����M���c��x !�����O���Cc�B]�S�Ç�+��YK���m�L"��<y2A5��0��Ȃ�/��w���Hp;��U?�Cw:Ꝼ#)ָ?���R��M���&oi�!555dF���_��q~�z\.���#˿������'���o�Ap����e_9r�)�K��)���O�}���{Ri�#M#�R��#z��c�k=w�؝[Y_^���=�
��f[�5����ݭ�\=�jM�ed�������D�1�=襰z�W�joi5M��Eǘ�Ψ�3��9�#��5��|$�[}w��v{��%J�{�O$(�4bd�R Ł����=ʋ�3�G��n��c��>bİTQQ���N;m�a�����p�w77����tr��0�lUXF�a��܀R)nz���tf��.,��Ex�
�
 �������'�?l�x���,U ����B�p/�O=x\�^C_�s��h�g���PEm����דN:I�2���z�m�z@�H/8'��0���G"]8�6�Шf�l�fB�C��&)��90k�ol�<t�a`g���
�С#�+b7+\#Y�w�A�_q	� �gr�6�2�����4�#P#SO��r�*���`
`\�^���3N�l�	���9x�������k�G!Db��^J�媫���Ξ��«A�,"�����{�Ҵc���+���+ḫ�Ήk�|f�	�u�����| ���&>��;"N���~���Z���P'�v�-��*O>�4�XyhܑLI<�#�!�3F()V%?����m�/�γQ�]oh�y��s�͖�4���jm�8q]�!}ʵ���6gT������I���p�M2tX��$�\?� ᙺ�v�۰vI����=a�A�:z���eGC��+����S�Ǭ}�?4=n��x�����^�M���Q�=�J��,x���;9�TYY��SO=�@ߛI��t�Cojn>V" �.  �SC��� .((�������J��+��@�s3�ݢ�gҗ���Ԓ)=N�JVZ�i��
��ܿ3����nR
��x��0C��C=��K�u�=�v�KDM* ��SN@�	l�����9���R�i�Z58+}H1��27g>�V!�5�		�_��J��J޷n��j���nI-	�,DC�F�0�lL0�~of�7��?������dl���� �,L�9uΡr�����[�nWuK{��TkI��U��s�=g;~��6�E���Ԇ�2ܕ�q����w���z��]�x�x��y�<1�@"ɉq���(w�
��]]ʵ�5Ljs�ߜ��3�܇R��������Ke�!	�\��F�< ]]���z�֕흽���h�/�{���L�e���� �X3���8: WrH�����9(R�}XZ�X��[7������s�ޠD�^k5�طo�F�!�B<1���FҡXt�MP�д,��~��Ͳ,��R�!2�I
Y��^6?��V ���ʳm��}�=�L��J�b��s�ѿ��3xx�X��,t5J4Dg~/e�t�7�P��U�b�U#Gд�3�y�p9��y�=���X �XF�ѥ0M�u���	�^S3jѹ�^vǴi�-����������z6��: �X�"lІ2W'a물�]@�h�T�nQ�k�8��f�4y�t#��]��m����צ(8���3�M_c%Q7�}=�V��ժ��7�md3
��{����.`@�X2��1�eKiū���#�ҜE����B�:�����]��@�1Lq���Y6�sLN����,Xxi
�#Vq1'�!��x��(U�6�R�{�Ĳ6�餌J \���둕��t�[?�c��hG3�Gc�^>\��B��u2A�:�<�<�߽�RMJ+KaZ��}�J�2G�(KA�A��2jhh���56졢P�ǃ5`�� ����9ƪ����j��:~�`��b
�����?bM�<�UQC����,[A<� 5��M�`�P���2inՉ�eS�%u}u@l�\(dm�ϳ/���*�S�7��k���Op�jV�'�o�T�7�~,E�I���&ڸq#�ܱ����Ö:� ���(n�4de����E�	"Կ���n��|r���r79�f�����4m���o�h�~� @G�7/Bbh
%����V@O!)�K.�k{��������!c�wtv~( ���6�E$O\�
� 6�Ѕ0��pi����`n:0ʙ��#�_��$��sũ֏wM��&�lz;F�ǧ�v�nF���{,���ŵa���
+C��b@�iK�.w�sc�.@�x����)���9).w :HCҬ�9٬�\������pګ`�,���q�J ��k�eW?��ݽ=LM�� �`Ҳ9�.p�����:��*�b����P��
f�R��\���fJ�<B(,N��ڐ@�0J4&1n'åDpe�#A�(-��,�c�"~,�}��T�#�����ø&BAPJ�Z[$Vo${4c�1r�x��R��5�=�^
C$�k0�7�IR���^^��~��S{sE���6���CL��8 ���"�_�
�&��kȿG��W�0�������s������3���+�N�ux��L��u� ��x��bQZ��{!�����X?�&�1dmʹ����z�4t��o�q�M�O���
��\r>	e����&O��̂ǒ%KY���v(�즇�
24�Y�f�BO����i޼K~x�3���B���z@�ٲsL�����^jй�ظܱ���R��+B@��&�"����Ys5����m�� �dm0ǳ�8�fCc��aи>~�� "�Q˦�L|u����㋡��I1'��O�3��	��g]]=�d���Pz `|}�~I0��
1@ ��.w
� �r!zOgW�s;(_75��D+�r�3�q��-$.	t ւ��M7�ĭGC��� .@���� �́`�DăU�ÜBa�qͽ�G��en,�q�3uw���?�-�g�y��e��H
���Z,+��J��[o�p\��x�"�%�H�8U���S�#]�&1������Y�I����I�N (ݴxn��.��LH�k��ڽ?��ښБǬ��{.М%�˺��u� ]�o!����{���dh�i�[}�l{l�^�q�<�%�׻���A��MTI �k��pW<X��~�� �޵K(X�&�B����8��(�W~��/X'ثX?z] �TΈ��{O=i<iL��.*�,��"�0�:iJ���瞣���S���x�1r������>ztm���q��    IDAT��ً/�w�ĉG	����_mz@��������-�D-�J�� %��PX�p�C  ង�P��ծ.wԱڛV�� �	�� `��]]��+��1B���Z
,*��	AaU�����ffԾ�B�}�	�K`����Y�
�lM@W��zI�tV���%�Q������y\�,_{TEc�2�x���6�����s�cb��ڱ�@d	�缀��ݧ�BA3ڽ�n�wqm��O���:��\�˵K��tv���x��|�qq�KG�t���p�%0�݌���PT���1^�1,1Ia��g��ռ]xg��)��Mn*3\cp��3�폊�Xgw-|�Yzb����D!(8�
6�.<2��~����{j(@Wk�V�ct����~���	���z.u��~u@O	5B���r�����c�<����V��<����~M���tF�D�	�y١;7#ed�h�J��5����$��� ���h(]�d��(��c�МS�RQq1��h�ԡ;!*�^��FR\&J�H���G��'��j����y?�4阦������}L?�_tvv^��'X���ƅG8@��Ol ��ᚄE�V�?��k���+��o���9��7���`U�4gu�kW�7�3�PUW�-��)� �p��0?"`:;��㽲=Xj{�6����,|�/P�2���:@ ���Q:@��b9�,�<�nߡ ����P�4�8�H�?>�9�Tn����̋��9(]q�zB�qm�`A�d��
��eP�&w�2���{w_?��|%��r%}��'�3Y3e@2���ऽ��i�Β3Б�d(lq�X�$��iI��[�7�`�	��M�={3�bU��J���8,n~�6n�FO��i&4A���r;�\0>�>�^�.�L�{���meZ+�����!�X�m��[�|n_�{(yh�X��G�*V��͉�0�sѦIq�;����S2���M���[osO�ޞ~Np��Zh�%����St��P@W������ظ������P����RY�C#�GҬc����Ù|jݗk��n�������Y��S@�Å��/�}����~���ݻ��4��eWW�� tX許U~k��S_OӦL��ѣ)R{g'�45Q�b::(j2�5v��&N�vi���'����=M�z6��ט+���d8���hob��=����kp��:�p���~�1�x�2�M<���dY �|6���n\�6�G�qzꩧ�?��'�����o4�,��a����C�r �31s�I�U�w���6�����hP���ր�z;�9�x�r��P��Ɲq�:��X�C&�VUݖP�6m�B�����i�6������U�:b�GyE)�����БP<G�$�bnuU �Q��b� p�#�1h� B��M]�G0�-4<�~(th�������?��v�i���*).�����Hz�<�����C������̮�6;[�AS-�����A1���5�܍Rf\��fqr~�:�*�Jx$��g �p�C^>@�z@)��I��yʴ,�#\���������V��a$N��h�t(e�v�c�s	:Ƴe����!mc�-��#)
��CDF1*.�
� "���g���e�m���P�sX)���D�.�>&1zt��?��À�����g<�}Ϟ=��4��eOO�<��|`����ƪ������Q5�t.���&j���Lݝ]��n����w�VNz�'�
�~�<�5n�i��٦jj|��r�HD,x�W&�^� n@���]_�2r���Y�9�Xͣ�`C}�Qt�y�ѬY�0��쫥��-~�V��.�@�s���W1h�8��p��غ�˽/FO.|����x	[�]�C��~�(Dv�T�7�˖>�cy�0*--���	��{��ՌߵbA�Ac�x��>^ݒ���X�9U!�$hB�s�<��l��*�,=�!��`N�c׸�=�d����!�jTD)T�B֥���'�U���=�2��tф$D�R�����-Nq�����p-$�{�ŜHQq8B�<�A��!���h�R2�fpL��T��V�(Q-��>nKD�O�^�R��M��w#EpP�d0�����'�'�C�U���Ög$e	� �Ca%XK)/I<������F��DZb׼o$7���4��K�y��L�&IqcǍ�X2@��-���W�����+Гy �����镊�@�ܐ4F���A����6�y`๨
�'b�� E"��ϥ��7!DKxw\�&M�������H06\�cD���԰f@��{�����a}H��ڿp( �������}�Z�;�5��2i*[��B�7h����& �k�Y4.���v�X9zv1O�`n>?��y�[�r��_�R�Dh�BK�.mN�2�*�m�B��Y�>@���Ll^��̣f�9�À���p����^xq� @��ܞSX�� ��n� �(.|�qI�3�j�jQ�ղ��<VY��!�9ElлgÀe�K�,ٿ�����fB�U���ο���$3�-B\�U�~��M�;[��g��'a�X���]4��R6�{����ݴ��Xi���ܖ2�X��˺o�H�/�*`����I
�\Ξ�ǒQ��)"7XB��v�KR<���Q*)B�U��ڻ�E1@���tSiq1�*KJ�w=��8RL��0W!�)Mݽ}D	Q��U��*��o~K[;�I�*���D?�\▢�X���u��ƢQ�3%�0%S1r��@�y�Y�ӝw����O�xʥ��6z}�
��O�����-����Ɗ�*�+6	o$̍��%���ѹ���ln�>{>.c�(R���ާD]P�p?�cǳl��O�AQ�t%a2N�$�F���s�1�_��I�&����&��sh ��]����Z"�vl��S�D���gѸq�X"^��: �ȱp5NiU�m���m���Y��,�BV�
t����+�k�ldx۹����2�y��پ�6����ǳ����б�f̚N�{.S9���� 56���^��������D��S&�nn��t�4[w����֏�>�V������g������WB�{߲�nt�����Z5����QP��cS����p��ʓ��yK�4�\�=�ҷ�*>�E�i+vvҤ�m��
�^K�z�\КD{4�˿�<�r���$����\	NL�����j�j��f4%S.���H]ݽlUE�uPQXʸ�J*�~�4���5�֯%�'�{4�-l��ch����jX'P��B�P�v}�f}���%E�|�dJ,�h��J�+���Ρ�gQ]M�M����ڻ:iǎ&ڰi55���l-���)
H���n&á��@ =��R�Bo������A�0���yw��rBmiI��'D3ȅ������ѰA]���M�����E($s���Nw�I�2�����#���:W�ྠ�� �����y�����,�}�_�	@ߵ{篺��.��㏙��E��\r���L�	��F t��Ea�j9��.�,(d�MUp*8�Y�~@/�"���ii��rY�����>��~�����m[v9+�t��BO$�.��cfq�5 :\��r������Хq��LR�zp��q�g�k :���:σq3��n��E`��9���ΕcL)	����
l����t����b�6�g��U�2nQ���
`�_� m:b@0��s��m���_בޓ���ǥ�m����4R��H�R&fO	
����/��x��|�=z�����M�@��M���0}��t퍷R���s�n����/?�a��4fl]|��t��9T7���WTR.���)�ttӺ���+��?��={�i���h��It����)'���¨�	��m���ח�u6s�ڟ����-B/B�8�VY�R*�J��$�'�����:\� tx�2	IfD��"*ʕ#A�X��Ʊߘ��d����;��r+�Y�� �D�Z*Ey�h�U��a@G,rUe�	@S����B������]t��:����!�p�wuv^��� ����X@�F�2H�:�e�25��Ww����5.�ևm9�G����~ ʝ�l]�9��RM.B���xM��5��=̀b� �c�;���f̘!Y�P4� ��ۘ�r��u��$,ttX�8�`��I{6��=�6��[��3`������>
�:6��I�f��|�<>�n,,��a?/{,j�����l��\�\��.PU=����m��W m@����:�&]��^����+/$��r�>U@�Ľ��8���n:����Dhū�п����k�N*
���Q*+��7�9�n��n*-����v����zy�s4c�d����i��Qi�p��TZTL.��;�	�)�ri����ʲW��e/Ӟ�;(X�д���E�w��UR<�@����ǩ��������gVj?|�CI�����U��r}�?���h*�� t,-{�5HKs�	��r�(R���2B��0Vԕo?;���!�ʟ�3�C营��v���H`��w���d@�#��	~�ɑ�VFBF��}l]��f̟.�w�=����������kؾ�W�]�a��75��9�����:�� ��ώů��&�a���n�Sm�9 �.��!�WY-o[�"&�.���mV�Hx!��J�3���Iq
� h�CAڹk��wWqR �����@/d�3������§<���$[yY�j�[.Z���oC���Z�H2�mб�.�	}YeK
r
�����^9c2��)2n�r7�~}\�1�z
4v���2��{���d��k5���G�u��޻7_����?�������J�>���i����$M�>����M�:��� �~�S�ɿ���6�T:J!0�P�ʋ�t�u�ӕ�|�ʇ������^�*]�`]y��>.�h"I�-����A������1pB�J:,?/y�/]D�#�h�UW��s�Re������i�jmi��a��_^1��G�1��^���5�ٵ����l���J�!b�e�u��4�~�%R���F���*������K>��6@4vL{#]��Ee�՛�y .,l�����а��5d����$
k�P��A���J��V+p��%�@�$�* ��t�G#�=Y[S��y]t�)�@7�W8���ݭ��w5�B��nZ t��`����Ex�576r" �p�AM�s]���4#��WcH�{ݶf
��_8��S�
�j��bacp6�)	�k-���%_ܱ��2����0ui]�c��qm�B�< ������jժUB9j:�og���r��k���<f�宀��)��ڑ"��q����k�΅�I>�]��,�
�LyH]��;/�[�~���pY��h�B�P�|�Ô3/��8&�`�p�x�
�c9S��WNp�����Y�!WRX�N0��Ѧ��yĺD�;�NдiS����#�={.'����g��?��;�!a-��'J�RuU97
��ڛhXe5��Ӄ������t�]?����/@<�pW���|�6�]C�@�����E^N��FӰ�*��(�7�z�~��oi��	t�5�PiyE��i��=��ǟ�Gﯢ��&��,��S����I��&RU���5�@�<EE.�C��:�|w�~�����D���Zi�+����V3��K�a�s�k�++)����9!����+�8F�Th�]s��,�V����UP�!� `�k8Fh�\.w���ɺ��g/8���Lq_�����w��۰mﯺ{�/�/^���q��٬��3 ��\� t%�QMT]N
�ڷZ����>��ˊ�J8�[h��^��+��D6�&�i6 6��,��Y��0�+| �7�q��ebTh�+��;w�沵իW�<�]-t7���rW@w�`^@G�c��=�%�D��n���ſ�������7!N�2�2��a�?�{�o�ɝ��u���@����O'�8��I��Ĕ�e��3LH ��>���߯��z��f�c�
�p�����O�Dƥ�VD��o����k��@�P0A� ]��j��۷QډPwO?��}4��	�ફ=�����	-��S���eb�����(B3gE7\3M�6�@��ƛ+����y�Kg��9�P:��/�g~�5��C%�A��jbeaֱ��E�.����u�6�}?����8@�E�:��\#��םw�I#F�R<�RK[��|)�z�mjܻ���(�C	a�����ԫ�c��a�	۠2T9�	�d�V�d-s����-�n4�T���d�M(fD���C��ښ��������ɓ%e���6=�����A�������q��M):�z�2�c�A��{<��Et���>
4Hb���߅i?�3[h����XW�%�ͭ|�#�'Ǥ�<�.9��kt�Cڸ`U��:6�	sf3�+�����|�����sY
s�'����_Y��ރ.��!ӝc���œ�?A���=',G�������K��rW�ԳS���|4�2W��-�|� ���^��6{M>�x 
�v6iR֔�X��r=�J/`�[�:7��P���B���yA}���2\�Ȝv�t�q��~|M�v�aZ��m��C����)�IP�M��Qeq�����t���@�H9�I-|���O����).�Z�G�=�����F��CE�1OF��8�H:n�����5k>��X?-�۫���ϢҲ�m�����W������.��t�ԟ�h"��V&�O���vZ��z�E��Q��s��g	�� �6���?椸��5����K��7VrR^q$���^Q�!�C���c	�3	��g���c��FÏv���2ۋ�<���c^E!j���ȸ��=4�U9b��xmM���.���F���2�z:���;=�777�54�y����R :���ٗ{�2����;j����E���ynTc�}�n�u&����wۅ��r^�jW���������F^�s��l@����ն�mЇ���J,@G5���9�t�/0���M���}�47�F`��ޠA`,|��@G;�� ���-`��#����BNرr��r>eؼc_,�|��k�{���X���+�SU���}���=�3�aSΙ�s5�mw�A'�p*�"Z��5���?@�����T�}T7�����o�e�P�-���vZ�p!Վ��k, $=���������;�(J^�%�\�5o��Ί,�T׎�o�6�=�t��T�'��������vr���8~ON��b�T^9���U�^���%�W"��(`Z�<�ld ��~$��ٗ���n���z����aBP�
۝Qx�R؄� �lD�wUJs�7f�+��6�O5@8c^Y3-�wˀx&�UD�w3$Q$T@6:�bo�Ii���r��s/�簅���������u�jmm����>#4h��Ăc@o��vh�臍���X��=�55�:y6���n��)d�{�jb��蕅I-E ;�7�0bA��{Pw���I�}(�;\���>����Zbu�}�d�ƅQO]�JK땾@W�t4g�} ������~t�y�3��em���
 ��г�@n�B:�^��ʐ��	t��L1�ω6�)����A`��>�R�C�PWʥ j��A	f��G?�iӏW����{A�w豈��P0I�hՎN�����y�R&���^z���$���r+��WP4��'>C��Y��l���f@w3qʸF��b��\3��n��t���Q TN�W}L?�ɽ���5��}��(JS0�&�B�m��	�>,t$��َ4�1��㰅��{~Lc�O������y�-jn@�w�]���ځ��wB�>U�h8M���F��M�֟���5�D\�;Iޕ$>x0 舵s���r	��>s�����#�����[�҅\x�1�v~ 5�92R&S���Ц�}K������U�߻�{�w�i�q�L&���Ȓ[ttd2�����HU:F�ׄF*�O����F���6CT�sG;��������-��ho�l�ڵ����I vhinc@Gf;�G��㍩���<���ךul4g��5���V�D    IDAT�V@��tq�խ�ڀ����W]x܅����	}v��H���0S,t\�o�k�˶�������A@�K������ܯ��zIbr@��8й��e��)E� ]h�*S�=��v���=G�m {��u<�o�cז�z�:>���� %�˺/4��\@�\�����3�{.w��D�}��:�h��wӌ��p���|N?��}�c�6�0-k�2�~��A7~�f���/��aU�����\�v��ߡ����7F��=��S���A�@�¬H$(㤸�Z��>�z���w�À*N�%�֭�)�@"Z?��(EKR��%��π��{1o��rg@NKՇ������w��ԗ
RK['��|9���m΢å�
@�]����.��.wP�>E6<�$�B�cVR �&�M�t�wȒ�P��{u�K�9z�^4�W�MϹ>[�'N��GN@���N�s�;v�ڞL:��"�T��q��T v�)�+����A�q�ė�� <f�NQʥ����~H�r\'�L�8���L(�8!�Is�(�	��Lǥәn%������	g2)�qҸ�7˙���p�G���5� �-�J�\��J%2�L��y:�����8�L&��u�<.&|d2ؚN(���N0�%.�L�9�ӝ�tfkqq���`������� ���nٶ������6l�@~�!��P�������n`jG ��^��L�e`���j��v��T �`�/�n�n���$yI�]��p�9*�ż���`�c�h�8��=�l�����LqC������i�6�rGkD�qn\c�� ω�k����u��^}��R��{�T� �XF5���c�L��zp@���y��8�e9��Y�����/+��t��er��K�/�E��/���t	M�aa��t�7���(D�]�&O��V�)��E�L��}�C���{wS��~
9i�,-��^G]�MV]�(�?�[U=��q�eTU5��{���g^����	���P8����$��Hu ��#4|D��=�s����>�|����)�]��2P)�#�����Gm8s�BL��	�2)
!�ŝ��=���~H�c�SIq���e�j�;Ը{7�З�����U�]��x5���p��8�ق�9��Ya�>3��*X��L��2�����fC���B	���Z�Q5#�.���G�������~��I�( 2}J�@�u���pD
5 9Fq}�r38G,���`�����A(6�L��0�{ʀ���Z,���=�3YC�/Λc�މ�_T0�|1J���o�ko\���mȎ2X��xGR�T*�H�3=�x�!�J�U^^~ߑG�a�}z( z͖m����r٦M��/��E���{h��]��-�pʃΤ
�҄��c%X.w~>�mu�8��7�
F6(�eAZ^�D1����M6�y��u~wU������.w����@�ɉ'�@�>�Z����Jtvw���vbbJN�s3
��,t :�v�+��	%����i�t���eag�S�k�en'�;��{���%���y�����/�j�<��h
�s�f=�n��:��S��'J�v6�#�>F˖-�P�h5�MS'N��N�{:7`i�h�G�5eRI�tޥ4i�4��2�ܢe��#��x�6SN�$�. d�� @2��++��m���>�<**N�����3}�n=)R���s?{���GJ������A��5��/]�4(���;�f�8J"���A�-[�: ��ڃ�.\���9��v�c�B&B�e��%�QK]�����.GR�q�1T�J�/~ײ6f�ˈ�Ů|.�%�1h��H�MQ�$
���`�-o��t!C��Ź��^y��Ufj���3B�Y��V@*�}?��(j���V
dG�ϯ�=���)�#�9�ɱ�RUU��S�N}�X�q�� ��[~���r�P�IZ;�즆�M��B��Z`��a����i�
�Ւr�Ud����@l��Z�Gciє�F��&!?#�Fϩ�1/�]��]��5)���ůIq"���9�D�~ｎ�X�a:%��5��ۧF"�!t�Y-tБ���:�ǲ�s�:S�=�����+�{a@�� d��^j���~�o���7���m��7��}�ݗ�?�,t�n��7�PT�/���;Ȟ3{r��%h��$�sԜs¨��6�'��	s �q
�����7�G��{��HPEI1}��o���PUm-E�)jik�{��wJ&���n�iS��EK��N�?�K���$7 ~7��&(T��h	�p9����`��r�-t�igQEy5�[������>��*.	��S2�Mn0M�Ǌ�(O[��@#�A�����&.�8(���| �Q�@OK����]-�)�j�k%<طX��� u��Z�em'�j�' ����1�����c�ecU&9�)o,z|p��1	I�1I��Y�F*�1����w �D��U&)0*�ב_i��G{�9��Լ�׿b7W4���^���\C���}`��<��0k�}U���;bĈ��O�����3ѡ�5�w6����΍7z�q������nn/�U�����+񆧝��^���y�2`���g�t�Jt+���v��9$��}����4��}m������nz�����I����Y�qu� �7��t��U���g�� Y��,�����ň����zJρє�8P@�g�5��>��`Ⱥ<����J�'��w�?��#ҫ;;7�
�_`�:�s�^v*�q/$�}�@�kt�z�	�����p�������������.�&�VP0PL;v�&$���޻�ش��?����K��r8e� %2i�����c�=B3�O��o���UT��i��7���ۿS{k+����J� ���3���Ϡ���Һ5_�r��o|�N9�T*)FM�������b� ��ӔHuq����f�>��O�Nm-���������G��t	�AL�2�~p��4j�Xʄ�����^Y���{w�@�O��g�[�����֠d�б����9���au�gn�RZ�a7�@�q�RQ����;�\@U�|v2��!nȒ���uN�%�����yL���R:	5��d#�Vy`��D��ki0��E��-��s.� ���-V���;���Њ��Wlm���d��o{ ��Sm���z����磌���������=j˶-����_���t,0Ĉ�{c�^���c �E��X\��M,+˅�T�l�!����rW�o{QZl�߭�%l������6��� ��v�S�\��0N<��fw��r�3�`�ZY�, �i�^A��v�~�i4���s��׮[���u�|"!ݿ2I���V��W:'�E�͸�f��o�<�Q斖��� {n6�Z����$����R�o��&�6����?� /�B���֒}:?��P�H!��>.������s�ǂM�VZ�0�_Xx���sY� ���
�1����P����� M	簪a4n���k�E�7�jF�Q<�䵶{�N��&����r����r���/����]���p"���(�ӧ���ʏ>���O�!����q�)t��Hly9,����t�g�Yg��u�]���g���۷�x��+��s�:����
*)*�ΎnZ��Bf����
�qY,*z�d�fΠ���=�?���K������[o��IqȈ������μ4ea��z)�F�L%R"�8�Ǝ����6v���P(�p7x	�����z^���0�u���;B%�[x���17��0��"c���z�u��;�Vvd��~�o �ē���Ն��y�h��u�������|�K|�Ɲ\n��3jԨ�N��χ��΀�}ۣ�mm�c3#f�����^��Ҧڀ�uƶV�º��e��=WX����<��Ç�9�����S_�00A�(�6���|:n?Xy`�t�^:�	+g�q:�|��TU=�ǁc�J�i��)n��}t@G�6#��3�.�"d��`�0QH�>p@�3L�������� �|�_G����ĳ��\ -�d�M`��^��I����{V�y����t���FY��g��Sq�	� ������F�eރ�O�+��H�
�����qo���;�_~���BK7�t�~��z���a�-۷Ѧ-�������\}��C�4,zy�&�9��cYi���Juss��kjnf��mS�LF�^���_��o� 0��]�`!'�)Vn��{4fb����A＾��|�Mj��@(���P��99N����c��R&���ͷI�\ �����x�1�y,/+�)�k(�Β��?���u�%H��nJ�M/cf9����5Vn�������6��6���ȴ
���I�'A������TX)��M��QC��'_o �|S���l2��=jԨ�>k֬��zwww�����ho�d��ݴu�fv��<ֺ��]]�L�XdC�m�ۓ_�=���P�� :@�
�/�_�I��W���՚5����`���ֹ�6T�Ie�#;��3��㏧�
)t��*)+�5_|I/��x ��|�.[��X&0�Qa�����^~�eﾼ�wr>@�������<'V��� z����C�|�|Y&89T��m��v�A,{C͞�[)�d��=����e�`
Q��e,t--��OP��Ȗ��O<�.�w�>B��� ���q���VӳO?C��F��1q(�7�t#'���7�
=TZZ¬q5#j�7��O��qfM;v]|��4�|�t��b�/{�mpU�1ǉX�Y,���P����I8�R�$ƍ�h :K��1������^���X	btd�3Q�G�gd7�d�'9V��.�UiV2Ǹؑ�`���8��r>�@����'�PV�X�\3%Lu�%����9Bq���|~��K�`>�U��``
�T�cS��>�J�A�爗(��%�~�]o���`��wo��Ge��QU�Ǩ/�NZWW���S�~:��90�Pg�>�o޶��Ύ�K���K۶maK�[�l�J�l@����1���s������5�I �ԛ�L�R^ ���+<�Zf�٤��Բ˷0���Ew'X�ˍ��fƸ�/y�6�[��Y�1.w����]��n ]��!�] �/[��+��(�����6[!@��A���Dg_�����,t �
~e.��PB�l�v�8]o�������!���`H,��o~U���d����!��t��@N	�C��k��i4o�<v������d� ^�Z��r��e�	X!�1�K/��N=�4fHԦD�H��3����O�?�8��j5+eeL�r�e��駟�1i�/O����p��Ph�_�=��3���UR�
� 2\2��E\��:���z�O�@qǡ��>z�w���SKcQ&I!��qt�A��%Y�е�\���?�0$�E��^/[�Y�+��U��2PN�&R�=�5%dAG�\�(����R��Ar	�B������嗶g�//`�=���CAP�^��j�=�`|0�\��������1Q��2��)�u��d2��:zz�6�����럜>}z�P�s�zWW���[7=���u9�n۶�A��+��j�Z�-D���>uA��j�:���-[��~6��1p,dl6�������4�zW�;/�V���|ce���t�{v�4q�D��cs��U�(�Hq}�f-�7�� {��,tlHX:9���@�)
hw{�Qz��W��6�"�Тl��p��ϫ��T)���o��J���[����7��"���A��Ԭ ���{�w�R�?�v�x+����ϵ�jC�F:����#7͜v���
Eز������SO��K�-��?���u�C�7@���ٳ�>�ZX�=}����E-�M�v���{�=Z�f��X�!h�g�̙�
��������h��"�'��ſ{�^Z�����)K2A��7ai#Λay `���wo��#&z��r���m�-�;��a��܄�5+FI�A�--m�%~9@�w�>r��9��Q:&�}Q���5��|^B{�C~�;��#���+�s]�$�e����`�Wِ��Mү?K�����.�;��F���>��� ����#���;�4�/�e���"�Ź��9�VXH��T(X�j:�H���x<�NE����DS,�T\\�fqq񎣏>�}(0gEf_��������[�m~���� t���؈ w��]]��l@W���po9�)��=��8�8����w�ు��#��lq�������y}}��q�ח��Bi�ܹ\k
@��Wd�#����K :��m@׍W�2��o�`��� �_{�5�fR�t�_�.�ƾ.@��o����:�?ށa����L���b x?�qΉ����s�����:Y@�MC ZV%�� @1Tn�z��Q�B�^
X�A�8���Lz���Vv����uc먢��&;��i����@!�2��)/)�=��P�^VQ���x��bQ�rHɠZ[�y�AG -`ۜ�.�����}��B����i�x��ۻ{鵥�ӊWWPW{�7�Lr]��̅�)@ךp[h�9d�����; �����!*--�<v�*����9Z�f+�����B˷$�R�4�BϤtr�P�]� ca1� Ȁ^���	26�/��$�g�Y *m� �
:��hd	@g��+}� ��������d&���5��`0��#b�8��A�1���-�F�A,@���0]k&�	@|�8��X�M�܌�
�L&�J�n�M�S�D"�N��`0�r�@�uK�@�?
E+++�ǉ������Y�u��_wvṫV�:6�	*���_�c�e�t/����V�2� �}� z�S -�aw���`�k�''���2.���u��N�t.� Q6%�>6��'�v2g���RRZʂ�WK�,�r@��MٟC�1�A�]w�utݷ������\}�Z�b�W��������:/�~�� ���^���^3�m�����rst]d����so?k�����#����`UB0�N>�e�nqFJ`�����{���VJ�����B3�9%a�0[�8�78+�E��3��@��X4Jq(��4S���˱8��cJ�V�����
������p��2���:b!��A���f~zOioz*EG}4}���S]�8�;.�u���^c@��� ,�t��`����s  �$�1��L�=��YB< g�ǰa���_�)_��vػ#��������vζ�Qח�3m�[���`�Z�p).*�)oPh7@.�vA����H�J�3IDW�bFx��� hݎ��9�w]�g2��㤓��$�s �N�R �t2p���i7PJ�T��h�adF&��5MI���~.*�,�����$Ͼ{�����ȑ��k4�T��-n �@�{H ��-�����-���B�4�|����nZ*D�z�M�BBݫ���W@��,/S�f:/t�FU/��+e�ݞP-t[	��\� 
'/[�8Xep9�=c.�m@�9�HfS@�Gc[��ŞB!�=!�k���SP�|����!�-�/S��.wۅ����Z �,ߢ/���~+d0�8���=�q r_����nρ\<��0$~).[�U�)�_�Lٲ5]����[���=��|��!4	��X�
.��rl2-�'�D�����<�� �W�u���K�b�I��`h���]&]r�ƤMp,�`+B�,D�G@\�� Ǻ�`���$�q�ǀ^;����@_��+�(�u�0�B'8���#ތ2W 9\��i�Q�7�S�/�m�!�7��w��@.� : �6���X�"��t��mنg1bd>^��G1��W�*X�(J����B�D��U���g�+�ꁂ��������1|��-����٣LڐN3��2ܳ�A�������M	�֟Mڑ}��PU�(#�d<�_�8���ZO����kZځ͢Ԋrmd�Jb�֩����C>M�S:2&�n1ű���F\���3��l]��0�ɼ    IDAT�QG��Y���/_N[6mf7&!L#\m.w 5�����MW^y�dˆBE���Ή7���q����d��(�١�#��`oV[q�sT�g+��m��>�?�������}[�߄�R֠z]�y��̈@Er�*�X˰��3ûZF��#c]������z=r �Wp�ĐT����YN��V+gh�����~�3�7[���BRc�6p�φ��<$?��UY�y���>[�	r\W,|�����K��r5��	�N�����ȞҲS~p��Q˽�Mh��wD���X�w.xdأ��������8��ѕc���q����L�X����P���0(�T���/ �!�ᆌ����a-��È)1 ��p�X�4�H5j$���<o�%7UW������q_m	@G���k���V�BGB��n�0�r�d}\�f��M��m�q =�,@n��sJF�CY5b�n�ޠ��s@�d7�ԯ
輁�5kV�+�� (nc���:;�q~���U!�
8k�~o��m�n����-��0���94�Y���kiL3�}�dP3��P�+8n�,y|M_z{�Rk���C�<�|�EF4�kZ�*\Y�E�L����`/ �ɟ?b�3|�N�µ��ې����������`�L��f���g�UD��@� �;ۮf��Gv���dA�~���U�`e(`�NY��s67�x3yIm��כs?�˺ �;Si)��>{�l���ul�7�w�ˋ��+�^a�{Q$�u� ���F�:���+��ʖ*�xG���ܗ��T
輞CFa4�{͚�N���^��F���G����GRMMuz��ɏ^p��_YY�O�\_e�>&���yۆ�{{z��:߲u3o4,�=��r�)�X�Kپ �_�Iq�k�\X&Y��)�^�S�7��`�V�
%�V=@���R�*��@-OX� ���:ӳ������
[� t���Bd ��8Q�py��e���u�UW!E����e��}y�n@�K!����������6�'�����E���u
`�����`�-{�~>�T�Y�v>�_���Ʋ8'*�pd��i�� �̑��ݰpޮ�Ұ�q/P��X�,p�0��9m͚/�.z��-�,.����Ȋ���]�OlW����VjL�j�"�ٿ&����7��m���3������5ַ�l��og��ܠ��+c����(�9��ī���yMc/ْ�1��9A�]� t���a�/ya-{y�tvQIq��Р�M t)s���
������=���
�˟��/ �	��'(���u��Z�5�7�ϡ�h(���X(����ԩ�������)�z���ѣG���8|����!�[�mD����߰�k�ְ����:����.By�-*0�m9�6�� j��'x��E�)JgF��֯f拥�a�
�n(#"$˚��������_��m�Q�R>L������Ͷn��s���;6. ��a,@GkI �z PB�,w����ISX����:/�:�
6jE�ǳ ��ǣY�F��,]eU�l�g��=`3�T����}���)SV����ZǶ���\<7��N8���=�y��V �x��超��B6�s������$VcIKmܸ�^Y��֮]��R���RnpQl�fݨ˖�7OB.����
������ܿg��9�j�txn���`��I�o�(��6�����<@g���H6{���x��@����܆U��ĸ�0��
�x� �5��rG��%KЋ�BTBk�$�E��ԡ�x�Bφ&�ˢ�L����]5
0�=�!���
ٍ~�g�����������y�>��@^5m��P� ~@��:e�?]5���7C�����3�,�M��?���y,�O?����mjcC55����@�I3��6��'THۀ�߳��ǩ �ͣ��n,,t���
Gl0m�*���G�jٮO3��[�63����`�,\�Gu�~��\����,w���O>��7 ���n�:cID �ㅅ�NT t��X �/]�T:�75[%&����vO��*�	S<��>���S��-}�xg�c^zM�G��
���B��Z-�zJ��!�d�->�:W-E�t�\t1�x����&�@�"��9gX�y�X��g(��aVӵ�HV4��[Zi�c�0�<W�ZM�ʴ��J?{�$C�Xu��~��j�R-�l?wSUQ��}E�����Uȳ����s�Ҧ�k��BMy�{�U1Y����s�Rg��aFTE ��(C��!e����rO	@GH�s2if������գ�Q�c�j�#�.�҈K�0��g]Ls�fF@���(o]Zm�yN�ZB�FUzM�x��Wr��̳�b���ŋ��CII�K��
�p��;�c��)�p�7��g6޴������*����ޮ�D��.�ѣk�荍��p59N31�Ԛ�0g���|�o�)��B�/xT�ۖohW2�%(S���`l��!��2W~������|�[4��D���п��St��1��?��!c�����Lc?��#�X��ʔ���Y�
<~���~F*l�`.V⌦����m@�Z����Ҥ
����e� �.K=�>o�SF3 U�X�
^���I@��b7k�:����/��cǰե�n��%���1���JBa<#���;��R�j�uI�24 �;�HRK�J�v{Ŋ��Ɗ���ۙ�vQ���a��}@�ׯ��y>I6��49qt�4K�G#!4����:RF=��q��X�*�wv�;��Vv4�@)K�s�2IJ���� ��s]Z��AT���d����^z~)��;Z�Iq ���J���ԡЕ�] ������)�l�A������!���n@,tC�[][Cg�u�9�$����}@g��%�	���ӧO������7��+a�tH ����~���s����F�4i"wZjjlf@�b�����Գ��-p=�"�Zc��������Ԛ��q��jbp\�Y�z��e�c�Tf~i��]-~?��O��nT|���||�a����bY��N���7溵k�7o�DMMMܭ�Aٔ����� :�n��V��Ub	F�)u�j���0 ���������HU�^O�˾Wd*!iK���y���Ɣs��]ۻ*�j�#r��kX�~�L9|��nNV8���	���)��B^x!�	|��r�m��S,�ϡ�xw7���CXI�oY �b��E���Y��CZ䖗U�GBE�ǽ�����>z�w�'���ۥs�Ti�9��f�� ����{�zϖ�{Z�D��g���hL ]_Y%Q 	�-އl
~��W�f��N�ˆ�t�!NA�Z1|�E[]�'�tz��j�K�hos+���_�֦fJ��C/)҈a�+bo��p����#�I^v�-f\�	1�i�d�Ai ��a}S��F��3�:�CA�����k`Âϗb�;��ស>}*Տ�>u���z�U7�n�F"�\��;=��lm�����Y �e�� Μ9�F���֖6����.Dmzbz4*Y�~+[��V�z�f�J����d΀X���6�Z.#��t�_K����ݮ��T��MZh�:>pVc��ː� ���Q�G�bm�����}<�� L�Fiq1'��g = �;���.w-Yiio��@G2��߃���}tdcV�LKW���**ؕimu+8��Ę�u��b�9��>̮CQȤ�3$�Um�h��C==}�?`�����o ܌�Yiij�HHx|JHeX�tlxF�֜���nqs0��U!���Vu*���;iێ����8��&q���QM�����a^S���JLқZ�ڳ����>�G}���mmR���(������\[�4sIS�v��*o��;H�Toйu�
�`d�ub��ch��Ш��Wl^
ܣd��K�����X3�%P�&L1fz�k�V�(�3g:ǂ�f1>	�@1�s�����З���V��s���u�K	*.QmM�qs#<b��h�2c�k��6T�#`�#���|e=hҒ��W<F`�DJY�0V<������z<*���w^��8�][C�fL�q��m�g�����oXx��u|}�;�����ræ����b@_�x���&�%�݆�fjjl��p�E_LJy̦T�D ��vu7��d?���KE������ϳ�*��զ'}�(u�tr�D]�:^4�(�mHXM�Z��؍��LW5�A Q\*�Qߺ/�2!b� �DT\�-c��{�E-�Y ��܊�|�ЮÖ�o}��T�BX��� ���3����� �91�K����;���a�bl8>�3%%�}B�u��So_7�[���@$��P&�`W5�K�ܣ���m��Ǩ����HI��]�5�����r�:B2~����ǻ)x����v8W�蚉P
�l�iy=B_4D=S/���JliI�����|0�ZEc������0R��.[A���1ڹm+�N�"A!cI+}'��&���ŀ�ƢU��W��_�m�>n�~��;Ԥ ���X7{��[�
�>��H?��?�_�p����Vb.�`˜�}�=.K�Ⲣ��e���(+ V� +&�-f4lq:�9����JU��/��=-�x�bz�7����z���P�' ]+@,�J����W������l~�D�^|��(��I�f�c���%�G{�:������elؕ���;�]"�O�nc��	���o�:c�=���À�������!蛷lx�����իWӋ/��«~�x��e��	w1,P;�EΙ�dX?�֥c���,�3q�|nF��w+�c�k����_#%�!D��s_��ϫ-z�Ӵ��}n�sq��h,��&�4.w$�	����׮��V�\�1t���8��C�$���b�ޞ,��%�[]���S��Z;~@W���a�B��\��Ϟ�� PŜ*G�f�k����>d`ܒ��<+ƍ�1،D/�e=l�B�R��\^VN��m��A���5Lf���#=��y�~p7�
g�#��ܸϢ�t�bQ.��\cLP��<w''����\c��_oT�Ӄ��������N$����E?��O��WSw'���Z��c�%���"JD#+���'�(v�TI��t���y�rk��Rċ�i
��&���o��C�q#g���	J�C�!�qwxAT�B6S�1+Z�N� ��JǄ�z���~\d�k�_QDҜ}ozwo���i����+����b�>
9V<����gx�N���&�.
dp��� ����C�/��<o$���H���|�\�,y)���P$(ʰFiJ&�x�J��}����3����W���À�{����~nǯ��w����a�vl�����z ��%��k�ꤓP�X��*@������w�ܓI�ד��8ix@��S�m��s��T����h�ȲU W�P�p �ChQ��k6nօ,V�( ��%�w�*�{}�M� ��s$�=�'Y�l���m޼���%��	 �T� Vv�� ~  �c�<*�t]X�:b�ljX�I�nn4z`,��@H�3M&�s�@i�N��� Ch�}��j�$��Y*�<�C�  ��c�UV�;�ޜ������6���7Z��b��u���EL��s�#��̜9���GL���|>A��Jƙݭ��E,kʶ��}0@��{�p����5�x;���b��B7<����GDܶ�B�|�&���~N��	�!8A*�q�kY�_
�Uq�g�j���
�
��(���HZ��5��s#\"��`@hQA<ÊS
t�1&ꁒ���{P�ј�N����`l� ,VUn�����tQt�P` �7�tв�_��__A�B渃]�*��{	��kZu�2��UY!���z��]���(,�&=���Ћ��)��=�C2�.[�:σ�t*ʀ>fb���5m�1c��W]u��h�����t	@ߺ}�ϻ��n����K,��N��O�I��2��]�g������4;�&`�B��������6h����nX�_�wlE@]��fӟ.��L�L����@�M������y�Ǝ���<It��<n��9�������6�]�Iq�~Ƽ���C��zl�;�GRܕW^�`�����������m���<�Z�f%��w��X?�;Hm,X�T�Q��o� VY�e]SZ�����@P�U-�=�uV5vy�:[�&�v�t�9s�,����u�X#�dWG/�{ｴt�R>?8�`�+���CBz�����7�Jol�VD8`�:����[�p��u���Gr�	zH�C)��}�����l ��q�3f��)52B:8v��'r�1X�KII�d�����c�=F�vn�0�Q�p������@��2��Ѝ˧,+�ۖ�>o��G]$�\��2�w8!5 �}1������ ��rB�=n֯R��Q�\����}��_=H��$���.���{x��h��td���[hD�h����������A�.
G�u���p����(��rE�J�ё#�9���K5Ӣ��� t�:0iQ����cБ���+��|@�s6H���@�X�iƌi�ӦM�k����=�
���!�۶m�YwO�ͫV��E/��. XJ��7��c��S�io���.����eVN�"�H[�=7����Ql������
�]�tډn
��F�G����v9�HV}�����u�
��:v���e
˓��ʤ�ڦu�r`�<P��B71f$űk�$ŕ�@��=�``P@GL���4s��M�az$P6M#n��F������)��>����������8	M�e1������ nq���
�w��ք(�|�m��̤�H&��'�=%G���|���Dܮ�&ۗ�uψ{:�=������=&���!OЊ�+�η���jF�����B'�0������<�I��8N�R��܀d��x(�!j�-~����SO�d�pq�Xp� 54��O=K/��"uwvP�`�{G)���ZB��X��q'����g�[a.�_%� ���~�t_��-}�S���~�z��%�$΁�� /��*P���0�+���d^�H0dr3\���=i���.ox�^��� ?,t���u�ٗ���6Z�t	�Z�{jB� {H�����'���H�3ƉX�R1�ײ8���l[r|���8\&0Lp�+�sN<�ڷ�|�}�С�S �q�Xma���4M�6��n������t���<=�#)n�֍��������{�^X����S��c�>�jǌf+�����nӫ��7o���mk��Ҙ�Ϊ
?������9ѻ�s�kTb�	�k���1�lV��D�dec�@9��� �]��zg$���@�l��2&�ذn}�#T������B�΍�C.uvw����-t���ba���9��s��q�
�hF���; ���.�3��..�ϟ��Ӵp�B��\s-�F��`Y�~�� B	��������k�6,b�3΁w���ʊ^x��ϘA���4a��#<W��}��_Ң��B?l���ɠZ@ �1�����v ����8=��#��4�ΙC�_~9�r�	,�{{zX����R2�$Ľ9!�r�|�jg��ѺS_�d�ˍV��>-Z��&O�F��~;UU���w�n�G~�$-[�
%bQ�L:�����#�1%^�\�/�{�)�r��%�/$É���U0��Ě�.Y����(��,v�t/Ԟ�$N]�%Ea����)�7KUD���9:���ɶF6`��X9�1t����n% zW�v�m�W��L~�>{��qIŐ ����������΁��	������c�ڨa�{K�������������n�L������f`�����X�4:�	S܌��hܸq�3fL���+��pw����_��C�7m��������,��=�.U�$CAU]K�'�B���/m��i��͟��F�����\�o6��;�~]�\u�(��r�� �5    IDAT�{�=�c}�C2��L'�8*Đ���B끵���J4LP�#�cgπ����7*\����k׉�}��b:_�
�;��X�C��+\�F��=%��-t�C!�:�k��n�o|�1�{HR�{���b���o��:�����-��?��c�h~%�����/>_�s��4�]�<�s���y�V����s��ۿ�u�xV�p1utu���=H/���� �Y��I�\����9i"�������c�nIyu����}����3}���²�t�M@����5�Dc��{�)7���{71��"HQ� ���t��uv���s���|;,�{s�����ۦ|�}�s�s��#�<�W_yE���A����>�0���׭@�����-��Fp��\����l[�Yzb)a��e��_��������kQѱ�����gb⤩x��ױ�jR񰔦<�|�2h�]�K�u�D�?�m-Е-�[����4��(�3�Lb��!��&Sbɍ��yO�
�@Z�kƌ�UrR��` �D�@Nn 񈉒��>�s��[�#R;M����V�֨%��5lؾ8�Цm;􍛫п�f��j���46�ό�Ď	o�:1Zvp2�5B�C��غ�cD�^c��m���	��gJl
��|��X���9f�{DɅ$#��Z\ �C��;v��۷��'�x���mT�����+� �իW�����5�7'�!�-���%ѭgh�%#'��Y��FP���ƻ#b��okQ\��u&�ޝ ���)j�o��`�}�|nnnֆ�����qg��)N~�nZ�����ڳ��g�I�8�x�2�����CP����+��0�2Y)w3e�k]�_�;�����^SW+5t�F�lߒ��uv�:���10�lD3�Wc�Y����.��G-)w^��yoY���3�~�G��_�$s�n�zCe�>}%B�ջ�8�ш)10�CBI3&"-2����_���D�N�}��3<x
G�����w&�v I�̶�e:($��uI1n��I�3��iGp߃`껓%��Ҿ����~ʯ�۸a�dx/��*l%�E�$u1�ϹۦTC�pv}��ǖ������x�p���u/#1��J �i�"5�u�k�JF�>x�I9~S�
��>���D0d�u�����3xXQ�a6nǮ]"g�z/#F�HJ�<B���i��J/��r�!�$���/��ls�}s���4�o&%�(Tn m[���Z䀜��wJ��P��#e���=1΀�1ǅ)���!ř���h[Z��P�T��30�<$�����T_g3L	qX�Z-5(0�yN�_m��L��
����S��0���.>�D�zu�)}��#i��3at:t0)�N�;l�ݻυ'�t�;?d=������t��++����P?�&��DZҗl[9�y���lԡ�B����:�J&�a��)nt�n�����%��?�V�1�|7=��_�#>>��C�`l���'�YG�A��(���CH��$$+X�N�ei��1�V����Nt$i��:�o�
SC__�^J�hM�cέ /�z��ɥ�L��ԓ�P1B�U[#)w*Y�Ɛ�Z��ӈ�1J�En/j�y����6E#�\r�%��fM[S�L���x�14��O<^��ĠA7z?�p�E Ԛ��6�L%c$ϯ<W��i��r��7�W^}�8B��G"�G}\"t���H�E@t{���w!��}�
�淿N��ﱳ�O<��M6,��6��h_��G�A�޽n
IY����}����)܄�`v�2��5��DǅG��nݺ�r�:<��Өh��\s�U�7ў�-iq��v���׮Y�|�s����"�,cp����dŤ��[~�:���s)ǁ��ic�{���+�Gu�8�tr�w�kf���X]�s��
k׮��|����^�QWW#r��jv�ii��m�y����t���#����r�*!>���R�nU(�:��ڰ�G�i����������Y@}�H,� I��<̢ܸpZ[�2�>ُ.�ŭ��o�ڊg��E����y%�FG�5t�V�f�����結��	i�Q��l�B�w�Q���&�1J��4��N�aY������Lc���i�e	�S�x�:	˽�}YU�>}�?���'�c���w�!W���w��QXY�����Ƌ��z���N�V�GJn2�$���W7�D���s��i�UAN�g2Zђ�x�tc�A��b�4�� g���>LתU@F[��������#7�g"�H�3}Mz����j���Ǔ��T@Wr�A�� ���ȇ���)���LM75��%	���Ѝ�&���t�����f�x�qQ�c�.��*o��x�:�[S�{��1F���.�@R��@&��H�J���W�I��߷�D��gd}�q���1cP\T����y�XܤD��棦�FdQI����h���^��]}�5�ի���3�nhl>�ɓ�Ƚ
z8�,&��r��4����\V�N ��xI���Ϛ)��s�
��i+\��G���%S����R���Z'����y�q@hh��Љa恌v>��Y�u�ة���*���Y �����Ǘs��{�����pۚ?#tC�2mn�X����%:L�3477z�w�ȳ�X�aMW;�] ̔��R�`۠:�|�#ZSS�O>�/��%l\�Q��k�n�VF�%��7^ôi�$+F�
���]�()�]���9O }��)x���0`�@�z��څ%�ⱈ���	�z�5�3)�_����&�;U����&�tp�"i���-��b6B�&Y��P�!m�S����9���]-h�P%������'�ϡ�!�#�h�l,B�Èd1�y���3>|�?������W��S@g�N�� �-���9���0�����+�o�����ׯ�ccc�s����	<��N��� 4h�2�����uғ�w)�?b4�%e�zY���|&�Fz7��|Ow�F]���+���JG@b�K嶂�BI�E�1��D$'�ilfcg��5�j � Q6�g�������� ��U2�t]�z����4��F3��O�d	�K�\��	Ho@���}L�;a#r�^HKv�u�y�0̣%�8�#��k��>��3�5t#�eJ/����h 9�llj��s�m��S-�����kVhF���t�\KGu>��#t��7� ב���L@g����CO��XT�YR�������PEŭp�Ϳqְ%���_���@�:{���{u�9Y��_T:��N�9RW:)��}���ǣ�++��y띷�[���"Uz�n�Й	
���Y_J�b��u�B�c<IqV����Tr�m�eW�����	���@���ϓY�#�:R�9�/ݮF�{���)���,�'N|G&2����ѹs��"X�j~�A��$�Q<����"L��B�ℓ����g_��UN:�(i]�D"��_��1�8U��)��b�J���W��3M���<�2���ߝ���2]r)�[��!ź%�N��P�	>��sJۖ�S�5�kD�bg��Q���mοI�33�Ap�a0�Ā�*�"�[��:�*`d2�"�#DQ�,�v��u�2��N�:J6��}�-}��9邏Μ�OE��?�����u����ۼy�666^>o�</� ���c	5D '�RDg��ī$A�Ѻ���!������&����1x�#���e�5su��&Ҵ��O膓Ԙ�9�$ݕ�cj�Lj�����9��5�ipTu��R�z|
��UfD(,��RtӮe#�ի$�ްn�l�pc�FFP%45z��xL�$�e ݇�@�jc�=N
�8��3r3�a�ݞ��T����;y�����9��xo����tҰ4�rd��%��<��e]���|dRkό���hD ��7ߔ���_�R���g����M7�F���L[o�ށ?�}>����ST3�J�u�y<L��s�r��p���54��'��[o���@�����AIq��A��e&�v�=���4�������+��.�8���L�RD���q�5W�C��&�c����ᡇ��M� � :ܕ5.=ٲ�"�s�]|��%���9�:�-E�H��@1$jp/32%��<�~����r�N�h�'bf�!��/��@I'N�frEz�!l��"��l�nW�
W^u9Ǝ��x
�-�cO>���FHi�� ̊Qq���FxBt���2%|I,`�Ux��g%�CG,e��}��m ����}���)�®�F�{�j?��~�C�}^':��=n�@9���;�_��Mt��gL���E�qq)?m�Sf�)�X������9�>7��	�tx+ڗ��~�/�s�����{@߼ysnUU�o��7o���I�H�Q��^8��,8�(0���DŅ�5/�;�S���"։g��W��&q}��f��?��:�鴙�|�>���΍Bϙ��2[�4�f�aw@w�:�}�e�k�@�ϋ�+WH��~�t�����c�E��cJ�s/8�j�3:2���#�J��Shv ��zv�����Dё��S�<7��v� :�՘!`ڟ��^�W^ye��о�;��
 �.*�g��Q������v�%5���n�Ȝ�����J����kUѾ�D|�;'��Y��V�H���ӀN#���)ll鑨�o�r�sq�on�رcO!��P���9͊���{bܘ�2�Qۋ��~+++���$�tN�b���n���������z�1�ma��;t8���*~��#���ϒk��j�˨��
˰.l֝u���`�`؁@ε缏-�f����+qT�_n���9�9O�g��o���&M��
YǾ �x
L�j��s���A�[TT��@��R���x㍷��B
Q�kW�o����p,�ys��������-��E�y2��ٳ��W��~�uef��#F�uq���S�L�O<�];���t�t�LF�
1�׮߀��O3zC��[:��uɣX���V>ֹ?���g~�{OK��D*�m�M��4Eqؤ�����%;qM;*��甞~���&��ǃ�;����t�f��+�\���g�������ڵ릆��k�ϟ�C@g1�y�a �$qj�OϞ����9�`�2��?!��Pi������НQGKuA>�	�Tmi������{\k�D�0ҵе��>v�4f2F�bw���|�Z�>��Xh����ef|*�Q ��P�L�z�r}�T@�!'���M��{��)w��UZWY�N��:&-�ܛ����8ȡyy8묳Йy��:��ꩧġ�ۻ���U˖��m[�Fj�ݺtEY�v����!+��A&�����Ji���/�@�w��a�ܹx��Wd���:!`
�1�@����������<>�b1�.֤Ys���C@��M7c���Ҷ�����C���5�w�}����U� �=Am݆ft
��ؾK�,���d��Q�>�1qһx��1n����+$� �؜� �~"QkՖM��&�5t>��}J�����dP�-[�P0oi��m7ץ(���,��ĕW^)\�lY%[��E��Z?�[��Q��F�DNN��}�7�z]��W]uڷ�(ϣ��sg���GǼo�y�E���	1j,ܾ ��b�|����e/�v�б}�7�«/����xU��~$���N<�d��?ܮ 8]��O��Ɩ�q'���:���#I�O��� :9,�Mt����e'S�3d�f�ǒ_��/~O�RS�\72pIF�IlJ!K �5���7�m��"ו���Т�!b��r-,�W�����O<��d�~�?�
��G�T�?w��������~�m��*4J����"��D<��6�n!�0�ڮ�<m츠iHYWg��Ů ��ӭb�M��5O�m3SO����v��%�竛D]��xSӿ���x%��nf��Q믧����Npbʙ�N P@g
��.���������A�)L7]�T-�3B'��p����L���UYmkz�����ikfd�O�C��GR�e䭽n쬩�3O=%���}�I�r�
�߽z��wa^>6o�$)l��رcPѡ�8r ؏ϔ'�='�1����-�ѽ;e�̆&)�������X�y����N�*i�/@D2#/9��=͌�\�]b~�����O�!�et��˶SV���1qM�QSW'���%�}��
P��#�+�A99b�_x����ki@��+0 #k���<� �lޘtё�S���^S�������N�ܨ&�a0J�"��6�pt�^|�%J��k���Qz87/7�f�j�Z�+V,ð}����/GEE��D"Q�y��K:/b�oЩ}.�l�9>��K<���0h� �r�/�!5��g��+/��p�tP�N�/�?�{
�[��)��g}&]U7����)�3��Y'mƴi�5����Im�9M��&Se&:�H�t+�Է*S*���0ڍ#�,x�D2�"N�C���d>�)�WR��~��ņ�㗒�g ���W��W�tҙ�������f?@�~��7W����,\�m��w&�|j����5zQ�9ݖ�Q���/3����H(������G�׾��dKDk:�u��I#Z�%q9�c<�h¤e5gZ�)���F1D�>��Hܤ�5rһ��W�=�$#�C;L ]�\�}ђ����O��`���U.�� ]硻�>�z(˝�.)]�e��;�S����Z�q��:R��κ�1�kz�}^ĤW:�G~X����e@O�QXcʝuԚ�;$��k�N��$M�1�L��S��1cF�:!xlش^"௾��1������R/�BMҶ�>�x4�=�'$k@g�S�|n�7��F���pT�5�F�7зWOt�x���3��5`�B �>ufx����E�gRG�˓s��ĉ��o��+�����"J�	n��� ��M$+�����BF�r7β'�V�,��|W�]���(�-ME|x>�ّLH�}ֹ�H٬��A�,�pϐ�]Ҧ8=J��Nbiaa���\��z���
�yϴs8��
�\�̇�2y^}��q\q���g�HI��ٗ������#F�#�4� �ߑ����(R������`\4�����8f~��d *W�D~^�dXJ/d�'5�/��JJQ�Ԅ��O��I�!]�[����1�W���u#*rM� G��!���-�c�H��p'�e�s�@��e��UeH^*��	��d >3�� ��Lʞ�׿��P�޽n9�đ��\=���?�
� �5w��+C7�X��x�;��|�Ra�*��� ^:��P����$a�ƀ_Uy�,r(	T$�I��F;kE{�#���0��x$�����a0�Q|�r�{%�d� �g��U�Q̎p�}��1�g���?�I�rs$:cD������3�`GPoj��PI{Δ;��I��(�M�1�nێ�{Lj�L�Sa#�l8=�4�k��C���T�9֑����#mi4\�dBX�M!���;���cԈ�����Ła�#����]��@�?�@���oʞ���s�5��;����9bh�oڈ1c����e�����~lݱ<���t�b	|���W"f<��������F��>z��J�+�|�Ui��ҹ#�&k��6>��ؾS }��������zwc�����b���@9ܲ�v2�唩S��k.��
��w|��������c��U"C��B����9a&�)���L�W���^tL3�{sm�#Ē�df}cȴvy���p��E�ޫ7Ca���|CJ�z�\��PZ����1�l�c����ǈa�p��g��_]C6n���'�:�Σ�zL|�e̝7�w<9�X$Rn|���x���0~�~�a��)@<��SO��W^}ӎ�u��mB2�$�y�ig`��ah�1}�L<���X�r|^ �MI�ݕb�������Ä	���mv64`� �4,Y�H��ȝ��L	��dE�Y��a�Ѵ�E��m�5�6`$��9u�%�5�����iU�xGu@����fC>�%������A�=쐣�...���!�?�R&����)�� �ꪮ6��4nw����������L}D].�����ǿ=��<�ΝsIcc�V�\QB+IK��I    IDATJ� )�d�z��=�;#1S{�IDcIcN@��W��>R\6�kJ��C�Y7�D�$H�a.l��FS���4]�t'���34P�x�;v0��9�}�p,Y�3��@Z	��u����Q��/�׆��tWq�����=��D�L�� ]�+p�����9[ ��j5:&t�eΘ6]����u�R�>?*��%a�kڹcn�y�A�":uu�`��i3�J�Dm}#���^w�v�����B�������p�xɁ��d�ǚ�9�
^�����݌���z/����O=�w&�%B$�G��1ǘȐ��!�H�z��׫Gwɸp{����r�X��܀*⌃�#g�����&bĈ����KQT���vO���>�=�֮Z)���<�Zk'��>��'@-c3�����}�7N@W���ٖu)έ^�@��~��i��ѣ���k�C�>}����s�̙3��>d���~��Q���<9��z޷���۰w�޸t���Κ:���KQd<��CP�*�ZTU�Ǥ��`�a#1x�hx��2���������D~�ј���^�m�t��Ǒ�ls-���g�}�����f~�9���[S)ב�2$ƹS�a[@>M��mKQ
�r�Y�
������	�Jv�5��d_���H�9k��3�n�s�~D3%@��jw�6G?Sm�r���=$���7���.��РA��~ء�z�54��n���v�Ѩ˛24z�T*��?�v�k|�]������%З�E��Q:����r�b|���r�݉�ۛH$�nw�Z����K$�W !�M&�st�|��˛r���d��J�<�;y<����{Q�"��T���O��d2����R)o2���2_S�T���2I;���T*%��W�&H�ݮ�d2�>�/�x+;v��h��$ }���44�߲|��tz�\XRC�Z�٩�L�T&V����|3UK&�54dTܲ�����&�e�Ҍ���45XҞ�2���i \��u@a����!��$-an�� �@��=�� �N���Q��D�K��tI�3�H�O� ���(�3�mk��M�ٺU-��8!IK�i��t^C����m!B�q�	rg�}V�y���a�M��Tj�S��{yi;�**D��]$EM'�;��ט_���$�1�%xo�NA�X�j96n� �
2ڇ����ݙ�v��y��]�������bL��$�sX
�iI?�X�N���]�w�o��v�6��Gƻ�B<ք3N9�s��
v��֪j��=��8�t
IԖp�ng֬Y����[Ii[�5`�Jy�����/��K�I�&�����9���C�
�{ 	��-��D5�6�H����gtk�Ij�I*#�Ҏ%YЯ��z�g9��g������C=T��|���� B�g�^,_���z��\2a�Wt�����⫯c�%��)�����N4��ϖ��QX�ť�H���x�Wq����m�0υ��oM��d���&��p��7�^8���D2��g���{B ��t�X'ر|3���6m%��]��q�0RO��3�,�t����L�UAܔ�����Np�2^�Ϯ?���uygfE�4(,�#���2#Ư]�v�ϐ�rs�6�]��T�4 ��K�!f�����l�*M�)12����dH�l~o�O�|>�y� 5� ��?��	��|� ʼ���y<��W�!����\v��39Ќ/"�|��?�����J&�Ǯ��������8�H$��x<�H$����d2�e~~�_���s��W?@�wvCC�m+V�(#����N#�=���r��&H�\l1}���FT����Jg����)�)PN��0dg;�[|?�2�M��W��T;����z���v2}�Δ;����G�^8��#ѱk�5 ����t�
|4s��"#tI���	�<t��[t��Ł��*%�e; D@��Bic��r��r:0$�����,����������òW���hW&�^={H�b���@�/2�(����3K�̊�˰v�:�6�w���k�C�.]Ep���L��{�}2/Z��ɔ��	�r����������A���Zm("��N��SN�眉�֭Q����`y�2̇`̙�<������h����-������9���^xAz���\2A�_�>����7w�<<��t���t7�2�!fX�?г��3��u��^�%�H�B�s�N�~���_����K�ŗ^��)�UA!���")'����z��?�n�k+��/w�	�۵�e�0#AǨ}�%L�1�?N8�h��T������ߛ�H4�y��c���ǌ�_�� �eI�G#�Rww'���a��q����С}W$�L�-ʁ֮@w����~f ��BB�E],)wF�L����%���:3�I��9�j�Q�[��-'W��)�%�)���zT%:ȫP�"mk� C��u����m]�]�وͨ���5S��n"�����Ь�f-��l�������{U�T{��	�^ L��k��:��y��e�4'V��������D�K�����P�*�HT��c���{��f��$ ��o����}�ʕ�TS6�x�鈡�Z�F���	
�N5�m���켑�]�1VvX�����it"@b�7���r��qL4�m(�5���f�+�3�W���w��]��D0�:�s��U�5�#l���(�Ѩ�m?z�kS����Q�o�e��}�m���2ӯ(\������WT&Q�+k'e��9�=H�5t��)J.�ɸ��u���/wS�`6�� H3|�0�Q��}G��hZ9l�%>H���m<�>��$�q~ �5ч�34ݶ&-�� ��܅{�{ �?]R�4�����ܭF9�^�p��-�6�$ٹ���=�8&�=��ǎ�٧����b$�$�5�c�+0��6��e�u�PS+��+h%��</f2�,���|0s&�4\<e:�b�q:�I��|� :k�$�	���a+��LBK�N� Y���q[�H�=�uE��C꿬�Z�:3%Z9r4.���գ�D�/�����

�D��*�{uꈓO�5�3�`�]�?�y;:UT����FIIl߱�>���^����8
�~�Τ�P�.H�\�d	�N��1��������G8���{x�簽z
8����~}�q8�Wg����PBHuO<�6o\o�:����p^}B"�/� )�ڦ�D�L�nX�V��/���i1�����E���uT�Pt`�kY���2�δ9��6%��+`+&_���!02��tw�~��^��)smi8M�����p:xjƿ�� ��IpZuX��k�aT[�Rа�@"��6�?g?_������Y����y�Z�#��5�����J�ZrrMnn��C����re��Z ���ϝ;���P�m�V�*��5�Ӌ%=n�������[k�;���I�k-I�ᲆ����~�Ş��R9=/�as���3f�g ={A���Ii�Vy�H��{��#�p��0�}^,^�TX�۫�
��,���z�"dۉ�:�*4�8�*]��j��f�.�e#��L��۔�:<���✀. ��;o�S4��������ɐ����I�3w��.��G��ߓ���%N�;��fFh�ʕ�>ƶ5��ɽ�x�e�.������E�N�Ll�3�˼9�9�m���]2�����x��W���0l� \p޹���{�.��[�n��֭�d)�nɚf;[�I�)$���������	f>�9�~���	_�����0�3g�<<��CX�j5�4�,�X��Jk𴆮�}UP�=�5��*[Z%��6�mR%��B��-mvW^{JK��y�>������O��N�
̈�?n~q���;`�ss1o�|�w���]z1ڶi�]5�x���1y������'s8ƌ���$��1^�x1&Oz���董��f"�Üy��̳Ò��[P��B���p�i�W��p{�";˶nڰ~�^�k�6��/���6��G!�2Ӧ�2M�3�h���;��ג���r��m
Z��I�%Pk�̹ ZW0�����^S�j�4RT�O6�*��}�	���9>�h�����h;��%�x����=E��:C���+����~�l��^�ο;��cqf������Y�>�����o����i�ɽ��?���m���g54�߾z��f)w�pR��xu�Cf�e$Zd0�)o�!e_�=��$�d/scUѭy��4pJFх`�Ϥ���vs;�]{�B��ME��4S�Bt�z�x�2a�o�j ��Y����)E#a�.2�:����I����!&���:�@@W�Ȯ���2�.�L�g����y�rHr�-��믿FY�21dd�S��[�����t?�=��nÌ$$u/��I$�����AG���4���-i�k��Z =�NJ�}S�6�s����L��� ����a~��)���z��Gv�"Q<��Cx���a��Cq鄋D2�n�.!�y9H��3�+��sm��0a��#FR�?�H�Ҡs
ޛ�2Y�^�e�l�N]��`Vċy��1��Йj�3B`�̈$�E�Dw�}�/�Mu!��j��O�&=�'��:�j'�?�b��7@��\c�f����n]��3�Wg<� t��n_.<��ܫ�}Tj�]x!rs�Q[_�g��&�7E�c~����I'�BT��7�	�\��s��+/�������������&|5�k�\�H�Ц(�>�z�W���L�����{SE��z�6ӶF�a�~���Ѻ�m�2,w[���j���yn]m��EJ<���u�mn����\KN���5ZV�A�&Թg�=5���8��, o.򜑚m	k� ��j���U��-e��9�pK���Z���K���p�S�s"�Hu0�{�ȑ#r�\ƃ���'�gyV����իWW8#t�|Zߨ��R���8s1h�
��X�7!ۀi�x&2o>�DӼ�ڡ�M������ޙ������N�碒�һ��k��e������PR�UƆF"���z9.*N�kf�$Z�����X4Ec��c��#���&��C ]�I7�5Z*����t����>~��\�[o�_Ϟ�����
G@gsII�4��P�dL ��1�$7b&�
�#Ѵ�� �*g��y�d?��7������S��ņ�Ui@��͕1�􄝒�(R�{HJ?�o�Ռ_���]��x��п��V�:t.��<9F:~�9^���86�A"o
�p�J�ehUT$�Wj@��FC�I�:Iq�7�M��n���+�D���L5�;��q���cՊfB�Bb�b�Ѝ�QwcIН��k��}T��ɦP���[X�du�xQ�j��m/���p���Ѻm����zܴq��+�h<GJ&��A�j������z���ѭs'\q���ر3v�@镗�!*��]q�<�PQd�|��s�^?�����@�|�I��O0C�E�ENL�p=�(���J '�/��U۪��ko᭷'J�w�ښz
C�*5t:S�T��1���CZC'��ΐձ��L��LG�̒Y{��S��h0���#s�F�tՅ��.3d�2 ����������ר�R�uFx\�Z�l�<g���ON�%�Ύ��VPu����t ���:m�f��~-}��[��k�	�k�Ph���f���ӿ�\~*:k�;vV߶nݺ
�`mS=�����f_��9�F��꼠���B
^"���\�΋�Mƍ�~n]���R�i+aJ�zݶ��#�����5)���q�i�IS�I�����_fJS1�����l�JIU��	D4���M*������q�QGˌrW  ,���W�`�-���R�tmf�~87]�۶��[���-�7R�9AqDn��V̝=�0ڻ���ѣ%��J���H&4��9�������"IQ�`UW���5��,((D]m�d/���V$a{�ꁳ�;�����1Kk�m�]w߃/>��L��x����.�e�x/9���;nCKPe��ac��~L�>.���}:�:�hy���7�Vy���pEI�2����^|/R>��!��]h�E���'�೙�ŧ�����%�](�<&
3qܜ�q���b����0x��I����|��D�dOF���k��]�]�or�ݬ���q<&:��Ԏ�rѺmu��8��z�.7��ӧM!J���^n>/]�������Sz�8��3E�uWm=n��^L��>r~��a����]�}�9�s��+��AU�7�x��/�=F��NR��'��HL����H���G^n!�o܌wޝ,��$Qʔ=/I�d�ؙEiuH�J!Y��aT�߀S�@��ò��r������a�.�>~�Γ�'7��1tp�,�0��u̠�`��iT�#m�R�,��ܖ"��`%��ݛ:#2�R޴��I#%�݅�}z6 �	0u�99R��{K�5{��l�lG"�<kwՑ�n,�a��=��<.�_�	P
5m
��))i�Ȱa�6�����;m���;֭[��	�ʴ����5B�Q�G��.ً�i��#�l�]��d
LHJydY��
?G��e��#F�AA��	y3����6��L��o�"�^�3dN8�a�k�9�v��u�6}����e�x������^i,&L����ϤC	�J�>t��0��A�8"t9O-hە˔/�/��	ȍ7V>�C�N��!�vw�~����:tD�>}0|��܉��)_���'���X߹C~���)w��ڠ��ۄx3��/��]�9_��^}zb¥ЫWOM�}XU�w��.���(���%)ek�x�Ԃ���%s`�[��n�����cxr�w�x�rƩ(,j%�/�#ϗ�\�.F��|�*	�����7�z_
�Ŧ�:����c	|6�CL~�5�4W\0��KdЍ��}|��lI��������~�٤ۚ���4,����� �)v�_�4���	]R�n�i�!i�Jw={���G�Q�Ơu�b��8	#�D�h�GX�s�Y��?�BT��nۂ#:�_s�dl�,[��}�>�T2G� y�i�;�c0d�H!)RYoһocȀ8�SEY��
�ǄA4F�ٞh�,]�Y�>�_}%��f����5��t@�p��8v�^vJ�+��a-��ߛ"�F�|;ȇ�ky�j�۾/�!2���v��(��Q-��g��N�+	�:�"���^5������X;n�Ѳ����]96tD�5�I?7w��!Q��]�]vJ;�ZJYg������Ӿ�/��НA^vÞ�����^���4���l/~"�J��M&S�d2ِHķ'�ձXd���3bĈ�����?�I���̟?��;vn�����Cv����L��2@NPq#� Z:�웞�X�v�=]���?L���ϴ�p��a4��F�E�����!)��pn,�?�ًL7[^���{�%ӣ�*o'��a��e">�l�2���
odN��#��uFڵi+:�}SC�a�-���e�N[��k�B۟��\�,@w��	X��g���J@��+�|%b����5�p�o��o�A��w������ٍ�~3�U��Ѹ�7J���!��G09O����6�߄o�/��K��r���_q��ׯ�QH�K�/�w�Y�+!:2�e�D>����o��&��Ua`��?b����+��>c����Eq��$��k�����@�)O"	��S@���Ʊa�m�A]2��@��>{k>}�=��n��*�--���+% ������`��-fK<fF��*�v۶�ܦ=̶з�p�Z����D�@K�ϲ	�\J���&�>�N�Y:��?��Э[W�B~AP�����P�a#��?�֮�kN�����pء�b���1�R|��llè��d�>~V��2l8�1��0>��3,[���v�1G)D�8���m-E2F2������W�,�u{uZ0GT�R�]N�s�B�&��K/E�.]��]/�=��Ɔ:�~;����ttU���w���jWZ* ��;���%��ɴ�J���癶NS.s�G'�g�M"IKZ� Dׁ��L*~w�K	8l�!��,�k_� ��    IDAT�F�^�.��U�� J���@5�~� ��>7�.M�N�#U��	�
���0���_���r���u��˕�qM�ܑT
a v���d2ɿ�&q�\�Q�ry9Ƕ�=���Fk�����u�f�����,8�z��;	�S����ait`�`��t]p\�!�{9S��E��ʲ��:��2�,R���(9F(�(�;?w��U�+�'@WGE7\Qq���<�@��yތ�ߟ�!>��l޸)��"�`Im��P<޶�K�\ŉ`L��%m�w��/b�H��R@�Dab�[����ƚaat&2J�}L*��١�=�{���w��ٴ�y����7aɢh[�
}zwǐ�DF�uQ��������[�@�@�����5!��u��֮ߌ�>���_��;�W������ѫo����o�;n�5�4�S�[2�cx �[n�EҢ���o��oĝ���?�	Oa �G���9��<$cI���C�/�ց�$�H�c�&)��B2`��S��bm�Kk�P�Hm�J�����Y_a�~�����(L\� ����O�н�zK��ֲ�����C�B&�ے�2�u�)v���'u�U�A���h�%����e 	��Y��iz�_�
��� �j���ϕ�H4A�)���u��U����t^k �ؑQ\\�-U���7�~�{� ��c�	��H�¶%�⒕�R[I�B�3�g�8� 1�a����zG-�Vm�����'����}$�d�c����]r1��艦�*+ץ�r�\�;AR��T�)��Ԯ�&�����A��D��L�kdN@���D�p���|�lwZ%�:�*$j�m�R��N�͜nI&�[�� G-� .�|��������Ƒ�A%��El1�r"� �˕��R�T<�r%�������Eq����� F����z����~�T*'X{���;%����\.7�c���Q��K&��d2�R�-�M�|Ts�:�8����,�˔�x"�H��I< _�t�D��$�c�c,Kv��A�S?�<~���Nݺ���իW�s �������Ùro��@�ԣu�憎����8\�5�q#s�t�"ح�ŉ���̎е��th����,[�Q5I@��$V1���Ga��R�����'�k�IY�T�c��W_-jm�HXj�tF�d�+�gk��)���'�k=[�5t>��y{(�<��шx�~l����?��f�\�9����CǏC��Fz��~^
Oa�W�Z��s2�x<�p�(䱍~�Z�x�S̚5���Ք#���d<n,\���q�Lk��� �vE^72�U�,�;�C�Q�JM�O�݅��D<�F���~�"�]n����Sns��%��
���l�D��q'Uo��hX@��>����e�r4x8n���k��M�p�e8���3���Oc��� ����}<b���ɥY��؈��+�*��<q�t��:ʻ���(E���hȧ=�q�~ɤp�
�N!���E,�����F��"��
��%i�i�ܠ�>8+!ɗk�5����DXģ�Ȏ׃��
��(���J&�ך����-�6=K�=*�%9z�v1���<�U��B>�	<0����]x���x������ޓ��.�	/e��z��cY���.h[j�teH���-�z6�1��D��	�Z3�~ȱ�w��5Mϵ�%?��N�c�*&��J}����غ��#��o'S�\�\��S������y<��D�O2�Lzn�;��$bn�+�Hx	��@  �'������<�'kp3�Ǔ����Է,Y�"��?���KR��j�*t�)��g��f+Osf�14�-�����n��UgIG�J�r�����d�� h�������3#��^6U�<�f`�<�� GqN>�d6�x���kIp�ϲ=�|�׎OT�
�/S�
��	�I��6o@'�N��е����d�[Ss��ׇmY>�C:��/��"�;F�s��sf����5+��M`ؐ�8�#ЦM�n^ÄF�i`+2�圥fh�^�X<��+�]��0i҇�p�WH$�ڽ�=g8�`���.܄�>��<�� :�CXʐ������:eh�i�ǥ��������}�DЅ�����'�S�.h�o�'�A��V(�� �t�����{��F%���c}S��܊�Ł|Hԇ���Oa��;h(��p	�/{�)wj���oǴ)Ӱ�j���E���`�L�R�W�GOu�q�ym��w�K���O���2t#��i��;A�e�!�hBz����G��\�|>8�.��j:�b�[����Iڄ.�qW@2t���8!��sd�Ǚ}�zd�(y$���R@sy	�fz�ԛ�p�d�z2��T	����0z�i@��(m_���?���C$����%Bg'E��^�/
O�7����)G�}K��S�)_��f�U�������O;{�����f��m��7��V&��䠴]�A{�;���l�.��V��g|��������/���m[�X�r����E��F��u����y�x�l[���tm�s~��wX{���
�j�뵵e�߲A=�zV��3���e���s�?^fp�Y���:��yL��i��Ш��92t9:L0�w�=��{�gj���;����;X���,R���A��QZ���~:<� ��`��͘:u
�|�El۲o#��1G�GIQڶ�=m��4D4���]��L��m���^��bWMo�9�|:.���F���}���n�ގ�����YI߱tx}fƀ����DiF��SN��Q�$�Y_S��~��_}	�7�r<6n.��Jt۫�����P�g��o�#*�)�ܧ̫���hp��TG��԰��w�������o��8���1n�(��2�Z�j5����\�a:u�� :ǿr&�\w���#�"k�4��כ����0M���;���ed���[�r��1r5��� ���P��S�Tͣ�D���1�n�ȨQJ��#�Bμp{O��ُ(��D�L���p/�H���	b��$���;'�I�~8q�\�5�%7�xH��~Hב﯀����{D(ǖ-[��Ν����v�u��6-�g"t��3vL�S{��Ȑ��⤘��ׁכm�z�.Y w�,-��dO��c��AO� Ւ��X��=�6��C�/,,��G��[G�tF�F��t��7u����腾_z^�c8KK�������,�֚���t����uc��3b#�[b��s�):OE�uN@WOZ7������ݻK���L�ӰsC�ӈht))7�v���d�SX��#�F��ր���mk4x�v���n�b�l�~6��L�˹�M���iX�ǱϾCDx���5-Z��>���m�dhF���}{��CǢ}yk��P�<	�ǲ�өwz$(��)y�q~H�'�1�a��1e��yK�-F0��{�AQq��d��\+ism�9�iͬ�?a�g�I�����۷7r��e6���kP�n�d�{�8���`��O��.I �(/� �tv�ڎ���pĪ׍��Q!�yA۪���[o��/�B�/�Ne�зgoJ����K�x�j�Ş��(K_	l�Y�����,��)Y)���h�1e�8Ud��ֶe��m�y��Q�%��HP~6�\ �7>�|!�d9h�5	��7���/��H�>�X��{�i;x�%�N��y��˛�D�n�˹���Xo� :,������_���|#�g���(�(�{<x��n?��_|��������g��]ڏ�k`2!Q#��hk�̝�) ��g��H�Aff8���5p�6�����vNI�t`x�:ɢ���}z��{Ĉqw��������x~��p��Ӫ�l�c��U��NR���~w'�z�������Ի�Yp��4�V��	�����Z�r�c���ݒ
A�o8i��t2�il|�4y����?]�g�B����1��(��H~��Rnݺu&���+ib>Ԁ�!����{���x��XC�\j�/����G}T�a1"�{c��2�h7�G��lf�-��1:v63��R��FQFӈ���
E�����
c���8ꐱh_Q��<���5�E6<<j�y�v����N<fʝu[���k���|��"Đ�x�}ӅB���eփ�#5����H)\�'bT�Dl�D���RB`	��cG5R�c�Ѹ��	��'(x�^D�Lʙ��WWW#NZ��ֈ1NfF,g4K��-���K4m� �c4�f:�i愔h��}��ß�vy-��̍�q5:��nA��!Is4�f��N&�4�����>���iv�hF��!��"c�1ЇJ�,��1�i��@��Q�0ޘб�&�0)��D�4 ؛l�����Bv��k߱�d���w(b���8�-Y�f~�o��V�ẍ́�nIq�d��)�:q:sL�@�6��v��X��ؽ)-�"e宩k�2��'<���:ojh��'�f�e�"𡢢=ztCYyiMϞ=~�q�=�}�f�D��?�Q�����M�<N��3��L�+���-,��"k5r�z�����S�F`4�&ݭ� 7�MU���-��R'�e7�SB]�
��4�����FP�Y��&U�h����n����:y��P#�z�)i�C��"�L54s��Q6�; >]�L�jģN��	Zn�M��C5�G�QL`���8��1h�6��ضzdL@�WP�	T�TnEJ�����.��&~�/�,E"����^q���"�º����\$M�����_��(��!�yQXX$�ں�Z���8젃q���b��]ĀF�4(����� �s�d����H1J$��9������ �?`��zB�7���Cr��r���Pjz����̖s-:M��:���뚖5��s�����E�V�lƾOk^[�3|:CA�\���,���L���o�����BFG2t8"�8��R���=�|�~v�Ww[�P�cgk!hy�j���q�7s}��̱�� Z �N0�����ض��Z���������֖0]�Ԩ�="5ۣgW�ێ^���x�qg>K6��$�79џ�o��|ǪU��]AO�=i�u�1W#���w����N��B�H�Q�m� ��+ƛ�����桠JĤ��.ˈ��^U�g'Ͱ�l���/�0/��	2r���X!5Zگ����6�u&�2f�A$����~�i��@�� �Ɍp3��D4��wϠ4ψd�쨳���)LBR{�#;�sǐ���N8���ұ�F[�mHR�$a��\�;"xX"��]��)�G��&�3��@ҕ���
�æ>-�����بְ���nւ�(���(�����oà��!d�����CÙg�&큢�6�]>Oޗ�N��d\�br��8�(�*�i��%HpB���8: G��k�Cg�V��i������N�NI�[Ǒ%i+�h�%���W@W[�ǯ��4���ә{>���[���5г��0��̱�='�v���Qq��~����^{��V��$�ӖiD�֮]+����昞z�"Bvh����%v��ЛOsa�����w9�X�;����WWQ�X�GΒ̐�ml���5ힱ�4�w�х-��{v���N8빟�����_z� ��)w��p�l��58@��Q�� �ů�YJ>�ߘ�*,*�K�hl)a�4���H�uTkP%��q��M��L�*�bݏ��ym����^&���K�AB�Km+R�Ν���'ހ_����?.*[&e�JCIn@o��ů7_u@l ՈJ���*�H-R��$�w�.8���Q^ι��'YQ�L��e"t[�tQ;BT�"��t����jK^��>*��B�]�@���8��E$ݞ��Qw��-)�")f���'�b\".�Y�������Й�@<���? �\|:�W(��m�fk�C;�0*W�gX>���̜��ͽT ����QSXHZ�~����m��#���s:�Ӳ~�����l��gT.us�$�3���;A_�����̻�]�t6�+����@�5a3l<6^oN$�w��;�}ih
�5d�e���2��η�?�][-cX��V9i��Tx�[��t�h��i�Į0;eE��܂\t��]���HA�����;�ٻ|�$��w�ڕ��ѫG�~�>�k�����񩬡o��|;�ֲk�٩������i\[��(9=u5`��9�\7t`mј,���A�S�L��u���Q����V���R��ǧ5mnv5��uJԨ
�D��Q�_��X\4���/�}�|���Ȏ�Mc3h�>���e��X��y"P��c�aʔ)�9�̵/of���z�S��4��h��i�$���(9�G�h]��ph;��0�酣�6�sP���� @�`����䴄oI�e+$Iq[�0���P[�B]�U�u�'<hhh4�"(FYB�r :K&rږ�L��K��P�!AKf�3��V-�����#p=G�v�jJ')fL�"��a����t
���1���4X�s�N<��C�r��-�`�q�`�^s.IK�Zİh�'u��:v8H�ǒ��A[:�E=>�I��΀)9�����}儲�`���r����~�D���H�?��gMwl�V8��E�ϛN1k������{ǽ��Ο9s�{���R��~V�=�%�z���3r:Vٶi:��3Xq��<nZ�9��ro��7�3g��p�0�uI݂$|~w���Kwt���O8��?������ӈ�ٶ�����*)�,��;���[��iF�m���e&���K�٬aԈ���<� ��`��6��������+�P�
?�Ȍ�Y��ᣐ7���IԞ�-[6	�w0����{q�_Á&��$	���ږ���n��(xAC�S�;]��N�
I���2���'�Č3�%��R�u���}7��<��L�4������D��6mJ�z�F,Z���_n0�A��ЃF�S�6R&�nӸ�n'�J;����'�2���f/�U��o�a��0vֲG=����r�od+��s��J��Χ�e� 'S�!"i�;t@aq�p(*¡8��7a�}p�ףk�.�F����h]@Xƌ��c�M�K�]�L\n�م[o�3?����B��<c�_�PSWk";������$ӫ�U����n��ʝ��ɠ�����ӥ&[RRP�{��4�����E��HUS�� ����������L:�=E�N��q��Ψ�����T�^=38Β��b�ݩ6�Βvr��n�39��q\��\;��ӑ����v�/,Ý$9��UVV� ���+��8�WJ�ހ̰�a�^^�N�GYyiu��=�?��3��9����߻�������h�_Um���իWwT@W�������^���Z��'C�����z�4��~���8�cЦ�����;z��հI�J^� ���	�k*_C05z4M����<I����R����H�A�С�DI;�w
X$	R�^�a����׫,$���W#�h��8��9��B"�����rz���-9U|�j=��	���#�ŻΝ�b����ߞ��w^C<^��bƎ����}���CC,KG�»7��ɲ0�IrQRR�.:|ر�oO��U�[�m[H��q�QR\"�����F��f���gj� 9�����������z���`+����HŢ2x~��ߡw�^rE�Z�8غ�cH��qe/�/F���9����}��S&�*Xx��(2�3"{�~���1����^f�G����	 X�5���d��|M�+�g��f𘝥�4�[I�l��v�[�a7[KY����۞��$���d�E�������P��%"w�d�
��<~�8Ϻ��|��c�%0u��:6��̼8�)}\�h�}��-ǩA§��#WU�Ml�/K��ߴvP䡳Ͷ�v��+�h��g��םt��/��?�������������/\���U���z��N�����<�a϶�-�&�d��8DJӶ�q��G�<��lS"FM���S�5IN����V'�p��&Ӛ;�a|on8F`܀Z��ջ�@    IDAT�jڎ�Ŷ(������Z}��sL?�:$J�#�� ��7���̙3E+Z�,��N�-���{ss�3�O<69��E$�uG�E}���x��?c��U�y"8���1v�0�����D�Ť�.$�8�٢&�����N
��N�Y���+�h�Z,Z�Fq��ٳ7�=U�����o��}�Dan:'�Y�^5䝻v�mw�
J�r����%+��=V,[/2h0~sӍ�ٽ��ӴS�TZ_���M���5�EL�듵���/�HQ��1d�l�cђ���r��K�1	z��|�O��r��7$8��f��iB�l'N{��;^�o�#�����$��]�C#mc��l[%���U�����#�c^�ӡ�tPw/�e8��ձ�s�㽑��� ��AHy�����&f]�Q�!���:ά��?3�+��i�{j��_e���)6?{�XTmS���Y�?G�����yQQQ&k��}�=z]{�	g��3��C��G��O�,^pbՖM^�fM�w�y'=] ���o~�;��C�֞�;�R�6$������=Y�L�� �Uf��n,56���ꕉ�MEC@c����ֈl@�Z'�M���#y�QgGA
��>�9���ؕ{��S�w�������-��Yӷj�8k�� "5v���7";�bԬ| ���ax�X��)���o���	+�-DYY!F�7�FA��6"�*�C�Ni�bM�/
��M]��" #�ll�n,����&|�ɗ�k�mF44�z�a`Ʉ���O�I���W�i�&s�l��7#Z魷�"�F9O��׬���܅�_~�d�	8�]z	�t�l�p`D�� j�>��<�H��'�2�x���c�K��*˽��2ٺo�&M��.Z��liAE�+*��{?TPv�O@��UehiK)P
�t��i��I�6�l����̼s�93��m���/�$s�yϻ>�g�����a���D/��ejjlṻ��[���{�m��;`��U̳�
�s���3��p�D�C��S���t( �6��\����Θa����q�Y��,E�Ow�����V� ����ˮ?1� >�C��*}�C!�k� 02��+!Cd��&%z~R��*m��PqH1FI�PS5İ+@9r8輸�!Փ'M��嗯��T����Iq�;��i6�}���U��l���c��Y��]$	;�L�ܰp�Q��ΰ�O�2�f͙�ޤ��������(ܲH; � qy/8|H��'��]8pE���L��*c���k����+����v������g91̲�6�"�Zh3+���b���)B�\32e���7�A�'OV���.��í�ӟ��������C̢%�҄q�('5��#����U�U��P��/�G�x�GI���t���^xym�`UT������/�@�gϦ^y�������ѽ�=@����Ɖ��쵎7ٸPe�����]�L�ڽ��{�~���&�Z�s��Wo��F�T����2�c��Fe�����Dc^�<@2�&P�>��jZ�z5���sQ�s�[ƚ��6�/�������\�ۍ�:$ށs�Q��Ρ�Fh��X�T�q��D����]t�X�a0RQ��T�� T��x>m ]'7�{��K�e� �<>������N�s8�z"S@7�����y3:�YP��>i�����ҫ�����N��[ ��n��������)@GA��1���%2��c���
�n�9��	!)��{���cǰ�5�H��JM� aN�f �����8�͈W�x�p���u]B�w�0p�<�h�HT X0`
X��vs;��Ζ��܃�YT��CՎ��� ���Ɛܢ9�%��'>m���
�K���i�˷f�i��G?��>޻��L��Ϣ�O]H�Ǎ�����/��\mjI�>^
�Pޣ<�9BU���;[h�ۛ�@�!�7o>}���f�'���|�s����K�*5��e��FmB���9���K�?����>z���y���g�g<�U@mХn�-8�]�wwO�;n�@ \���!������|���w}�7}�N=����+�ړG���G�T�9��F}���%Ze�"�]^3�ĕ<�t��1i�r�W��K��C6��ψ�
QZ�̤%.��AR]Ƈ̧�$��� ���!E{=J2+Vii�v��1VD6Z������w�,:�ɘ Դ� F��9!���> � ���A�������B9�O�C���=����É�(�����b,w5ۘ�L9a~K��k	�x��g��xgɰ?��F��'��Aa!N����y�t�dpbH��@�+�j9R�BJ_�l���1Ћ��MZ1���v�ya�c��B>vd)���q�վ��7��
��x^�c�8�n��;pƵ����-!QF/.�?3��U��P�a�Vi�⭙\������g��;!�G�q���,�'��/�������-rRF�t�v�K���\�#����ڛ�}��_d'��f*_=lD��墿����r{QÄ0��t�$T��M[�Lͨ�U-��U�AI��,|8���:hi}\�N�Op���#���\���؇{}(�7�r_�������zv�}(z?q���g5�_����ޝIx���3�����-�
�GO�Gl�Q�.���K���6~WM����c~�#R���7F�L��.3-K�T|����2���H��_�gy��zY��#!@�C���f�ē�'e"�x�q���@@G�7ѳl�������Ǔ��Dc�:\���/0�*����6����w�'?�����}H����v�86{��,(���.Փ7��>�T���"�"��8���<���*� Έu2�ތ��
ޙM"��10_a�hh^���$b 0Y
cjԲ (��"?4|�E�(-���85�1����AUZD�>*�v�j'5tn��1�U|�C_��/�N�t$�^yI�p`�χ��2;�����T���]��}Z��!B+.H�����.���{�^Skm-�����1�9�'�i���'�=��j�R�[.[ᇼ��n�;V5{#
��9���_7�*&$Mg�����K���\{��T�|.�'���F'E)�@as�&}�baQ�JYV�SR�W���Vqn�����f����%��XB��"�^o{Y���6��5�����>�̡0!֭l�}������X��o���?VH>�P'��t���>��kQb*>7脻����.?|��uN�m�	z���;t���VEYȊ�,�3yA���p�������/&aՒz �)�	""[�0��ev�o-
��gf�w�G~���ͥ��=,W|�5��_n�q�	�)�	!:��R�xB:
84C�����
	� q�<�m�,���d���BN
�-ڲB� �ײp^o�ڌ(Q�{��0C3�3XG�h����x��۫r�g�'"�c?h���7��N��Ṯ��������|S0�I%���)d�`|���M��l�4J7�̈́<�6��աv'`���9>��|>�D��o|��8�U4bڲ^+�hmw&�K�6�Ӵ�G7<�K�Jȟ���%R�Qu_�a$$56���R���ӛ�\{V�By��w�;��ʬ�B
#Q�k��|�VyҖM�X]���Lsw&@vG�����1���: Gs�$� ���Y�jh,�f\a节M-�c���7d�<�������fN���p;6h �S�>�?��-��te�zw���p/-;���σT�M{X��k�G�D��~s	I#��3�R������#���H�;{ZH��*Y�����#6�I��+Q"m��3Q��>W�S9Ͻ}`�G�[�AL�CS-1��&�Db��-᱗M�cƶhp���3H��p6���ǻ#\M��XxZ`���Ⱦ\}��C�ӱd� ׀˸�qb������5�~.&{�u�G� �*}يbլo�wM���3���:9�u�Hd���Xv"֛}Mv�2Tѩ�3����.n �ﺹ�@��f &��
Ǉ�r6��䊖:Γ*��E�����hA{����k�	��(���e�|�w��(V5X�l�{_�C���%2����[T�/���@u���s�����qŞtܟ�J-;��2��x����è���^�NL��ѵ!y���mC�y/To.�;�e�	Pخ���U����%�߈G�U,��|��NTՃ��nci;��>�[������]U���.����t�Փ�e�Mͱ�#NXE�̴�sVן���.[n]3fl��v�2�����G`��}����X�'#tD��$0��y2�Y����Oo�k~kn�/M:.���iKN	�M���oM���{>�����)0T�+�Şu�Oc����e� ���鼶�>E����5���_���rf{Gٟ惵��5�5���ʮ��*��&�-Ē�8o�߻FoI9x�o:��&�ml�e$�2C$�Zg�1�`i���q>Pg���gD����I���j6f�!�k� ����$��kw�!Z$g�P}Z��$�1�4Z^O��Ƌ��*5��v�3�}�@����k8':�ۓRik)�����U�z�,�M�e�s�}�T7J
�0�}�v��K,�sm���(���;vd+�$��L-���|�މ���k�` �
��Ě.'�c6�\�5?ɶ�~T]�l^{`�Ӭ"��?��tYE�N|�G�hj'裩�L������9��sԤ��<��At���̈́��u��X���h��aC�?;�_�v��L.q�SY�xٰIBRd�!k�����Y����O�-��Q���X�(�S�~�9=k���;�V���V��5*���\+P�u���Wb������$)�'�	�G8'�����I�[�F�0[s	՞i���4^t�:q�A�_�M\V��d���U�GJɻ
����p��q�PRi�d�Uk�k�\/OTT��ZoH�W�qJ(�G���/�	YP\O�)2��h(��Lk:�2
J��%�p���d��(�0j˯����@��ة�� ��O�2Er�P4��ǰ���������e�T�o�k d����������z�Kں��֥>!�y��&���������R���e��8�Y❝����슍�����ۺ�M^�F1k���`;���N���H㾣�A����xJ�ݢ�
�1��2Dp��ӿ�ܙ.C�L�;,��ްcW`x�l��+�f������R�'�*�O~��m���3K����Fv��$�V\�5
/z��z�_��Q����l��������=�\m5���O?�&��w��`� �#R����B0�}j�z�{����;��P��K�y� %�e������;�0ls��j������o�Y}�@�5�zFf��?~ف�;Y�Յ`TE���ҩm��/�Җ�s����%�ɟ��4�K5߾}��9��x~^�ʎ�*3�7$ ���G>(��p1<�]���hf )�K �Yu�A�PJo�R�ЌӨQ�-���ш�Hr6��	���ӥ� h6��S jAͶ�( 8�lYM���Y���]�p�:x7�l1�}�,�2��J9�W�,����Wr����n=؂���K�)0�x�+o�5c���x�����z����mnQ&Ϻ#��Xn��iЍQl� 쐷��x�޳����'?%�Y��+�_2�|U<��kDSq��'{E<��u8��~��m[�?�jA�fC(��H H��%L���8[�A�2���i�E&�u��'t����r������"�cB�օ����[�'��'������O?(;�/iL0�������~����X�/0��jv�����C�]��'/x�GKu�D\`|���_�$���|r�Qm&���=�o�{rI�pKֈ�������2���L>����w��)����p}��N���E�����ՉP��P��%�5c��������_��3��a��P|>Qn/�_πH�j����_��Җ�7�Xp�^�׈J�{�D
�u ۏ���a��5v�ʒ��[���l�q��XBƆ����DUhMe,5����_�s��>M��~�W�$�{w~F��D��J\�D��fV��b��O��r:��*�p�w�|�?��`�?����*��h�Â֯ܗ�6�j�ke������&Q.o_o=�cm/~��F�>��[��o�9��J�A��S�g�Ҥ!���*%Z@������|��s5h	\T��4E�(�'��&��݌�(�a�o�̗!��ۤs+����3>�V$T��$S���qB�����eΥmF�vUE%������%t��+E��r�d��?���>���+)L[A_�8�J�XO'Y�4� ��~�t�φ�]��D�춢�;�"���r�ޫ	0���1zu�t�|�Ǉ0�hM��������"�s���X wJ��?۷�h;|M��nv�����{�dt�j�;��j����
cW���{
�]���kA$�S��v� "��[wA�N�Q�߬���<������+�uN�b����<�X?����&�%�\���	\A2�I�^��dh�$.��
7������M5d0������S
_>�\�h+_OϊO�beKaZ���}R��F�����������ɼ����r}"y�w�ؗ�a49%n����ϵ��"|�!����ջ�'��a��E�^!t��o�u�a����Y���9P�hW����E��I�#\s�H�c��]��c�o� �����B��g��Z�R�B��[��z����##Z�o�W%��|6�_�(���&��N��/~�؅�5�|��[�p��C�S�����i,�˶|��D=9H�
zU��N+S�̠g^U�a������{��d�������H��;�R��ҵu	�f�3Q�o�N��܌G}���G�;�W&�l<gE] ĥ�IH�Η���*i,�3�Qz:�t�8OoP���j���f�0�`3]�Y*��~�A�k�ci�IL$j�WN$�����v��{7�i�s��'�� 6���^�_��'�������������o;������p�ے.֥>�� い��h�\��.�s�҆��[w���3���>~;�<������QU��($��'U���2	�=N����=��׏)������[5��L�L .�L}�366]�k��o�(0���r��Z0@�"�&�]0k���L�`�^��ue�̛���E0q��9J}B�OѸ�����-Bf�B��=!������3\G�(���qQ����[QX��-9�%y�Ϸr�;�\�qRK ��D�����yRl��M�Z֏� �.>���?9����'���ݱ��c������M�O��q]o)&�S�)���Mfy.ٲ�6
�^�1�_¤:
�(榛��d�3�C0Pq�:bN?H���mMXZя.n!j5�
��Q\�o`#����N��J��/���~?;"gsH�)x�Z�������a	��gW���&%�x��D�P�~�6���eᇋ�g�_�"��xNi��cgbާL���4j������c\db��Q�pΏ^����D�Z�
��C%������a�W����>���s�^�𰔚��-=I�f��UD�8�A�Ht��P�mJ��L�˃�jd��|87�A�[^�|D��fhR((�>��j3OɡY�3 �b�ܟ�:{}_�����!Hda�o��ɖ6(PBG[w
��5�����hyM�3���A�ň��yD1$_Gj��5��=�#(Z��������_a�$(�GZD�7���Z�Cs�k?����H
��12�&�eZ$��b��Iۮve�Ꮨ��_��� �ϝ��Ï�˒K�8��]�?G���I)�ח
2^`^3����C���VV�I�g�	}$��x��'���
^[��u����P�ܐA�ű~>�n$kw�0GU ����n�zIao��grI��)���K�(k�MM��#}�d +��i�I��&C��I�=�B�d��䒣0)�l����Vo�p�&�Ƴ�:!�E=LԵ����7�@�Ӯ`�?y]l<X|p:�R`Q�@8�ש������3�X���� ��6Ltյr��e{���Q ��ZH�;�j�����%�v��e�����*
�x��]�U��sr<�R"�q�����b|_T�����4^9�|K]l"�R�;�:�I�ӓ�O�=P�^�l!�������D�b�5�+]q�غ.Je��Q�W�?e	V�ɍ��$K�9��&�O�;�&��s�~��Y��hi-<��=�����J�m���1�6��^���yr,�u���)?��{����Ұ㌪����&΂�t0!F�?���*��Բ 	��r��O.y��:=Ud�-lbWxVM�����gZ�����]�z`�Aj$���I������O.�����^�*���N��7)9y"t���f=F�"�Q)2ypMV���߻���;<J'�w*	�e�]C�����-������K��޹>*�����=W���^�BKEhr7�G�<�"n�nn����LE6��m�����*(�IG2_���:��}O�~�U3�\&Hz��G�8O�X�1�Xw?��r��7Ԥ�]�%����Pv	z�y␨�]t���>�F�\�A���KT�.|#�7rnI:����Ff�ٹ��^Wa|��r�Y��>ē�*nc����c�k���F�����H�KC�	{y�)�t����
����&#w��%#�ڔx]c��l��~�����wG�GFq���$�׻�.b��4C֐���0��6x@h6��z�,��
�3窥Ul���mz'�'��:<�?��o	�)}��F���<���@䢌�q�Ӵ��>:�����GK.s �+��JK�9����Y��B�^��²R ��K����!�2,AA7���V����C���~a�U\�A�ZW4�>M`R�2�&A�Ư����x�~���K�y�	�Of�>�X-��5�f�������A�X�Gr��c@.к��0OlS�Ħ����-���St1}y����w����J����Wvipڸua�q�r\��
|	�)�\���������V�m�~eO��3׶��K�z$�5S��$]�r��}��V��!~���o{w�ա�U8񥘆uffP���iOO۳*� _.�8�A_����a�P�K�J���Q��)�P��tˮ�-���f0�l��2�s�h���Z��,Jh+�AD���.�:G=Z�h���z���c���N!h�y��4����h
L��P��jSc˶A)��,[k�c.S;��O�B'�'�L�(T:������H �}��H7���%�'�鉋�=6����k��d����d�����N�K.�9$����[��7Y�Pϰ ���4�jpHr�Y?�e��S�V�xZo�='���<�.��|ۻ%{��K��ّ�����~u��/�(.�K����W��l�������wλ��b�noU�`��k�����$�����L0��v�G�4���0��G�!s@�����c��;2^Hb�t�r�P"��9��JjY�h�F��a��6�L�NH�''R�̊3��-b��7pN5�V=�.H_����X�G<��L������>���0�7V��.(���w���+��#P�5����XP	�~�pBL��g��Tk�����)��Ӂ�{��%%��<j���i�C89TP�ͼO�c4N\
�Z���R�L��Xe�u��$F�bp��33�Ტcl8D��H���S�k��[{��=�����	�����7�8�'м�
:,�|D�w��S$�P��MQ|5����-��|��؂iv�Տg�s7�C�(o���+].|�q��Z���qA��)������ʍyL��!Dzv�D�f\p{f�\�'��o�N��N�J��h�9S_�*���G��Ɉ��k���f��ˠ��p�V��SHp����dbX1<��=\�N����M����7��y"���ԑ�|~�N�q�x�L<�1QE����ȏ�׿�j:�j��:(�ݞ{1S�$�MB�
���cS�}f4�N���Wؤa_��2�s�+I,��u �)�H� \����i�j��]Z���jhT�3��_Z���",�����<c�5�@�?e�b����h���ň�|�M4U��֨�t�S?�ɰ9�+;����?
�C#綤�B�����S���2�Г�tM��*C����3"�]מv��}����0�gT�>`����*�M���.	�҅b���]Ӕ����v�Iğ.��/m7�c��0�Mkɮ�nhО!��}�X)<N�:�A�q��Y.�7[E�7&bb^�ɕ����dp�g��)Q�׷�MC#��O���{<e&-���NDV���s����I�\�vlp��V�|Nuk����)j]	���L����6�L�Pfϐ�A	��"�leEG��L��I���f�Q��+��[�)���)��en�+h��ȱ��+���D����T�Y>�!`޾-!���.�%�Y����arV�(�9��hQ���rH������vL�BJ�u���l\_ǒG�YH�{W�~[��Q���h��z�r)��O�vDp5!�/
N8 �s�V��<?񜾶~N=/&-f�ߎv��б��z�ٳ�7|���E)�kKjk��#��`=A��|���Y[Y)�{|��
�s�&[�������7��ͬ�	(6@u���{�(H�p�,����j|�p_�P#۴�q��w���N�����YD6�"�Oa��c��E5��V[i���E�,���7�*�Ey��,Xn�������U���<���{ ��G%B�eb�1`D�{�?���.6��&�M�\lGY]��&5��r�����:n���2�۟��L�~3�k��2w�����Ydd���w�֗4+�Q�R)�ʞ#��tW-�j�
�E��G�lc2Km��ˁ�3?]d��{Y �ӽ����G�n���j��>���=ۘE�rM%�O��w"��B8�!12:Hɕ�FO�kVWl3ACQa_!nm�D�(C����#���]�,e|�y8�]���S8�b��R7G<�L^LHҠ\�gk�����D~�&��kC�$h���s�	��b�6Յ�|�v?q�K���Q�,T#���C\����M �����r��`��xFaA���G����>Y&��q��4�r�EC�"�l�h�����PM� �i�c �ռ��J�'��#�[���b��mv���J���`� �}+l��&n����~�0'�&!�#�3����>���s�*;�L���ca�ų�:�.�P���\�p�)�E�3�(��leB�ڣ<��\�nI6:����;N��@V�m�z�8*8�G*#R�5#��N�b���>�`�l˯��i��f�7!v�Z�	)��2��~�T���7wxI��Bn�����2����/�e�`D�(:�α������@1"���e|�:�����M|3B���<)s���6c��v���͵	�y�$!EM�G�ҞTs\�cy�y�Z�q�5q���t���)~v������ɩN�;W������[2��f�b�[ �7�:$�V�n��K�֑��� 7?"��h�}eۯ��t���g�[����2��Mq����Y!C
O�ju�
L�\K^6�S��o�!j%��w���j�����F!�ï����o�RQ�S� �G�j:�P��u�?���C�9I���~�2l����β��c�ᒂ���	0C�)u?�$OE�/�'�rp%���6��ޏ����D�O�=b)�(T���#�{s�27�p��(L�"���T��;r��x=pL?D��B�,����t#	x	�R$Q�������n9�JC	+�-�"�?B��K�;��"�����(R���4��k02�>������j���=�"�۽���Ab�8X��5���'�Rc'.2������Kd0�ofj]������TS�8T�#-�%�p��Vٗ���^�=*��c�	�}�?N
%�l��+�M�OH��<ӻ�=�ܜ{��+)W�z�LT�k���s��R7��͂? ���g?���m|Ay�E)�>���Y<N3LK�8����#1�5{>7�'��䝩CJ{�$v��4D�|�a���� [���?4�7�I�K�m�,���V�r�	���M ��T���3���=�A���-j��Wti�-��ݍ5@b�"{½w�M�eՔ��1ge�ׯ5��R�^"2J�0�����$W���{!=����1n��S�������=�<���w�Ej]�u��&�F%�e��� R�4i���ɦ�j�rK�wB`L�k�xI�^����ZL�����z
yE�ϊ����!��&R;T����$D?��9~A�c�� ���G�����su95�|�k����Θ����P3�$l�+�:�&�G�e�z���{�)}5�jO_(�Y�)!�f>6>�Y�9�y:�P��8|����Y���,m=є}kz�
	�P_����J�-p�,R��L�IOsm?t���7��{g$����2J���<h��l�h��8���Y��ӑ�d�g9��=�-���z�x�@�o�lP�P�������|!$՜n��§HH�D�!����-��{F���˰'	0�	c+1�,7��q���rs�B�;�"��������=�s$z��n����^�I�T�oZZZkRR�Zh(j����K�\��(�(���CO����g�� z�ḧ�I���L�+5o���}԰�L�7&X0�$"b″�����	�L����;sc�1gVV��P$0�S�[04ܭ��w�=\���;�ȕ/�w�{"�>'��kn��ȳUa��PPG��pL1��B�t3�+d���-�ڰ��3$:Gŕ��Af��].b��je���̀<6���c��d�5���u9d�cC֡�A�*�+^\H���5S�Ųo�~5��;Z/���>s�i��}W]��e��O=,K�b�����$�҄(ؚNF@O����,�n�[ W?f~�n�,p��y��lr��px�\�r��a���HF����4^�3.�p��ٮ w��Ƒn�}b&�����l��[��J��1��Դ�n�+������&fM�*���|G`m��竃٬(
�k����Lt5�{e6.((��4:�����������G��K�)a��P#)E�c_�RIQ���V��&7�pa<`��\�IK��|"l]��eO�+�=�m���X˖RNV-2�=6�<�cnX��j p)�]D����3Y>C��$�^�ԇ��*���T�����,�����"��}�J�筛>J�dR��W�QY�� q�m�y��|#q��\J�zEWV��9�aM�����ʞ�8
f�B�I:��?r:�v����C�nF��O�X3l5�����ŗm�e�����8y����ǋ�Rs�u���0�\�}:v�PߊC�@���K�e�s���b�#|�i]3���C���,]&�N�.O:��"'h^���:4+  ���nJ�I<�߾������'#3�x��8o��h����ǈm�X���8��~U�=�������Xf*����5�Kvn����/##3o�8��q���v�?��g��
^�gV��m^����8�C�{BG�P[z����ޚ��\;YÂQu�3�s����� �{\����L�L�����+�kt��4?g�\��|sU�O$¥�+�SO�M���ڙ ��m������ܨ����)����v�%ڈ���H��I������z���L�D��c}�ޮ��H�K�� ����q�t��(���7(؅=�x�>Z��͛w���a�^�~�YO{EyyoWБ��q���)�u��& P2���jA�a��O�s�L�5��l[��C���|��}��H���M�Q6wl�|#�$�KR����o�����~�qi��pi��$6�h������҈@�KQU[[��O<K?��0��Q�I�
��I���\Cc��u`]�SQ�M�S���������a����M�@O�'��:OR:����!d8"�2��>�Hh��ہ<m�*_f������~�7�	8  f!4Һ��/��������.��vp@X4�
寊n]�Zϔ�.c��y�E���,db)l�іm_�X��u�B(O ������Q4�D�����\^�����y�2Z����g\��.K�$���������HaK7H�"��݈T�tD���$��ʗ�Zk�R@ẇV�)U�k ���N)C�Ut_�HX���N~��{`�L�J�A/K�?�����u=<�2R�Zs��pҢTM�:�C>g}$j�e�����+�*7�n洌�;W�(>�����A��⢢7���4�fwlFLTx84�ʀO���۷��'�,�P�N��L�3fV��}��~�=��\�����Ov!��`ԜX9\d*VN��U{����SoCכ��Fbsqd84��tI���k�t��\&Z=�_�jm�a��q�yy�.v�$f&S����xY�I������'���~��l)��u�0�Նn��`�r�EWS�G��v��D
n�O&��&�$q1O0!e���:W����߼�<�]a��ʥ��#��/��"J��w����3esK䆵8}���څ4�/ �u�/����;�r7m�:��\T�S�;�fm��kY��^�ܤG\�<G5ν�7��j�&a����K:���~��3N�ux�V�
����?bA>'�բ��Uc,ԅ`"?!]^
��Lᦦ�2^+��Ih)�~"}Zsȭ�s9������wu�xچ5ē�;:�u��
�?��ɘ�e��s��~�7a#j�?��`�����0-����u��U10X\!xj�j��~��u��V"4j�O蛝`����kd��}������z[DL+�}Qdx����$��?���[���g���[����ݰ������\�^o��X�"���v�����!���� ���s^h{'��\z����6����/�N[/Ɨ���}���+R��NW�Ǳ��c�a����TQ�WtdP���n�� cm�ۦ�ɚjw٩iE ���\>?;���t����<���#���`_��/��ٰ!�ր�4�o�.����	���m�.����SQ��2阴sC�g$��f|X�|�Vn͟f3�/��96�
�B���-�������ğ���ۍ6�e����K��Y�ư՛�:��#�{*&��Wm9&5���y�Ӄ�e�7��&%��t���2YYT:���m=�!?�5t!��u����Qv�
��v�X����;r���Y	�=^�����ɛ���W�1�򷊞����O{�Vs�A�V$���Z�TʕiN�o�M?�陝\ԩ�܍�����b�:��e�h�:Q�9\�c���e�W��Ɩ� �!�Iy�$����֥��i^���� �N.�0�a�GV�n�F�B$��E;�n����Ru�⎩�q]H9m o8/����e���I����"�!�8��PB�G�*dH�tcŻnE�[�1MV�hU\��e:LX9l�1���7�s��3L� kCH����Z��:"�� ~ߑ�߹e�˜����ݞ{���}�����e'��P���Il$��#��}���-��b���ɡ1��L� �˯~L*��g}zm�*=/i`L����v�:�Ʀ�G���v8�1c��
HU��8�
Ӷ�{�,=�s�̏|}-��(u�c	����O��q������!ŷ-��1KE�/�A��@�4��r�����MO���<A��G�^@L_mL�+�H�w��{bK��lIP���}� 勃2�'+�)}�(�O=���U��Y�[bK5�~�%3�=u#�P~��4"^������%��_��q��rѓ��A͟%�o*Mۀ��j>��C���(�>��(D�׳>�D����bcX������lBt�����Q��� �c4+���V��/�_��'�s0�r&����Q�]H�H�����	���}�l+ V�������O�ۑx<�L�]�Kʈp�lT8��������i/l|P���!����~Oj�@�Q���̤dm�NF�`2g+�Ԯ�24�[��#�=����!U��������y�w�����2�=¤p��6c�O�豳1���S�n���� T�|�Gb.7�ᄕ���y-$�'��}q���,�s\������E�b�n�*�S��vM��-Ӏ8��-����}�F��:N��.���,���5Ș�ϜJ�rNo�=/��K�9��l�E� '		���M�C�+�Y�Sj�7A�d5iN�͌7�9��r�0o����wh��{�x	�}�]��L� �Rv/f��xQ���h%X�c�XK�[�W������F�w4�����_�N)0��sͯg-�u����tA�����;���d�k�n�T�؂`Ɯ�ܮ�#vN��Q�:�'�k��}�������ia�T�Z�+X��"G>Fjf�r�C��8s��5g���9Ȥe ��J��+u0���6&���X���#xE�G'�2�/.�Q�K�a[�iZ*x/�.'}���1#��kf�#a��S�}mA�f�gI2��F����D��Z��Ŵ)>�T���%iC���L�li F�Y���2o@��K�\��Q8�j��>��"!"j��=r��M�-hoP;�y��ǵ ��ŵ9	��}�X���%ѥ��+Yi�SG�_�bV6��.���}Z��~%]��#2=#�;�>M �u�*�cħ�a��kUd0S��O��zS�����D�?�",d�C�N��_�ݺ�wm��3e�-;jo����l���}��d��57�&�0�����o�=����{���>�d0W.@&_[*H{�oW���|<�^�}�"lK�N:V.%nI`X;߀�6�Byt�>��"�i��(���d{�q��վ��:k:�gU�H2�n�%�=6W�V[�����Z�w�y��$ze�x$�'��N_s+~P��).���>q��?����6P����
��()+k�'�@p�BR�0�A�o���?�������ӓ�D��[�=�@���7��G������J���cqγ�9�"��u�H���*ñ%}�J����n��n.�n@V����Qh�T�e��p�v5"Xf�՚�y`-n��u��!V��~��d)�)�T�?R6ɯ��B���s~�'�
75q�&GT��C��f�X=E�[������A/�ȱ~��[���)B*�Fa:��):��h$��4���$��u�wʧ���!Ӡ����:����)����J^�W�2m������O��/��/��Ȭ�aq����u���^n�b0G�Fhʊ�w�O�y��?~��^U|J��T�k�68�dy�рTH�x�۾�&ې=�s>I�\f�L]O:�Ly���C�V�ej��KZT!�w�:tB�y���}bݝ�:4�:i��g/T"xH�	�ȗx;����"�U�W<�L,���f,E-�`3�NG�-W����	ID�q���z��l7�Z|������}�Ŀw~�tt�&P)�af���)��`���A��+�S�d���F�7Z�5ά���ɶ
���Ud������� �iLh=	,R;@��w ��Ǆ	|�G}�B�[qs#���f!58���q��ż����wN�y]��B!| ���U_}�^9�w)k���wڝ=b���:�̇/�B�>�᢯*���ğ��j$����Nm$U���$Ζ���EB�X���E��-�o�^Xc�e!x��mU=0����=���P9������A�g� ���Ƀ�JYiY@QE�	;��
�O;��¨�9��*��������H@Бۣ%���{�GGN>*���ZhΕ�5�Ͽ(Nq�e��TB����7.��X��}�t�J�
LHu��R��c�O�{��=J�y]�̇W\��zΫ�k\i��a��}8���!�IIE�P���z����O�K�J��=ܜr����y �g�P���8N��!�
ݩ��&��(��}���7%���V��i1�r �j��Q?פ����r����0���F&��ݑ��/XX��N_���@�*`�u+�hy �LK����%h{`֒���#��r��>_�~뭥5�7�i)���̆���;�+T�T��u�0ۯ��p�h�1ϫ�R��kyu!�*kMG���+�+% �B�)r.�*����ht�����`��'�C���Pe��\����_�miv��o*E��~�ѽݽ1B�mv��Oj�.չ�-7z/�OR�	<�HթIMni5_Ҩ�OgL��}�L��G�3�D�D1�&k��h�o�g�4~۩�B5���ʵ?�����~j���������B��{q/^(/�P �H��Rܓ�E��k��E���|y�g��ϝ��5����^�=W*�u5$̀>(,�˳�,����y�<9l�����B��T3Ŏ��c&����?낞�t�S8��W�}��IZD����%p��aL���d��!�s��vXp�/�Q�L]�� e�u �Ia��&��=O�;�rm���%j.T1��|�H=��kV�^�{�Z~<�ij��3���4�^����9����ۖ �Zݗ�J���w'Q9\
}(��I_TQ*��]Q�~t$��̳�]-���w|��s�U�m|�.�y>D�v�*�ǸY��u<(c,�@�9�[G��>�m��B�L�/*nR�c���~�Қ��<�[�B��L�ebM�oeV��I1v2�}K]�VѨ��!
�$>U[[Ud��P{�-�x�����btK�S٫�Fd폢e�2���N
��ZHG��{�z"�.%D�bv@�0����ޑ�쾩�Υ�`N��r�3 � ��\(h[j�̨ӂ=����1S�!k�)�Ab����ކz??� �XA_�]0	�F��ї�m�`���(��I�����́j����'�r5� �f5S{.<CZRSI�cPP_J�e�ʫ!� +�-M�r!����]�h��{�8k1���:Ff�5�9�j� ��F]�0i]�_�̪j��js�ϥgn�D��a���Dv�?c*3�-�hlA�ů�G*�I�C �D�I:"��J���'���H����uKL�7�0�l"?�3����G6i�Df��e��g���~�D�>��"8������0��`�Ou�s�ӹ�z��7�~�D�AJ7n�CD��7�D?w�8z#����u"�&�'���`�TJ��r�UV�����^Io�ޕY�ycuH|��п���)�D.>B�9�D9�ޑ��<��7
9@��tZw)�5ឧ����������p���3Y�\R4m���m��cN��<�ݻ.�p
�%�A�^�u�'MO,3I"����&����E+=1M?i�h�Wag�
�NIc�ٯ��fAx�/�1�Н�Z���5��`cg�6��5%[���š)����T�$���U���fK��J�][����픦@CO
t5�ފz-���f_U�jI6H���T�0&`A��4l��5����	
D�X���ݚ?��d���}�IG��5� ��"�8E���X[�Mcls=�PH�����pE�$��e��5{^̈�w^�i��0��Ҫ'�zQ�4c���z�U_�[�-8� x!˧@�&���5�=�����Ǐ�.�Ȟ�����Wm���`�����X�k�^��+y:�#�4Ψ�1og��~�� ������Qgv�oJݎ6�Ғ�k�>F��,�^���I�o���D�8�8�ߦ,t<�f3|FS��X�D��M�xʈxӾ}��}�]X/��=K�ZdCHwSA���('�Qi�G�Sk$b�� ��·��T�?�|�>�ov�%z�"*��v$��er7l�ׅ�vŗ��Z���S��;p�{H���u���q�r���$�V��7�ْ�qc�qy��l-h�u!���Ǜkl<5���`s�I�CF2rh!;=g�T��^����Q-l��d*�bߗ���Rp�B_�x�������G�2�Q���$((�v�|R��62^�����͝���N�[�˕7{����W|�M���-�JD�
�>s��I�&�{/x\9�1���C���m/�QȈPFMa.�Z�x�1~��M�,��W��]H�nmm=vVߝ�<yX:;\	��� bq\BKY�����s:�G��p�ܻ�P����њD[q�������yCzG��V��eU����d�F�'����<S��K���N:]q���Rb�P-(;�`�O���a qr_�ɐ�:LDA<ɪ�!���(�|��.���a����O����Q����Z۽������b�E���bB-�GL�HK�;\�N���Vp��[�%f5���&��Hn{�A�'C��N��ҫ�����BK�1 �>K�Cgr�Zr��C6[s	�A��a���5�n&�]	?�)>�tL�}��11�W8ݤw��)Q?��`KxK�����TZ��HVy5���ˬ��JK������l��6cPWg~��Kl<�����g_t�wZi���0��ec;��.�����&���ֽ��]�>"��	R7��^.s����gc��B��+亹?ՏPo�C����Z��G�t��gi�1���Ʊ��9Uv����l̵*�:D?��n�a���P9����)���|h���4m�b��I��������&��p;�[ʔ�ߪM��j����p@nя��jC���%W,�O}�����*k
��F�e���=��˜Ɏ ��Y�.��9�_���p\���?�������U��ߘz�5�=vlL��E�̖?z����fΟi�ogP��꒺���"n$��{R��g�GtFq�x���1�1�ă�\7����Qw.���0ZygjQ�����w7S��J��3�PwG�d}���(���Q⟗Ǧ@]s�L��4ߣ�.Y^6�@�+���Sƈ}����}��}�w�����I&�4_Q��C�C��z�#��s�����7j<���ڄ�����t��MҿX�BY���ƆI�pTķw�|�\�ƺT�FP�o�����EL͖�>rP�����T���UvF$WHC�P'�JC �S��755�>)��L�c��ħAu����x{��ݵG��$��t���-��v�1�4�u��0N���jޚ5`V����&�r����[sc���(O�:��^�G��,����s�' =�5s�WU�w�X�����\��b�]X\�m-3�2A��ǘ��*�\�����yތ����x��X�\\�TT��קP@���J��#(�n2/���Օ�G�|���Z�ƏRY9;�U��.�i8�h�A��C�m�2t�N���n`�ۇ������w
Ą()I�f�'�/�h&���|�~�ռ�\*���V�_�n��ʿ_0W�˖���^�c؈�4L)�\��{ig[T�"��X��ܖ/=s��̫�W
	1
��A�ZɬZ��	iͫUm��'ǭ1�7��	Ѝ'���x\�����c��#��|�&�<����0]}��vz�AL{3&�˪�y4�nz�������y,�G��p4ۮg	9QOfgg�R����W�'�D�P�D��i>|�f5�^g�=4�V��D����m�����A�1-�L��|YǦ�	2�/�[���F�ɜ�����O2��\m3���1k��Փ�jh��0J\:��́&@3�n��a�����RRF���+�x�z[��e*1[vm(��S8�9ۤh����e	�_J$�h����--Y�xh���R����`�YZ�T�ǞԽ#H�O�����s��dl_�UB�xliV�: �Tv'�r�J,o�mX	A��W����h���Ӓ]{�rr(�X�8�t�7��[q�a�fEqq1]ԭ�`��۬��X`±��ȼ�T�~����;�����/�~��{��n������T�^H�W���#Dv��0��i�5�ෙOO�2�wQ'3僱֎?j��]�1�1�Q�pA���c7����1���R�L,�h*G}�0���ܧoӄ?F�֚=���0�����<��ii]�@v���K��Y֞�7C�Dى�\j�!4�J8n@��\K��(Fˬ�>��\��u��Vg�f$��l)�%��3�M�:՗W�Z�����ΝI�.�/��Q�6���<<v74�]�1�3��������{-N�u�{c���T��w�K���9��7kg����S�4�|P=tpp0��?k`��� ���;Z#��̙�H�!y��6C���B�sc��1�OO��|,�B��M�����{`�`�C������(u'2f�HKa�vz�户S9t��\W���/���[;� ���A����		P�G�"/Ҏ�[�.1�q�"(����ڀ�H�M��;��X��d��!�w詯��D���#Un#�������-A<��F�#��pp�j�=Y�)P���V��7a�_=��R����֗���<�+Ys6�L�*+��ʐ���,��_$p�����.<��O����5�I�&��KϙL�GW�)�~r���}zq���̢�7��Q\j��|��f�@#y�F�D��)t}�ܕ4nrG��,A��!.9��t�����͌�"�Oz��s:�[/�Q�䗋},��b��Z�.�@O��R!s!��ƳM�A��������t��4	,"$p�lژP��ST��7G�涯vk���!����]漒�S`��i �� Ĝ_[�S���20�� @��P�]6c���I��Q1��T�[������m�8�k��76V�P4��#~y��[�hw>��ʩ@>�(R��@dm��9#�3f�ᲊ��G~���7B����sd.�W�O��S��4,8�b�� ��:X�f�m����P��KX!8f�x����hW����L2x��%������&����_x�+Fe�0�w@	x��U]���}g�r1M�J��~���*����=���Q��̠l��V��,�" �:���qC9khE�5�G�/�M���r��+�h�(t,/���^�ٌ�,0H�|�0�X/�g�5X�=�J{ԗ��<��p�s]��{:�SZQ��Ux's���0�[g�H�)����;�e��_���^�#b��V��PU��g��t��rT2"�&�7܏��,l�î#ʙ���>c�'	��#b�f#�%�r������&[���$��P�?��'�����T��f-?rNu������X��h����J�C9���T��A-�7u�]�+�:]G�B�Ɲp�.�u�.�&�tf���I�%11�ͧZؿ�1��4��ǋ0���k�k�?�_Fn1s,`�g�5$�^f��h��Lk,�݂����]����K"�Շ�Gm~��t����H^��ƺ��R�+��m" A��M���ˋt��t�J�{�u%���z��=���si��Kzf1�������g.�XW5�T`~�NIm�X�s��L�[�Iż���s�X��<d���{�\�ŨmS��Ύm�h���|D<7X�I�ĿǍgm����8�������90|t��}�2I-(,T&s�]5��+�����T�s��y��Fd0��"0@���Y��P��xY!��0m�^��>�|��r��@���~�Z�t��5�Y�}r�7��N�����,U0�M��$ӟß�%�O�Lۦ�&�ϭ�,���#g�J�	N�U�ZG���V�ha�^Y9&����^$/F��-L@��j����-=m�nÙIV�(�7y��C��co���و �1������]��q<����㡩��pKq��*�r���(�o�b��N�,(h��"�QN`�e��Ѹ��r���<����h+6���|�II�5�D�Ӳs�֔@�[���[]q?�'W�-s��6������hkkk���\��|����
f�����ɜ��U��w����*80$?E�fw�ˉo�w����b#c1M�Yf�T�>j�U�����2��}I~���_���{^
%����\-��o�HR/pmj�a�mHa�ӋV?�=���|��eJ���l9����3"\��������|�OHi)[y��WMdb�wb/�bA�qgW���2�Գ����>��/�c..E�����4z�}���5�;2��0���~-����rr���^*h/=�ji&�ȹ�#q,f:/0�Ġ�󹿆��̀_tu!��
��l�D�I�A��
y�OC}i�1��u-�Ӯ�뷁2	���$�I�9�?�(�x4u�X~�%?�� �ڈ��"�ă����#\����СﭢX�5n�=:t�ʤ��ZwQ>����[bY�����I7-�>v�w��O��/�j���Mn_�ǅ1E�'~�[�-#���2G��F*�A�~��������/y4uc~}����Ȝ���Y���3���m9ƛs�� ������S�O�(?-̾��O������,����T~j��'��5,��3ib_>�����[�)!��l �-��U!���n?�D�ch�������E��es�MV�;GQ����ee����C���
X���4KW)$�tS�!�MA"ؠ�o����T
<y�
/p#,�-��jS��wX/���tmJ�ᣤ?σ�?�A�fK�1m�my%�8�?����l�������|��;$��ۗF����]�dL��롆�W��,�"\D�
9�q2��.ddT����L{]�7y�������^���بY�D��gZ���V���q�kyܙ0|
��H���O9Cj�Մ�����2ҵ�z���>'R��R%woY�pjZA^*��ɸ�=}߰U��;���N�󸙡!}C����:�Û"#���,�k��?�����2t]=�_��U�$yI���]h�X�ł)�4�^Gb�ˤ�����H����&�`�V���b��ww�����$Jo�?��44���&���{@���:�[V�I�hU׏�f�s=�gO�R$��E����	�d\�c�V��{>��MY�Rq��*s�	�9���R���إo)e*7.ß��m�	'k]�u��d�W�JfM��F	�t����\k%����¹�SQ����@���&7���X1]�0���i}"���Feb�\�_�c���u���t¼�DC^igq���OB�x�e���d8�A;�	Tc:¶2��]_�L�2(ŉW�O�>��M%S�t<���`�*�wWRxF�'w��ܕ����:������ӊ7��q�]��k�������>�NJ�i+l�Yf|	���dv���;P���:���ۃ�X�IL�������ʺ5�[|�M�+�ofaD�d"��a��6ȋ���s1��.�D~�o�w �*4��)���8��[�������^j<>�%$��mhLo�+_����?G��(��bꮓ�~Uh+�� �&%9Wci)P��X��+���cjLh��F���/�0����=X��u���%1��,�b]B�����"��gwM��耯,9�Z�=�>pY���~D]����E���[�y-\<���nA�)K���N�H�XW�榬��`�����9�
~t2
z )?����W�ܽ�֠�5�Y�t�w���o�;�"5p�Wsw�m��ߑ�R�i2(m3���G����ʧ��gS�l�3_U�$�T���(}�6�0@@q �l�B�q)�"	O�_� kDվ3S�z:�DVN͖�O�0���lz1�B�\��^����<V�٣n73#����ji��s��($�}>��}������^ֿp��Of���/$�f*sQ���ɺ�Hvjy�:�%�c'����9u����]_�	Y��V(|5�A���=8Tϝ��苎-�����vN�������N`.<�46ƒ�Z;g7���\$|>�p�*��H���B�`��>��+`��]8��"I���h�7)2#-;í��P�+ټz�� 'GΛ������2���Ȕ:��y�(�3��E�������hb�R���c^c#F�?nHz�6MD&ACS�4alJ�zx]�E�V��L�W��AD�7�IZ�(�*���KI%���~C�X�{�V�4^�x,���υ�.�/D�%8^��\����b-b�'������e�w���=�����p	����:��2����P_�I?\w:-Tݵ� Z��ĝ}oP?�Y
v��y7B��=�|V7�b�|�yp]m��p�;pk���֕Ѳ�ԝ�-�H�,[�	 �vVz��ޟH�c��]{%MA}����rKt}��L�9�Qr�W�i�>�fs0L1ξ�|N�V����
G[�m<9�˪�aE��tm�'��x�����D<�,�@&�^���� �Y�ĈH3$ۈQz�g��Kwㆽ�VcD�_EE&��i������[�G.�=_����OK��׽@	8�]l�Ң��Cx�ֿ��������/�4'm��|��*P�{O�6��7��aj�>�hi��x1�A���ły�k�o����5��\�N2�m2�Ǭ�L�iI|�i���ԜN������$?�H�)Ȟ�W���;Wك��L��k<u0���	�կ;��?�
sƁc<_�ɛ�o���u:�8�X��_�٥{0�5[_��߯���]�Q�ڋ�R���|�`SA����*?��N6]6
��H�NO+ȇ�q7���y�;�����ߍ�ѧ�;�yez�p��	o2U�F����8��{+� �����P��A�Y>��%��1��؛�?�X�v�1��0wL}T?_c�a��U���P����]� k��Ќ��{Λ����� 2�iX���-�~x�
P��
Ќw��O�1��f�a��l3�-Y\Mv>��o�'����+�ʓ����Z����V�_�|R���/=����}5�x[j�p<�y^*���"�3�K��8����繹��>cZB�n��ȧ[�9H.C�9����;�ض��(������7@B	�bY<��q����p��J#Y�_�s	�9)�CL��jѭ���,X��{X�X��T]�p��C���gO���jȋ��W?�RU+�am{�FH=���:���f@�����f��o��>�l���srrRsu=��&|q{�Z7q7Mɡw7���`�?��C�������U��u���F{܇��%UfQ`.`.y�/O�}�tM��ZJm������`u���C���QR`t /4�{g�#�n=U���\4=�D�}��y��:�B�Ft�)d�Z�7a���#���B�M��xN�-��.�O��L��_�M�;0�гs����RF��~��J��\��2>aVͳʹ��/meu~�#����1v
��c��RL�)mEG>b���d�\% ﹶ����e��L81�����KN�B��0�9L\@;v�yڥp��,-/�ʢ�Ӡ3;�[q�!�r2��a"���]1��-_ lC���nUaHE��깘��'�
D{x�]�������<�����Z��{"���Rɨ�ɏL�n9��T���s������r���}}�EVVV��;��!��������'�8?w�x�d�V2�W���K��d����M9��;H������>�M�Wg�f��Ddz�좐��*�܈��[N�P�Yz�I��	Q��Ȑ�yP�����X�V��>�\�|�wz-VN��PO�#t�@�wQM�U5�;{k�>V;q&�hp���;�VJvў�;������M�$���ן'9����=e��6SK(��;�u�J:5x��$�i\PL�B����Ǔ%�H@�!�EOJ�)׫=�SЁn��𿰄�_�韢��HI=��^���u֞������{���]JL;���ək�o7�,�P�NҨB٘�,���Y�G�`��.���98N�<�r�t4��ѹ��T�6X&k��̿���}a���ل<JA)\�5)���N�HV�	�I.�1lm��(�J<���٫�F�u(�'F����C�B���丹R�8ŗ`ٝ��yY��
����4ijY~�N0�X��3���d�Fk\�x���|U�2�q���3��d�9�/M1���2v���d�{=�6�qq�|��r�Q��=��*�.����d�@�lI�ku
��&�r�����N��wt���Wu��#�����O��hF����Z��"��2�S�5��&*T\]{�?jk�DIP�k�(
!��y*M��]��ʒd�E�mC�}��b d|��4MmӘ`۔,T?JS��w`�U򱉕%1I�\�� �tg�|�rB4B��i�o �����Xf��c��J&�*k.�����2���rt$��=��1��w�U ������]���u����#�!�F�����)!bq�/8��s���<�.�2݀ :g�%��qs'�i,��h�2pk ��)��$���R�1�\^-d*ׄ탉��|9�|qr�o�q�S~�Zx�n�tB�[���(+{W�Vl{�~��,�z�Q&��p�^�������N����/j���'��j.4�iF��w�k�k�k��6���e�Xo�|���29�&(��>%�J��*7�W$%�sǫ�`�1l�7�Ե7
�3��l�f��Ϛ\Tz ����̮-p$ޢ�z�!�?�Ȼ�aD��"��;*��uK4)�[�o�v	n��ڀ���I��v5�(+R?��:=d��1V���<��~ �_�� �.���V��\0t�*��z���++��gepʄ5�ln� f�5�/�������N-�:|��$V���e�NQ*������d� �g�*��N��͐�^wa����y��V�
�����n I��[��ce���6TB�Q��q�a;6�����?�L��in6�Jї�t&�cO� ����+�*�������-�j8�a�n�`E#�֟��,��Whb�Å�k��)[�Ua�s�ˡ�F����&�G�/b	E��z���Ϊn���..���!��s�]��+@m�Wʙ)�3�����]�Ai<�fx2���6jbH��Dx�_��%�#W[��}��n
��ݼȕ�QԺE@У+�Sű6?�p��J�*[����C[�g��Z������]�Y~��k���fk.]?�ե��J[Rjk�<F����-臊қ�@���|-:�}gx�I���
V#�ٱ_��B��ִ�W�~'u짫琢�]���7�qIZn�{�(�gr���vI�������.���-�ks��4�q@��G�Ӛ�)��tZ��b&kHK�`G�$�+�q�J�r����#�bB���׺��v�ם��j��I4�w�B�?UQC��V���a�:E�3�	w����5z
?�e: ��g���J���#�Ũ�9���w��Z�s9-�����_�۴[������7��ۃ"Q��&��	ו���%��3�4���|ڙ�@4e���$�?�GG�f�.{Z�,Ʋ�)����A��A|�l*Ǥ���Å�B&�������e�����$C�w�
�m�Fz��)@�#���C����V��۫��lSv�ɝ)�;��8;�Œ���D� �>G�۵c՛A(��;QzD���f�uD�fn���F��vA���ը����Cz�G8�_���<тW:u����L�����
T5c���e]�OfA ��r�R�Ʊa��}��m<�|sϼ?��x����əd:��$Wo�2cc������fM�b��rdӲ����ԋ�wg=!�6&�%ܻ�0��cYG����=c������������B�L�01�l���_�)��
!��U h���x�B~M\:y�+a�7�9w�q�i�X�jZ�����6r�;� 奛�E�P-�kuf������is�4	��a���b�
w�{koܛ)K�_J,���]�+M�M��`�U�9S��Af��߲�m�%f}���U|�}��A�AIy�<�Č�d]�}a�OB��.�K�F�;{n��,}��d�4or][�1I��*��1���wm�
?���Z��z�a.�RcJ��&-*'�5�0��Na����o�F_+R�����6�d�7���ҷJ�Y"��4kn�g���!A��:I��%�7�Qǲ/�\{�ݔ`���{'C^�������6��������L��c���s���>�c,�_D�i�b��淇D&GR���%~G���߹`�Q�ȺO((������M	]{9��� ��:�څqZ����n,}\Q@���@m���{�p=�� �Z�vb��u^�/ϣ�p�7��:��Y����FY@S��w-0P��Pg�^��o��|_���:��.����d��Z:��k>�:Y���||�'g��HU�1�f��z@�ϧ庸x>�%*��G͒��ee�I�6N�Nݳ��G�4��
���5Ka��׸��rg������K?�"�?O"<��u�?9�1��[��(�* ���Էjf(XQv��~Ζ���x�'�M��H�1����@��+��}��}Ș�|�YɈ�I���g��x����,]�Qv(��Y>v�k6����t�乚t��pP\I=?�\��'�]�ar��R7�7&��&O˓5)V��.j�F6A^Kd��:::�w�m�]�N���ҫ�^�YB��8�(�9��w�O���{>�LT���eƻ�*t�yd�.T�+J�a�0E�0?\r�~#m.�f��!�.%������sE}�G���15���
�b�*���N���$ַ�ws
Y���<'��(trL�"
��G�Ö����b�6��-u�z{{l3��S.�  �3��iw���y4o�<�C@"�aH+7Kq�����)�#�%���Ak��W�N̂A�J��/�}��/�"V��O�je:���[�9��L=D̑�C[M�0������x0v߇��I�8�<�-.׉G�EU��A��8-�)��cO�#��n�0��t�m
G���}	�:���D��J�����,a��m��C���B���Io�/�o���:<��Y^��xT���,a����C?Bm�T៷q�7H7h�����Ƴ��[U낶���hB��T:U���������H�^Av&���m'�pצ�iM��^?' Ԟ]���n�Q~�%��!D�������~�4�85�T 8yZ�c����'c�o�����}���J��~kdh��sӉ��D�-�L�V�ŏ�Z-�͊�,��n,�#���ɠ�!	�O���^/@�!�+Mn� ��݆�)�`��{ޫ#�ѧ�[2��l?,Ϝ9j�3@dݺ�_�V���v�&yՓ&^ɿYJ�U�Q��',��;+��2���JZNc^[�@�'�.�R0jP,z�'	�l�;��+���J��ל��' L?yQ�ݕ��/�RT�Аztf;
.J���X(������!&���	r�I+�p���w�<&���*Ӷ~��E*�~�<��v_�9\��t�u�
��bj���K|�b����9I��}bZ�_���of��A�x�[`�H�����Vٕ���1��5A��/�ʚ�Ѥ�8�Jq���z��;�t��h�)��du�X�[57��.�*�	P'L��p���}>=���dfت?�&�C��4��r�b9�g+����7��tﻼN�G����b���K��n<)��Vȿ6������H���+(�B;Fi0�c��a�.[��z�K���h��󘶓���1���u�ܛ��d�HJ��_E)%��K^q�����nU^���[�B�p�b�|#�/�;d���]�I��<���+����%���i­:��m��t��{����7Nr�b�
��V�'J�"�"&x�= ����m*����Z������N���F���B��!c����Az�4!���;n=��Ex`ּ�,\������!-�3��K�T<f�F��W$wG���1�"���\Y�w����j
��A���D=1�dP�Z?�jO����̧���Ŭ�Eq?jp}��ƌ�:k��U��ښ���a��KֵF��X��J��e
U����b0]x�5о�q��#d��Dm�����Q��Q��o�k��F7�nR�e�xTNG�GҬ[��'�͖��8̙Y�J��R���1cb�p\pϩ����(0)=�;��Vv� �`rK���r=�'l���v�8��� ��=9�k���;��(��+��AW�W谭���~�&M�$�e�5+��;�uG@"#��yt���ئ
z_�4C���B��j��(��'�\��������/rM�Q��#�0 *��U�ު~o�� cH�(��|���O)� �̟3�JR�J�k������t`2݆�Pi+x�P�*�0���z~:�\�R���S��!�*���i&��Apȋ�e9�%4W����B���rʿ�E�~��e\�^�G���tI���c�kz�L?���1ߓq*�;[s��%�4��,F��N)����g�� 10�&�7�lKO��²Y�R�E��.M���+���->C��6�"�E��m_*�~��O��o��ԍT������+����(X�c�g�88:z�|Y�4hҹ4�L�	���2�Q�3�OeD���~��8(�����GS���_ɿ�N9�+�k<�,�//�L��gӾ����U�^!��ꈗNS��;�Y>��r�{����Hf|:����L�4l����J�,Xg~��ĵ�l^��~h4�3�{��1?"&����h��Ʊ�T�_��Ӛ��d����]+�)ic%rrǢ0�-0�`X���E��#�տ�Eg�0ڹ���h�ɶ�5��ZE����:m.�E��mL�Ҏņ�R��:--�w��	m8��~����#Q��&kQxxl�N��<����01����bx|x8���u1�7�TB ZjE��Gw=��N�%%%M�_���{N.��	����r���� -�VQ�u
V|��ž;{.r;}Ԧ&�k��Qf��I$��f6��Q`��������W�����dO� V��>2��'���u�M�7��X>���|�q���:�f�W�\+�T�Q�`�g�&�vNi��3S#6���#M9=Ý�r�ί}�i��@�7[�ێZ���m����:%p��.b���V��ēO~k	4Znv7� �m4�l����*>>G9�ʇڶr3*�Z� ����Ls�P���g��T�wυx�ۭ��7�ܝz��f�>� ?,�'#��� (�ΐ����P����qe��4�Yr�E�2P�r�������Ȇ��}���3�+��D��_�6�P3���8��⪫���G�=�����O]�'q;�'�D�O���}�!o o����
��+1L��,���00����ɹI����OU41¹[����'#C��(�����D����ۋ�_�3�P"S�\�������A���A����Yz��aw	��QU�T����� PK   �i;Y��<���
 ��
 /   images/d75681bb-bbce-4690-8af0-fbed32c25461.png @￉PNG

   IHDR  �  Y   "���   	pHYs  �  ��+  ��IDATx�����%�q&葙כּ��/�4��I� �8�D�H��������>�c�&imfu�H#���(�� �}5���wgf��{�{����졺��ˌ��p���s����bUW�-MK�Q�nW�,���C�uo_�F�g��79Od��@v���pp$��TbE$�+�1Jŗ���-�
R�?������!���W�Z����j��^?�{�������fY&1�{�0�������=���U���2�OПs�k�G�c��V���p�P���^��횁���C�����b�_��1�����\h�î�_��+�|�&��������k�o����C�D�����C�}�������_�Sf��GLk#�>:��_-6G�L?��l!�$���)��i}_�r�?����]6ꖾ;��W���g��=�[�x�y����z�R%���G]�:D�6%L�S����މSVŌ�k:*���Sغ�ߗ�<�������>Q߷��[���}��Y�82}��(�j�oB�=[ǚ�������G�,$�|��<�K�;�*\��^Q��~-�ݶ@���d�M|̱j�����(8F�>���N�-����,�+ϰs(1�#���,�7y�q�M�gߩ�j�;�/W���˲��l���|5�=�.��]��>|���+J��Mk�1�w�]��]����o�����{̿�f�����5_k�A+kACr�I�殇ce�hv��_�7�/�H��962cv!��}�y.����Z�}YM�#�Tk�S|k�y��J�~�e�s�Qۊb��:וo���{5��1�����͕B=�F/�]���k�<�UO�f�oɾ����������g9��Ki�2�:��ٕ����~�P��G���<�+>B��.ym����B���mw��&����ϝٞ�{gUp�'����vD_�����[g��`o�,���c���G�ǌ����ʧ2�R�m��;챜�u�m�AF1F̄�"���+�$��O�+�6lJ"tl��h�ds$�ס#
�3�U��ئ\C�g]�-��E�K��xUU����/��oܳ��L %R|�^�u	�p��zU�~�H�����$�u�^��Z��x�o�b�7`Bb���^�L���ܒ��Y�:�H��6����4�v���e�8��� s:?�l��ޱg��\�7�8�w:�o0���׆7T��Z'D1���Ӭ�f&/���kJt���s�X9��O�]�G��m�cq�[�������\���#�F��H�� �2��+�Z��V����p��▪�4	3lap|�z��զ�f�7����<æ����a�6�|�i���{аX͆f>Q�==�CQ��"�?5z{կYO��sa�ןI��XHE�5�_H��sၲ:� [Ϫ�9�V��{<��ݼ-@�RNi7[E&��&�mA��ߡ��N���N���H��R��󩘣�s��:K:�U}���r�Ě��[��qt0��1mi\Ya3ݐ�J�H'��{�������;2Q�WfK�=��^x<�Ȥ��¢�����U��7�(כёJ��J�6qh�:�} ��6g���|��}�ch��r��O�F�fGW���F��dW27ƙ�L�c��e���2� :�KȪvp��}��
�Jr���$П��lB�*��̰���
Y!�o'Wr�YH�h�H�>��7�C��J�>�vrv�;��~�DP�v&亮�"���6�u�j3����\�Ɨ��R���p��0��0W���k�6I��2߰�+>�ѐ�۾�.'��P�,����gu��|.bh@L�� �}���@�$�:�S�&�!�(�!oH��4ph*����ʵ���Ɂ���U�Q�A$g�Q��"$�3�&�q���>p��c� (�/� �=��3Z� �m�ڿ��A+�!M�0,�`ړ���i��UY���I�U_ٟ��%�Q׶n3�1ƅ����9��Ou��8������f���Xifp�W��0�!����|.�!K���g�[Uekb���@<XF��^������YL.��}4���e��M������͉�j���z��t;xP(9J.����NZ��z�1���Д����=�	�c
,辤�B���$�����Ў���!����mZLx}����T�g:��1�n�� X4��`((��<<�WZKz�����s��2G�j˙��C��e�d1+m?�'RX���9a�Ak�m����']�jny>����y@�	N���7��U�Z�����A'�S>���#�	�v���m�������uA..v��MLa�\�-(|ͪ�1R5�YH\p
���q���m� ����a�c�C�c͒���o�V��R 4���V/8���I�s�{U�J�جM�t?�'7k
`�Be��4�H{g����ȏ�Y{&�_�u��c2x2�w�σ��Ε�Mm�I���}�x��)�B7i�r{��L�'4A-{�څ�2��<��#9�) j��m�4s�Ûe�h��wK���uMn����`-)���>u�t���������mNp�3bzo���΁,Үe���{��hr.CYHz;} ����]�,\���u1��o��{3U�%�lD�|&�����s\�cM6�i��iӻ���cm��{�ӯ;+Mཱྀ���t��dVf��BG_Ք��^�/��T��SY�weV�ro0����T�ϟڔc�ǚ�-��B<�2�J�#C��G7��?��=���W�p���&Y��vgѢ�Y���'3���6����T�0���&L�;��o�����Y���M�FF�8y�)b�h�B<�.Le4�	�]%����7�ǅ�Q�B:�	�d�h�����<@OR�Ɉ��6R�hl�F�����0� ���,.�hT�7վ0�\\z��Jx=Z����gX[�vc��=�J *���HK�\��k�i�ߒ�uRzIKp( �+d� �~t� �b�b�H��\L�΅��\q�YF�@�Ǵ��ߴ�H��GW���;��R�4�Ql)�$��{�&:��	�r%��4�f���+�|���
!���Fע>j�����B�8�)�M�Y���=�����e���A���i��RO "�h_ʞ�21@$	����eu_F>�� ���4F3jY�8�1�;��G�����3N�c�����̢�ef�foU����V�Ϙ���%2�l��`�	�?ă�s��]������33�������Y0�f�L!`����gA�p��lZ��R��$,\U"��Q2�I��_���ւE�	!��K���/�&,+h:�n�d��\[ZT��L����{��̳t�3$i~J���Kr���f��fOua.k����0@�v���FI�F��̲Yuf6N!t\H���?�u5�C��H���[��f�6�����M�bΔ�3���c��
�!�8��9��(�:69^�k1k?���lw5c�Kܹ��V�.����cwf	�xݸ����:*%	�eў���&c�{�����e��u?����	�>/�a�38"�3ӫ,��fm}+�f�[��U�h��k�x��19H�ӈ���	�P�36��E��09ѝ����4��\2���l���̔�V<�y`ky4��(dPw���!9��K)�h�(z Ԟ�(Z�mS	���i���(&�.���_�94�S�`�܎��s9itht;��"���fc��,Th�3H�>�mM �U,���5$�E��5|����6O�!P�؞J�8H�gDe���ݨ�:6v%s����8X��桌��\vh�6����_��xР?�ڃ����Ttɢ邔\��x����F��g���u���J�%X`�s\�d��d�A����N+�\�@8WA������,����~L1��_��IܹՖ��X��w$��g[��iɒ�X�����doZ�[���?��u��l/K��*�R03�zk��A)U�*�	v����C쉾ާ�-M}L4��"i!��e=k 7=�8a���&ߦx�e���������̣��.h!�b*?8�Lt������lv����0�[uF�sk���:]7�$��w�ӑ1�^Ǭq��bn��,�i��k��eh,��3��d�;'2]��49�f/9��u��y�"Rn�c���ߍ:�͍�+ؔ�$W����[8wfl��C��n�(�;�r�W�8d�T�'�HM�z���M.NQsJPrBr�%s�����F�d�O��1&P	j6����5��6{���y�낊P7oǿS�2z��(5�%w�t�]|�}�H~jS~ь$�e�sdΛ2����,ͷ�9.��V�-��9)��YT*S�b����H�E"\�=�Px��nH���y᪭����ō9����� �B쳈��Bq��G�=2f���as�� ��e6�>�oWcA���L��,;R�B$�Y�kӑ���,
�cTC2�&o$�yz͢�)������ܟS����"��\�?0U��X�}�AY��

�uV8�3'��^D�lV�Q�)� VE�D7�,�\wBG�I3����lR�׵�o��2Ƶ;!������Ie
BP�$G�t~+K����C�^�o�[���b�\S�"��ׂ.z�W���I��Ԯ4�R j��)�·��:p�SH�#b|3�L�0�8S]��|������ѣO�'3��) � g`A��9m?��=g���pcm��1HNK�q��4{���<Q�Ȉ1e�\���9w��!	}��B>U0ہ= ������h1�s�L_I'̿�o�o���Ì{�`5ѺA;�Q���,�cA<I����� Y]�˔���Ȝ����H#{���I�cN�Μi7�	v�<V��󚠀�͊Ά���Ra��j�4љ?���b0zp���r��*Ω%s^0�ͬ��Ӽ�H�N��y4��a��+9��ty\�)Q��GH���.Z��$�[侱����X�JlL�ut���s�Li6��Ȭ�w@{�vJ�$�g�A�#V�ي<4a��cb	��'|���̃�q~#y���#��g�#���[��`�.���46�����1����G����Tu�ꓖ�PPg�#��6�=�Z]�WW��-RCAL�қɝA-G;���o�}�tn&z�N�ä��d$��RS�����齘b�!��������ߐOn�H�]�L����"մ��p�������n�oDn�L����T8]�V_�CO|�?����<��` ��f���#6�,�G�<.h�:����	N%J.Rd$!]��nTg��scn�<k~�Kps��t{E�Q����Z���n�wȆ�kG'9���'K�Ift�SdBP��O`��j<_m� (��B�f��`*�o��v��9;�yCR�͞��#��4'�y���ً	�S�X@�|?��85���Z���p Z5��}ԆemJ�2g-���-#��T ��(�����R&:g����S*1�=$���7[��S$��bɸ֞��s�@F?K7n�	>�q�ɗ��p�m���
5E2W�C�5�8d��>�~^���w|�f�ňc�˴�"8u�v#�e�}>W��Z�S�戧��<TZ��2� ��)��`�i���:�,O
�@$[++��y���˩�+��{_pg%�����o2��A��YSǅ��@O�3f}��:���lV�Qw��5Bf!�F�p���2f Yw�@�\��b]E
�������(�Z��1�ܟ��;n�D$�
g�:�[��  ʰ��@�ȺH�?��H�L	� a��?��%2�=�Lm�e����S���/U�c�J
2�ų�:�{_m���3-�v;m4:L'��٠�����Y0��:�Gʊ��fhRMb���z�l�`"s�C����}��pt��wǤW��b�Sݴ�P��^K1�h�u���É٣�8��b���,�P�G��R�W�E��c( +8�����2��Μj�	¼^7eU,Vcs`�:Jڇ���%�j�Y�Y�{gE��r��e.sa����=������N�4�D%)�L'=9�)��A��@�ޮO*�{�������Y��N��	��,��3�)[����	XC�g�׽M	2A-�#����Vi�5����ı�ݲ$�ǧ�%@R7�^8��gD��n���չ��4`��M�x}3���F/J#Sg;O2�h��.�R�9'�K��[�Yi�K�t߹��괳��f�Z�#��H������0L5��y�4��?���d�:����H����x6]�t,i�Z�<�n�|��H:Q|�BH�,��{���u��dN��&��+Y@w��[c�!(Qx����9U����'K��NǍAQہs���)����<��Y{�V�5��XV�2ˬ�f�էz8��˃���HRƕ[ٛ'�2�{��=w
P?� Q��S,���<}���CFo)g1��z��lE��Z��Ñܺ�-�oܑ��9P_���I:���/�_�;�ʭ�Y�u�_t���-fz���_�������\�JX9�wIF����v��񶴪�������jǡ,w2Y�t�����h3zx8�eg<��#�Xʾ�`��3����(�uT�5g5��DՍ�	(.:~3�(��&g�U̸׼^�иk��
t���05Ц6Q�ǥ�"d���l�J,��� �5/,ʹ�O>��Z�����Hc�2f]9^��1�� �!�����(!�Xc,��<J�\�+3�5̍�|��TTD��L�H���0��4��ƈH`�x��7qmT4*��jp����k76��wjXb����rN a�K:ɖ�F���-Z5
�x������iVf�@��<�]J��t�����Qk�׀�4* �P�\��A�E�eU�i��g~��c��W�(T�_��9{Q�j�YC�+���t�1��s�ʭV�r|Y��e�f6(F�}�pG�R�2Wt$�ɱ���q7�� ~�����M?Z��Z� ��:�=�P9�.5$���,}�=�>Y��B�Q.+61�c/�������3�"�j8�p�E��g;:<�|�S I� �c��0��vˢ���إ2��gD0o�	s� O�u������u�Bc�@v60BZ���n�$N���Nb������A'��=iaϛ��՞u��d��]��m�6���V��ޅN.٠%���uPX��%��Ѿ W��Q=��Fp�	�R2s�K��L&�LqJ ��e���y�����T���t@�^R[�y��2M'#�/�tV�N�~�e��!{`�r���؏ ��Ι��,��1O`�;[�e!� +٦h��$@T�p2����t۪'Թ�R籶̥1W���z'��fNK�/��x:ӽ�Πd�؃c;Q�Ф�3���"�����ht�vw$����&��~E�j��l���p `Z�VcS��o��"�^oI�]�T�|Y�F��ԖJ�ؠh���Q��:��=�̽�5L&��c?�V�)}��,3�����@iR�|ea��E�ű��E�=�fxF<[�c�����:�R�U�t�u��
����tr��h��ս7O��e��]f�s��+gC�6�D*YH5������G�T��>k�ƃ�^{��B���z}]��C��
�*4Q
���1�/�{T���Dꊎ�kl����9�~��&9�ф�z��Hj�Q}��{���R\3�&w�Â>�>���C�E�7��p�@�O�6?Z�T5K*���u�᎜cd&h�>�sw�uW>��}��		���چ�Y��Z���
����)ϼ�L����%ɉ��*x�uK[�I��1Sg�^�$��j�u�t��i��ה]�^�t3�%lm�a�$�Q';����o��́D^ԥ��
�ڰy��P�T�~��/`c��D8�']��iH�1��R�=4�M	��F˹k�YO��~�W���x"W�J��&�HA��qA2]�� �:&�X���y�Y�1<0GnG-M҆�d8�L�5j�D!Dw��(8���n���h��4�I_��OGknS[�B֢�bC���c�C`[�և�I�~szk�[s)G��7��R:��|�T/u��<s��<����Ǘe��:D�g�+cϴ���lyI�8yB�:wV���c�����Ʋ|����W�ޝ���p �#}�����>ѕ;��7ޕ�ߓ���`O�k�JD7��-U��H5z|�'gO_����ڪz���U&��Z>��#o}r�������V7�R�?����UM6E����� 3'��d(jLRe�/k5�TG���&	E�8EgŝDs-"b��UX���8(D�F��JE(��[�#,��ɹ����E��;�b���`�xTf����3���U�xiØ���C�ײ�W����Q_�����S ȣ-��3�#��ZU%����H/蝚nq*I��4�}>(VD�f!�;f%���`^+"��:KF�B����3�	a�!R���~�JnV��!)Hp|�A|��G�>3�׭�j$1�"�i�*ݴH�e�h��p4���,o�O]�z�1�[�h�������Fh~�;V�>���QPֆ;4���P�:�n0�s\��M؁Z�/]�;���]Xg>f�N�X6��J��vn�ҝ;wt��\_����	,dY��A	d�֮�Q�JNh�IIN'p�{�T�S��In��W�xx�u§'��*sA_���N!dq��)��tMt���N�3IH%���P� Cp�-�"Gg��C������� ��AE�8�`(�I�=4�j�{:�UY�^��x4�� `A1��P�cFfF�����>O&���.���2I=I��et�� �t��:'=2% x�rJ��{c󘾯%�I�'��`�0�X����0�F�����eP<z�G0,p�@�F��ۗ��{2RǢ�����H���ʪ�9�$J��%YZߔ��ΒB�z�ʣ�֙2E��\�������N�6�ũ:�����X7�7��N���Ir�]������(���:�r2�x��GK��t�z�e�G˂-�t�K5�ֈ#� W�p�UTP���w���s]��m���lL6W6e�@�~ɂ��g��*�;b,x��k.sZ*k�GF���]%�XN����tx#���.��i��c'��W�����t���x�vUn���=ە2�!��q-�qʰ0�f��Rm*�Z[�h�6�rX{�	AƩ:�Qu��pGEo�5���5t{�_���ڮ�S}��?�s/K/�3`�2x��أǥ3��7`:3q*{�t8��YG��\��^�]�#��䳬�DƊ��Qhh扖��:�T���~E��:���wu#�+�(ԩ���t�?~L�BW���2`��>�D:��Di��F3��}j4SN�bM-��U��u�+�V���ϭYXS����2���.Zn;Kk�{��^@Aml�1�r���X#85�=2�h��j�#dƑK��Tv�MJU2��o�V�d��� �To��nа]�[sf*3������BCME~�"u��(��mx7%�L��r�,5Mѱ��F0�`kuS���v�gۅ�;�@V���Z`��q�]+�`C�g�(pg��.6z.z9���j�̏%��L�]7�^e��"c�2˭v�A8K��+v7m�co��+�b��Tq��V5��Zƺ�1/Ȱ/�ͫ�\J�^�/Fca �C�X5cr$��Ah_�utOl�GaܔqM7^d7�y�)4��kL��?ƭ�An(R��`_�[�0���j�����gІ��5u*]"�d�em�-O�9.gW{��ZA$Y�vʜ�R�^��C����i={�s��嫴��rK�NE����`�o�ۑ��]���wG��������ɖ�%�W�hV<���9S��Tw/����|鹧�g���Ǒ��I�fa�*�O>vRNl��r�g���-F�fj *��
��)�e�jF�kW���^��ݤ%)S]�!�6a䲴,K�) ���b-m��;�լQf�b$�N�gK�a���u!�_X6a�@��^�O�*Zn"hq�i��E<+_��P��ϊ����b�'*t��(h��ZO��C���oӓ�˜�G7It��~E3Bf�w�F�xϑ�YV�bp�3��a�h$"��^���"���i<�yU�)
��.)B�N ��#4�AFb0RC~t��#�J������X!;C]��z�ݴ��珔����WjlJ�"D*um�j`ID[�QeYT�8��[R�ք�yf6M��0e��<bl���>�k���s_�z�1��L-�#SV�%�#��K5�ro1>T穣���wT�Ki-mI�t�j�Hy�VEa68.�����x��Эua��^�,-�ǷN��ም�uU���D�ٌrQEys��u�U��Wb��}�׽�3��̳�O������϶��ey	}��;�c���N�p��C��
�M�Is.:=u���8����T��T�H9��C�g�X4t�4?��ʬ�- �GZ�������D��g�o��t����P��p8� ��ts�@Ƈ:o}���h��M�����	�:��V�봸W�v��J�+'On(�ʕ˗��mKm��9F�j��gDSm�Rv "Z�QP]�`3��Z�gV�Ƭ&�Ec����Sq�����YYVy�Sx|�/��Kr���P��ړḒ�?�L��oJ�]�N��2���=(���:^�:"�ާ�!��6��[�#�PX���iZ���� C���tB��=S�=�Cx��S�؉g��ڲ����x\ZM�;������|t�
�[]�KD�r�n�Oy�,5P�����G�1C�P���œbo���\��r�̓*'X�}:,��0&���-H!Yp�>�"�5&HA�N���ʚ���K���*'��ˉ��2Py)�]^Y��?�T��������T�i��Q�'%(r'�:sg�r����S�%e��.2�(�-(��h�8X�@?�C�ߊ��l����\�o��������!�t���ѩU��_��T���R�C���c�ڱ^���C��l��u;,x�Y}�������3�����-�{��rl딜8}N���'�©�sƠtdР�sF	����ڳ������@���d��/�
�_}�Ey�⚮������h_6�����e/峛����>Q����]��̆Z��D��'�1�.�6��rFg�` �R9ʙ4���0Y�A���ڌ�#�����YE)�=yVN�_�U���H��[� ���U9�i�}��l�Ӎ{Mu���� UC�df����U�m�����޽#/>���:uB�^�&�^�"�����eCdTۊi�����7)��!�mr�4�൙���hA�����dp(+����pAVW:r��� �>��p�y$�������u�.K.j�,z�%���75�^&�@�����*o4�H)�d)��ΐ����iF���F`&�dK��v ck���Ǫ긎꽡�Q#�cWS��V�ӑ`s���,��ڤ`#��A��%��o���`���B0$�$k���7��2sӃ�*���r�@�%�p��J��g�eQܮz����J�\ cJ1�H�|_rBU�awbtH�/�KMgi��^���r��ڔc��ur�1��t�h8?��5=U�}B��ge��x�P�I�۶SΧ���p$�������m����F'�L��j�/]����}$q�#_��|����rRAphu�J�Z;6@0�JK�镶t�y\�>�N�ۗ�K\;��x��PA{���cdݰ�'ɤ�-���k5�Q�r0r�$��B���0�lcO{ϳkt�u=�Vs��n�	�!�: "F<uS���W��h�y,R��`Q%�yɅNme��oka�j�-���o�s59�n�S!�7?P1���p����tU
-�,�Y��&8w�R�t_i����l>�~E�H\p/C��X��	�A%H
d<�R��@_�t*T^ږ��Ë���0|���IF�31u�Mkn3��sD�������{���\V��F���R�4��,s�ϟھ?�
��^��n*��.�:<v�*�)_+
�1���p�����}$���R�s��^G�������/��}-�j����G:��@�8!��2[O����r��'��r���p Z7����Ǵu�S9�{�S����P��աc�L�gȱj�y�1ĸ��m˺�o��Wԩ����S�q뺌�Z��AᬭFt��N=�b���h:��B� �QDk����'�VF #���k_yE^x梜9�N�|��֘�<���߶֏.ߔ��oU~��]RG�����r���3D%	.M/�s��T�=�z[S�rZ�� Wէ�E('|6���Zã=y�Ԗ���mq���@����;��Ho�������L�ww���H��<'���"�5K�h��>-Ҳj��ݖ�:_�y��?������_䣏>!Ek����O)G������1�:�ϚC ;݃�d�'͆�07@i�j���a �7ԽS�X�y����w�$��{����C6�bN�>����V����������Vtu�Y[�[nm�f�p�$��"��h�QDF��~�kG����

kh�(k��9;�0w�lĈ.n5� �/?�|�O�IE�mխ���;��|zG�Bu��^�*+���n����25�Y�l�!�{�yZɦ���x]N_�_��q��!w�I�:�g�{��*� /��I
�&�jA�$H��T������1@������ȷ�Ջr����z�k1V�{<ܑ��<%�F�\�~]vG
�t�ۈ��̞`�ؖ�Hn��	�D��'��\eAIPa��FFͭf�(�|蓒;��q�G�T~����/��[+|Z�eR�u0��Cr73��?����P�FO��q�(�����!���k��fs�x�3N˿���rvkM����ܒ�vP�yK����Ef`fmfz
����h���CXhNe��$����>��p<���u�|酳����#ȬZ9�0���>s0��o��߾��w���f��L�ě���`Y�t�_�Ĉ �=3�W��1�(�U�&fF�e�em�1���?�
�_}���p���+��3 �X�F���Wˍ���ݩ�.����'Uj�d�A	��NeA���k�ګO f*���<����sg���p	�^wx�Nf�o��lD�����y=0�_�fzψ��[��7{b;�N;�����Y�W^zB�8�"G���(�l���x�h\�o��H~��o�B#i�$��M��E^�3�j��Ӛ9��Ϊ�_B
���}��98����b$�F̉+����9<��%/�~?��V,mA�=�'`��+��,�O���^�}�F('##�G5�i:cXc��flFY��uTן>q\���)fw��ܕO�^��IT��/���+s^��6���� �HB��E1�җ�@���o�Z_��'V�d/��%��p9��M[�� C�H7���֭C�fy�9��;�Ĕ(����@*?j��aK�n��(��L�:59"��{~��!D2u�؉M��8n�/GHf!3� ^i�nc���9�1)>TCt�ގ�VO�f*,ځ���z����ޔ�^|R���"�+x�P��̙.2!m/0��tTTh&C݄�����A��W���#��"�\����R�=3r.��Q~&�C�Ɂ�ء��!�?x��(��$9��t�H)���5�S\i� ?s�7oٛ�)ٝedE��L�h����M=}R6�GC:�-0BQ�
�ʘ�ǌ�J�e�q|�E!N����c���z�]9T`�� �,��wH�)z+��s��g7�a�'��:$�0)������`-��[�`�q�z�b� ҡ�Cy���<s�)�Zk�.�!Dts�	�F�Ȱy��+��t�V������Yt#'J�_�槣C�\��7��3/���7�ʵ��?�f DsH+�7y�W����9$%�!j�
"N�=-���+j@��VS�c� x��QCԑ��C��;��?}���*�޲����#���U�MI�*��CL{�%�d���F{v �p[.��|�[�˙�ˬiAres\�~��pl�r��o�YAt���U�l�՜�:5hjje�#�j�t���������[rr������#�}��l�<�J��a��Q|�=S}��q)�¥�
E�d����y�wܵ��}���NO^|�	y��tu��]�ftzQ��gV��z����D�+zYS���d��L���_R�*xփ��h�6����4�L'/@V��f*Ȫ���;��3ؒeY�FK�J0q��D�9f�B����^����̮F;��iď��Y��s�T��x����%���	����#����X~��wI��8ƨ�He ฯ:	��
�)Ԕ�={F��ޔ�O\��	��QP��T��wp��d����r�B�Q�8U���djkYQC�Ǳ7X1=U:�"�c.������k��ol�)�p=FV��P�S�,�T2��r8�I���Zl�c�92�?��gNn������'7dymS�l�����L:��{�2����۪��Ŝw\e�������駛�n���L�>і?���j�W������g�ɩ�O)S�]�^3Z��)˲9��Nt�|�#?��b�:dfd2:<b���a�ϣR�Bu�}2R����}rcE���L��t�]��*���Y�����M6=���N�Ϧ�n�<��N�YF{u��������N�S��:XyU^��Ʋ�,�X���Oݑ��N�^�@��`��m�������`�#q��e\�F��^fdD/��s��=�prU^�ڏ������~� ���t�]u^r�5g�����rj�T=��r8�eL}������
�W�_�����j���B�4\����{r�䖮MKe��>��jc�Dk��j���V[߇6~~ZpƐ����%�޺H/�iK8w�u[փ`��j��Zk��l,��V��ޓ%��H`�� �������� Gv�����Sӓ��&���T���u���V4��t*y�ٓrl�+�Ͽ�P�~�#ńYZ;�zfd��b0Բټx�ڃ��~d�֎��nI*qg�� b���K0~K^θ��JW_��	w��za)Q����U�`0�CeA�D5�bc�Ɲmr��ڨ��j{/8��%|�ag�AUP��b�u]�K�7��ew���Z�3�	g5W9��}��26��NX .��{�ͩ�d�!�6��&yL�ʥS�������y���C]Õ�����O�6�6B�/�?��9螕1@��`-��S��ȥ�ߊfÝ�O��)�s_>�}(�UiA؄_<P��>��D���{����,kcH� �>���M��[(�v:t5�:��괞�X�+�G�(pj��?�2��S�k)@SAt� �����X�{W?���9/����ȥ�'d���aE��n(6(��dB�RիG�N�d�J�ߖ.=!�.��_~��,I�kN^L�[l�]Ńz��\�����Hk[�~�4�{�0�-�}�0���Ҙֹ�ïߔ��zm�Ќ��L\��1 ���}21+Q������Y��K��`�@~�����>�o���03�-��I͈_����ΏdHYW����d_�� /=A���K��u�c�Z_bTlooO7�
����݁�����'7��,���Beܤ�Ӹ�<������f�[���L�X��s���ۯ?���Ț-R	tM��ݪ�@d_��/_�K�}S
eڎ�-��qg��]�-����Yޑ3k'TF�3��ɹ�}��N�XW����r��2ptG=_��,���/��L$_k�һ
VW��H,���Q�Oy$U�9���s�E�,�O�����(�*e�������l!�̔���7'����;���tSL٢���+�T:��v�e8(e��D?D��l�ܵ�%�ohB�X�8l���TP�SK<DYZ��x<��߿-O����+ϰn�/�f*�|rY��'U�WU^�w��� �P2<������Z|�њFG.f���c�Js�n�:�[�vum�r��M�"�����/��s����6�{��)롌�e$ؚѤ�	��ſ�V�F-fa ��p4`#�����T�Sc�5�AC�h-�kF<�;��:��;f��U$?�����������*PG��He��hlzJ7PG��N��,$��3N��cutMG��Ou� h��@��o��=��ן�/�_�ꏿ�*�{�c��ݑ @�����Zg�8�D�6��|'%2�חW����S2ڻ���d�Qe��A�{*�-F��1BD��7#�>�D�o����Y(=5n�jS��)���,�*G'��꼁��tV2���ֈ�范�� 2�����N5	c���.k�*�F�����:=g{�c����&c����N��s ���w?����m�#�{��^[g0��u���ڄD�̬�Y4�a�L��-69���^��W䛯^��_~Rvn~E���'7/�#���R����������P�(���l5,��=�P���g�ȟ���K9�L����9�nK_�����-[jF�gjdz*a���L���;{Y	�-�5jDg�՘ڄ;����ZΝ;��~O�ܾ#���сG�/u�O�FM������(�2Y�w�`(��?�_���Į:|�%uЕhN�z1����!��l������u��� ����%�j���_HV�7��<��w��t�w޻*�\u��I	h���%k�Oh��1լg0����׽���������W�|�]Y)*9���P�ݮ��)ݧ��#�<)=4`�N��LJ-3<8b5�ֈ�n�cjv���a�D?�h-43��`�C�6t�+��$�w�Cy�G_�_�����z�Ա��})s]3Ş��#�%�<x����+�^�ͦ"�w׮ԩ�J��տ�~T���ߒ��w�}:G�-y���r����P��7o��x���͓�A73���BS���ߥ�훀GL�I�������=��/ߖ�W;�lz5�jO��rGq�E9��&k���q�Hն7Jg՞��>ILͱ�qY~S}~e���X��yW\&\b�sls8��H1b=�X1�Wo�u���{}��W�T�������fg9XnV"s�05�R���`�G��_�U��ۨQ�M~����M�bg���M���N�n��d:d����7>L�?�P�9K�T�w�f�w���#�a�յꋃ��������G�4�8����宜9�!K^��������Vm�	��u�?�"��33"�-�۩�U����y�"u�d�Ե� 07�}F߃`�Cd����
�Ol�ɭ������Ń�:cޱ��޾�������S��F
T���?����o�xI^x줬���/��7��.�z'
2�_�v����|l�//�����'?S� �յ�c���y�D�ㅣ�Z�����������/�c[��V�ܳ�_��3���Oj���w�޽m��"m�o�I�6��Arݠm��;��VC>���U �d�x��?�Ƿ�ڽ}��#j7�2]���8'u6��>��4L�"9�읹��Ȥ�Y�pW� �B޸vE�UZ��
��zG�nO�m�T��� ��<�_=eM��S�/pw��x��fܞ��Z�dc�X��'(�V!Ua���M9ع�F(��6���\�rU���Б#5PhvQ��M������"at8�B����]��w��1���^zB�B���N~��U+&Vp����
5�υ�L��#vIE,���
a�ٙ�l
@�ů>�~�{�h_�t�V:-ftA!��׿.�]z\AJ��"�Ր}��W�u%�S�摨F+/�l�Qd��(�o�F�{WD	i}|���D;�	j-Ёڇ�@DQٽ}g_���@n��U`�J_����:6 ؼ���\*�b�q7��qh��7ü�C#L�}i�/��=��O"�0��|�y��/_b���������"ځ3�t��S^�`s���"��.��D*j����n�Z�����E����ǲ�}�T�Ӫ�KuN��@�c����i��`D��t�JD��;Df�э�GĴW������W�M�!�@��Ғ����� sc�׀N�3k�T�1�7/)��@������jIT�@L�*ޖϮ�V�{��D�=E�/���{��Q�/:}u��	u���1��u�ͬ�]���j&��LT��!�F���P�{7d��c��+/�7�;'[�*����R~��7�Iە���*�]�V������*K���tn�޸*{wnȾ:�p��;�un)hP2iT�@j��D�f	C����2=�h�V���~��<OT����S ?��wWf11$*:� ��w³Hy���noI��%F�f*��U��mR�����MS�1R�4 q�-��Z���V�XZ����ё�������Q����Q���io�,Q����l�nP'a�̤5�c7%U}�_�v�SR3�5�B��#��cr�Ʈ�����ꚼ��|��X!�ß�m�OY��ME
"�~� hQ�-~`+��7<�D����Z�.�R��&t�ѷQ� [�F�mՅc֮���׿��ڍ�E��ڨ�����i��� V?g ��y���h ��c���΀܁�_46B�%�d�%����)�y=&�6�HW���Աݝ)�J�ԕ���A�� �+�I4��Ugı�D���T��,�0��3q&�����:j�
����.��^���|�̾�mi�_�'W��֬�W��bwL� �#��!�Ĕ�SPL��*��g���G���|�}u�dIu��GK�n��9f�!�%�����uoL�Q�T^�0'g_&��찉V�Y�9[��$����N!�l<���dX��-��Cp	�~f����{Rl������@�|�C�5}?Je�e�U��≢ӧ}FC��������붏YWذ)g3Ba�	c��S31[
v������w�N�*�_� ��X�o~�U�����S9���=�F6G��m�`��L1���������7ߋ	�v���2�x�\9腀fKj���/���~��)t�>A�z����W+��e:�$����)UL-�D�z6���^̣���B� �����BO�=��(�#�ŇW�i�����)�oP׍��@u.:`��4�.�M�A�R!#�)�}���?�[j_~��D��yy��)y����
y��k����rkgW�c���-Yrt2���K�u���q0c}� 0�7��3�;����m����^�vk�MϞ>)_{�%9w�M��.��Ԏ�o��a���ٔ�jMq�aW߰�2�E��N��I��T�r�j�?,�0\�Jse�9�\YR��"�m4���E�r�l��P7#".X�0�btz�'��n�~U�n�u���t����$Wr���7��B*g�>��7�D+�~��c����N�R����m��]�n���yC�"��TAU!'���Aj�[�},��C��Y&�\�4U���(�t,E����6�֖t�Qrn2Rg��+hF����r����\�o���������T>��Y�ܒ��:j��SQ�b��&kP{�����#�����5.;"������U|�uxc�߾#'�Wq}I�^y�Ŭc5�u{hԂW�	r����"�^{���vnc�y��3���8/����*q��)�*�'֤
�ݵβ{����'?���ۺG)H+B�RA��p���nPXt��(l��n!bψ5s����NwU�԰��/ޔ�p(�-U�Ϝ��H�����[�Kgy]�N�W�n<��!K�#�6���\:B"�̣�-ݔPҠ�.
徻} ���骈��x��ݻ��l�9'�8-j���h,���' Tɬ`
�NIʔu���P# e���<2�f�j�0ZR���4�y��~6��^�Ӫ��&PY��3���Gr��uW��j�
4&At �ôǔ�<�[�s>�.�5�`k~� �p[ݎܾyM~���HO��=/_}��(@�O�}���M��C59�ѻ�"��f.�r�Pf��#:Y��Wl<���f�G�r��w�V�po� ��ɤ�q8�j(ׯߖ��#���ñ�	���1���޵l%qj��f�y�z`0<2��;{�1y���ıU5�-�9��jZ��3R%Ic��V	�?�a8e�X��Ddt��z������3�'Bd�Y.����(�y����A�m1:>O�	a���E��2 02Ը���c3�a)��H�=������W����7�F1|���ew�+U�N�,�ãC�v�Qafs�C���H����И��*�tDz�8�v�Y���y��Yg-ٿW���)��������w��m�sI�4�-��_����E�K�tggO�޸�ʡ�K�  �Gn�ζM"�Bl"����x�(cأN ;f�o�	_KT��˧e��9�l@O��~��@��Qʚf��QO�H��Jt.;p6�kcuX�@JG��߆� ����[�'����ml�����u�ٚ픥����Y��B�9����%Aي���"Z����s�V@��@�i�#H�ӌk�SG�>t�Ś�y�F�{tZ�Ӫ=#9W�v��żε2�ya��wn���N�SutP��>�Wl��5�BP���9P9B H�����Q�FO�$��p�֚:�6:�N�qC��)�i���� �G� ��I��kH���9���L1�T�����s������o����U�O�˗Ϋ���������}Q�"�ЦN��YG����3^��B���g�]`-lI�;���y/��Oٞ~Iu!EMG#�"�do;��~��I2��W���ae�{�?[�]%�i����(,;� WwuM>�vM>��S6���}��멂>����5��a�s��r'�V��))u�с���d�N�N�'�f	�@�1�����Dv:�NB�NzM���v����GR!C2����#��讽��/w?ە���Gߐ/}�K����j�^c�ҷ���c@0��d���T����ǚT��tS},i��:I%3O8%����Q�[�xPO&�As�єXx2C�Eeβ����X�JK�,9b� .�	��eH�K��鍕5�)'�W�+v��0�gGQ�)�c��q�x���M�k��rZ�oDS7�L�<R7{��=p}�c
D��P4׺~��d��[:.4z�Ժ�ƹ̎Fr�sU�?d#�����=�6?�&s�B&�S��zjaM8=����T��9���p�F�R.
3x���� �-p��Yx�kPL{�*[G�U���j�Z�E��X�0�YV�y��c���e����;䲣?�ʥ��Р&�N�Q_���t��Z���
���BTg6F(V���rzU� =G;���-�p3Ӗ;�bje���n7崾��N$�ŏ��AcDX���`ّ�{H�<#���t��@�L�MF��
�?�rG��c*Ēh
�l=R^�)��2'�gJ�w,�=Bl"�FKRE��
�oޕ�������{�=+����0we�wS�����2]Z'�"}�ϫ�|��j�����{����W1�&]�k;���;�m��ć70�AKwM.>wA�a�N7�؁�0�y�3�P`�����;�o����<(��"�x,���a��ik���dD9x�Mv:r8�H�A�$D�?�qO�쌥����`K�����Hnp��G�2��=
dZ��$ n�h(x����BW��/dw0���W�YY�o~�Yyᙳ2�޷Xd�޻����M��-�߮�e��]�x3AG`��3h|n3��17��n`.*p�פ.Jn��`Wu|��Ԣᜦ���]���h� ���Y�R��c��T1�`�gAW�.bpѲ�Т�0O���K�>�� 2A)�� ?,��b���UG���݁�5��}�,𘏥�c�
B?(P�7��TV�W������1�yf$e�Y������$ܲx��6W{���&ׯ]����
Z2�ګ�˅�g������Z�y�c��%��P[mm���`ʎ`G�T�#N���ڠJ�sc�����u����T9�(����%m�=�N� V����r��e�ȳ�@��0v80�CS4�Aֵ�Q?7��k1{�w���y��19{|��>���-����g�1�/t^��d�3�xGt����Qe�-'��ɓO^�6�3;ג�`C[�,H��7)͚�*�z;F�gֵR�A4m����J�����k��L+��qB���2k�ġ3[��S`%/���X̱BFw�k8M�)�4��M-�X�E��<4H���t0��q��.��'WN�����������;���%����ϯ�^
Rj�ͻ�ZxkoW�+�t���c���gs������9uӂ�� ����C�UQ�έ�t�/�HF�����n�^��@�G�T�m�d~��"�Ox�S��h����lh� ��&tQγL���_�Vv�y�ÿ��|�Kg����'?%;o]�}���#h4P��Z����6P�+�O�ߜ���G��\���a�6z T�X��kCƶ��Ɲ{�T?�W-���}��M�[��;�aб��f�p����������B0���z�٧Y���;��}=�o���<��&����Z4�b�
uW�߂u�=~lC��<�';�����\|�Ea�,����n,n�ʨ���������� ��t8a���D-;�{b+B~Q[�V0 l�Ù���[Z��}�DZ6Nƌ���7��)��&�u	��d�
kJ��;b�u��x�
�yk�,P��-p����k����פ���3����7���/	�q0'�Y�X��B���c� wT���=���%i+F �os�/���%Y�!�]#�~UiN�A��l���=����@�:����� �2��n�B�A�q8��NPQ[��@yO�#|
�'��(�D��,�̋y�1�F��:2�mٽ~[>?���Y]�W/=%A�lwH��.�%�!Fs�*�����RP�y���i�-���!7<⣶I�G�������Q�1Y{��8^�*�i��L찁n�)D��Yew�R��k@�A`���^�U�,<f��:(Ǣ���l��.k��r�N�T��PZ�tGu�&(�п�u7���V�K:hG���@q������}$Mcp�-I��K�]綠C�PY2�FHa2����Ý#��2��zYV�Kr��i�o&���͹��`�7>3��Q�B����>0h��b��Ζe�Y�KƘ�ϱ54����L�{�rf�'++�L�_�
�?�UH� [��N��e�U�۳\��DF�@ ���<�CbS��P�ƺ�U�r�53�B���z�Gt�����8'QG1P�\@h2_l�������҉�� sQ�s����kP��
�ݹ���g�e���?���^u�=�^�����$ꐚ��vU�hu�����9��}e����;;�*��G�7�!}�Aj���G�ߙ���휍��5w��_��>�%?.Ũ������3�i+���%�������t�D��݌(4AK��)譙Sg�y��㈈8���E�ad��C9<� u���uPz��T%�u��4& *�}����B� [��nq�.�Q��y,�p���3��a�2��*3�9&吵C5�RٹAH�Ժ�۝e�9�F��!Ã:�\S��	���m��������p��N�L��8��ݔ�����Z��� _�tQ��-��L�x�cYު��b�`m�Y/힩��`D�m&)��"z�r!�['����3R��_B��vOp�6�XWG��#�v�ʈ�^���Uɺ�r�`��aCГt���tA�����D��QGs��ը�(ʶ:$��2�ߗU�gę��zNФ���ܹ;"���W^�'q��6��6uP�Cv���.d��\�.�x$L��1���fu���ǣKT������[�y�_ސ����*�㔝1d	 �x����mJs�&��a����+�0���c��X#̹�<o��Ȗ�e�v�����ޓ������ۮ�p�H^x��lml���xMD�IO0�舛�>ʗ��{��(ݹc�Gt�PS�s��
^�����{�~5�m¬�8�V7ųC�@��FX����[��v�2/-
�uB ����!�.�D�AC�"c ���u	�2h�~�&�sV?47�ڲCxNd�c@3���s��G�3�sT�X 8Q�艫�{������8֖��.�؊��9ݓV���t)����������-�k5-�\��A,�ao�Y��C͚��Y��B�gq�( ��IyQ�`��3�����Ay'`w�iM�˂^'�n�-��p]8���o~[�S�%<��ꮸv�KE�N����@&�rq���&��f�AG��`Ա+([A�N�ݹwO�Z.G�c���,-u�����-����(Ga��>�ZHn��ұ6嬒�s`��|\x�(N�<Kݞ��i��D�S5[�ܓO��c|%p24�.�+��s"{�r<�Qw�OJ\����\��&�3988�C����Ϛ��W�{L�}F�I�N�eMx,�M�#k� ��p@y<q�<�����X,����K�Lh���Z�3�,C̹s; Z:�`�T+;���"}���(Poy�q�`W^��)�j:v�֭��Ch����^q6�co��|�cڢܓ.������e��L�������{������0�����fWV�"�t�]8�!��d���5%]kstO��'��ӧ�����<�`8G7��1zй���z�f��$K,�;�\�� }�Y�2=ݣ�"zf4Ҍ�=(�7�~�܃��������"�	����f;�Z�� -���ܽ?�f�ʕ�t�{?z�	Qi�/���sO]8(Lzq	Le�B�V�
�B ��g3�� \M���Y:��xY���;S���)��D������=�ǀ�Ya}���T��t
�5��i�o����ZA7�#��/����Rz�6[./0�9�w�ޓ��X�xlρy���Bc_�+�eG���q�Uyũs(@�K���ٹ&� I�����[�j�W�����5�{6�������d�B������|t�}ypk�>9 ���\L��XK/��1S@v���SF�+��̜U-���/J��0BH�>��tF���_S���dgi{T��u=�[����>�	�L�Ăq!sU�f�.ڔ��sѧ^�%е[��l~vW}X�j�|\�����Um�� C���~ xjqy �m������t�M�6(Є�)�� %�� �Z���c[�N��=GPB؋�d��́j@qm��� �M�UA����E6P����a6[p~
;�(�Ј�+$���-m\�q�S:��C:n.�~=��S5"5B��׃���g�|^����i9u��Z��r��# C�>"�A�*Y��B�;�����ߑ��u�K9;�[�]p�	��K��V� U5��1�8^�w�7�3tcav�x��r>�;�a饃�P�6��k.3M��D�YF�Fe9�9z�PD�X�NS=����ϤT��L�BN��N�m�|Q�ih��U ���H����.�t�\���bq���)��JqRQ-Y�*	"^9?��e7���!X���3����eg}]���r��M���.5�o�%�T+�`�A�ϵk5�Σ�Q*܉�N툫��:�*�M�Oj���Acs�ϥ�j�h�J�ӗ�7�wȨ:�u+$�H�+��H���{yv�L&���tѪǖ0�F}��G�Y�C�j��ӳ�m��V��F<���z��laU[$fI`�e9����9����@�Dk�f@�jX����E1Nes4�l�+�9�!UA�*{�C��htf�"��X�	�G�G��|x���{�mɒ3����1
��KYc�`����V��.��K`k�ѩ�	�Tx��`� "�X+��A�\���S"����ϭ�Zb�s�43p G׵�	e�w��d��IwȤ��| }5��!�ҩ�r�~l|��:�8x���bgpx,f)�o*����h�1Z��R̆ɨe0��R�8/��Y�*zdU��e��b�?�s�����fs��,�����2���Hѱ�6�1 ��K<��m6�v3��s�iR'⥁rJ�I:Z�4h���x�,@��X�PB��j8{��l�W�=����G��1B`�`��6 �-s�!PyЯ��ݮ\[�*�qN�w��O�[R�] x��{6�q=�����_~L������+���f���I�km��J_T0�|p�3���;Ao�絨���A���K9׿�����"e�fsy��h�5`���j�2u���|��ʔ���!�Vפ�S�<�gB�ણwa|2� 6����f�mNL��� Ul�}�S�"���/M�Um��W�?�����9~~.�fO¬%'��_˃k}������H�����6;�L°m ?V]��;�
�5�U=Ȭj���Cٞ/8�%�:s�����c��3���$�����*-�40��mN��#0��Q��J]jި?�Xa��غ�˜-6H*��{ �����^(\)r��dV1�7����2�9�QYu�8���>��d�Ӓwܓ�ӑ\ �T�5� �tt)�~���5�r�Ɩ�k$���"n"����@����c�Y���O��;���0*���}^XeL�y��0)0�/8��B�s����3���z}C}�H�_�̫~��/�YߐF����C�W���6fP�zd����$��M������ ���^����Ϗ��S���gT�d�����+UbƸ�k�5w����b��@�i�8��ǚ����G��%�@��M� K����oQ��������D��1D���A�l4���7�U�Z�|z�qch���Nƴ��C6��ajY%[����Tu��zJ�[�*)��H̊�2#��]*��mOJO*��j�s %��Ϫ���-(=��7���/0������l]���@�֗���=����D�yAc�p����'�v��(�CC`<My~�36�M���b.Ù����P��Z�ԉ'�9
>�b]� ����}��$Fx�:p�~T:a�A�UB�IL�tr�$��9���у��zIZPd����	��+�wt#"beX�5�lh���1��ޚlo�HD�Y$m֬	�p�-O��P�Jg-�J�h��
!2ơ�,�
��Q;�h���Ձ|��7��՗��^��nߑ��^�g���� �*�aE)�*l��(�:�^v3�V}z~����C	t*����i�����IƝkW��ut߸֤Q�[i�/�K����/FCVf��lH�N2Ku�uMP=��&ג�ͪ\�s
y�����'ّ����@���޳��#���B������ŽnB\�B�wX|mF�d��<�������#fO���y��i}u�F)������CY��哏?��{_�'!2e���+*6�Q�ؐ��z+�uU�ZmY5�������$ФF���3�����yG0��I����ڨ�t���o��Ǻ��LT@�A��b>�ݝ�&�=���^�~T#�c��D���� d#^��x����З���Q�[��X��VÝY�R�M
M��H��2�N��؜�ڙҏ|�>c���|Ɋs7���f����/l�;L�3|���_��&A
���||牁
I
W�`v��cV��K;Mݠ[(uG�?1Z�Ld��zi%`�&���bM9:�˟~���ci�-�h�[o���Ҁ)�m�¶�R÷�F�P�41$lQu��7����ߩ�:�A��RXI���p䨐j�U�E���^�U�~���l�-�p�����)y�����\��b�b�҆��� �F����	9ː�hG� i�+%v���L˚�ޣ���\QS�����ipV�=%�N6���J1�*�����w-���{�T.�ޖ;kz.�	-��䥱l�eJ��
����N1��� �J��M$#�&Y��e*뢈Hg�VY��l�ITW���oY2��X�(/� ��z���Y��>er���@
��0����A�x �쯻�~��\JQ�U"ș���ׁ/�SȱxU �6�z1���s{��r2-	V�f�)�4��2��7�uK.��5�h���� h<�X��]���o�ɤ������֭�,���tp�Ae��B�8#�q��s��1gg�ᝤ��m_x���L�$P i��R�VXy±H ޅ�9V6����5�3�M�ن�dTm��/ zHN��Zp茡��1�	�.�I�1"<M�V3B����JJ�`41)�P��砍@Q.������*Y1��
ĵ8��`vF!@��޺E��������xT@���ܽu]v�����Y� K��J�tX'��Q��S)	Jv�j��a�^��+�"�zK��bC�<C2�ZL��Ol&h0����4I��}�k�wݛ�V7�z[���2ɏb��~���*�.���?����ݖ���v8�	��m{�3\%��A��]�	G���"oЇ�#�d2��1��P������\��/���u]G�~\���!E�ډ��k�0ј��U&Ah��0���h��X�����Ͽ��9�BLQ��-�CK�H<.�|T5C0C2���A񸞐&�q�֐Ť�i�*S��5��������-�PV['V�{�XV��\�zk^�A�f�!�U8	��넿t����8���U�^?DE'^��y��g�#��x���`2�f�C:3)�LL�F`�R��uih5���NGºS���,�W�":a I��3M�^��h��J*�N�h�,2��O�R~��gW��m�x돡[@l���4M/ͮ\h��#���|(���iЪA�6Ӟ�(���q�Ph��sh5(+��%�Q]��^׆"�~\��Rf9�����W�\>x0c ���R[���ը��&i�bd�W�5���^è7D�`� �+�NSR���L>��#��4�B011f�7�wu98��c.e��D���_��cٽ���L��X�
yxMg��bk�֘�s�W�@I���Q�F�|x4er���2�@�\K�9�N5u�y�"_�X/�$�ɮ�%��I�Y��f��J�����L� ]�ڒf��y��,U��9��A��� ��p���Wџ�U+I�M�41d��4��|i��ŔC�h�^�L��&~�i �?:�O��L���5軺}����?�10�@��ֵ+��4�D$�)�A�=v�>����@)���J��=����M��Z�g�\��H�6��W�{�oT��FY�6��-�w��A�wi�~�
[g�A6ß8m	���P�Z\�D�=�ৠV|ɍ�@�Y�.����K��?8�����xnj��U����^1�(P�;|ߜ�:���s`"��l�1���i��y��G��F�� ���?9��gk�7v�ן��1�3��_b!��6`��&�,R�
$��G�.�pZ��j��4���)� �@��?�v�zUi2��<��!�h$���2g`�>�#�E�
n�U�5�����ȣר�~�|a����'��)*����^@p�����LبW�Дw���
��EY9ӒIz�oH�7;L�:�#(ڃ��V����� �c�D,	�+�nP��<9�ō5J�'������0{d�2�F64����P�O�e�	-#G����Y�EտY����̫	�S��	�,��+7X��q03�4hcP�A�*��i�:�v���H�	P�{׎Tю�c���&fe�k(ռG�Ea g��N�'��&�����@�U�K3�'u��������qVa2��
ך]�a$��IG) ��b(�@���x:����7[}ȅ,��9�����Pz6fKSlD��9�0:A%bA�f���{�"+)|�i��l���ͨ�Yq�<��wo�	{������癐`fq�%��ggzTZ�1��s�YͿ�W
����R�M0�!�
>���Yn���j�a��lf	i����(��~����@�
I^� ��*�zN� ��O������v��l ?>ݗwnɭ�}�8��{�~Y�f�#3d	�)�6п��������@��̃/�"Ih2��s���+X�B"�ibIE�U"w�Ql̀U�����x��8�>6��W�Y�'�ySA��n�X}�`ȼ0�- X�'�����b��XM`6�L�'�f���n��0�-Ն�5��{76��ޕ������D�

�]���l�,.Ne���X�ǟ���?�I&f���-P�OkU��#��AA���R�v&��w�?��dVc�wfB[��.�R�+ξ���6��Rt���u��	��j1_�"~���Cro�������s�HoGbb�J.�b��;/��(��r�f%)��^�z��Q�z�Y�eH&Q�Y��K{��Cy��i�r>��fٔWJ�Z`Tx&��U@zχc���(VNm"v��ĳˡ�\(��l�y ��B��w}����P��ଗ<0t��%c�l`ɠ�U�d0r峅^c^�k�Rkue�Օ�2J�ؑ�'�Dܼ���du�,�
=)����R�׳���f��\�D�9�"�gcV7߾}G�F�4#P��܂+��f���v�+F@��n���IU	0P��wVy���Pr�t<�B��ښ��]�������U���|!�:����C�h���ݻ��[������?��A8o��(n,̸�Db9�1X�YvY
K!A�:]VaA�B�K��6��?�NO]�*�.md�W�SDyq.�r� %��S���_�@��� cb��Ӏ$�\�3 z�!�R�pD	�=x1 n�"Xc.���WN�S`�o�9?[�a*֣��2X�Ѭ��&0��B@�������
�f������Κ>/��&���GHI�xl�hs�5�'�y{+��
�Jx��j�ͱa8iP@-��ps��do(L��%ED�+������)���T{��x��t{���A�a/����g3���G2�!Hi�$D��� �|V�"�	�Q��kaT)���	X+��^�� T(8��38�;fŊD^�4��MQf��*{jb:��&���]\��\�)������Xڰ{)�=K�h�\E6V�O�Bߍʧ V�I�-����X�����2���w�����Q�4T�Gqdt���ܔD=�0�����A��*��S:$�љ#���e��75Ks�ռI���w���X�e:g���n[cU��x5/7YV��i���P��ʣ���Y	1���M�̞=��$7��^�t栭�NA((3@�8�VKZ͐t6R���,rf^z�Z�X���d�$Pl����g�a�U�9�ש�ތ�*Vܭ��O
���������QF����9�Sq�j��`+�-Ѕ�P���Zb�'�F��.��y�b�"t����.��G;�y�U�/D��C�X�⌬χt@�Չ=#�?V�3�먺k��t��k�@�}��<~��j��?Ę"��ov>��٫��7��/X���5�%(������U���BU�0
�E��h�D���1�}��l�`0�\P$7�>�"HE@�v��rS����B[�~��B�f�*��T!s�EC����݇�B҇wa�XT���b�SP}� h���,%�5�=hw`'-H/��90�VF�3�N��5��1�=��-��ƌ�@Wk�Xku���u�w��|���D�F��I*|.7�]�}z[:��g�g�*˹��7 ���GX�m�����K��`��Y2v@DP��7��d�4?Xu�@��Zz�Y�{ĵJ]Ӏ���F�+���T-VU�����拸?$�	�!. �UX%��l�9@�k�(�N�w��������յ��Z��f�d%ۿh��Пq]��;���������G�ۧ��J�Cy�O��/�������1�M]�������n�#��A�8�G
<V�b�*V�
�BJ�'�<����>�1f���"5���17g����h�?>��㪪�U,���+b����2V�WV�U�(埊񞄋W�Y���,�=!�U�+RA��8h`��5�?�K��zW#���4���T��|�JLAÆ�9�15���RK��|j�T�굎����щL�ޒ>FO`�1N*F s �K9>���� ���� v��fH�`\)
a%i�<Q��A(^4��x����@���[V�+~�;�R�D^q��.�i��3:����e�sf�J�^��s�u��3B����⦮Q�+D3:�^Ъ�8ծb\�.�B~vY^}�/bx��:P���9 Gc� Ā�\d\�b�i�d��rSRd�QS��#�������OO���z��|��[���o|2�ӳ9���g�Au�.R��r����#Z^�pel��l��8���K�pe�r��+�V�y#��q~�� q��G�\�]R�$��:}�3&�Uz�tT��R�^���V`�&�m�t܋�����@��>�t\HZ�3M�5����6�#p���c\����<y���'�.M=Υ�i����Y_��`8�hYrN�|�����|q���F?�� @뿠�n�GAYEs�xj:��Ta�ti�SDW&���?E�Y���`�%UokE2�:��
͆�F��2����{ ���q90���T�@�6/��1P�Y11*����%�A9��Hw�"����p?�P�vgIÊ������Z2�D		�C�,��>{�����P.c�.�3'���)����XuG]��,��֟��[�k�4 *�*L ֟mU���DF��2�z0ަP۔�HI�4�j�3h�]>>;c�Z�xd�ѿ�Y��(���y��K�"Ƴ�V`��a���3f�iK�Б�ª��^�Aʙ��z���3}�4�>v��T!ƺP`łۼ4t�������n�T�򈉍T�t���9(������>`�~_CA�����%�2d �r��82����� ��Ϣ�	n�I%�?#�)st���,Z%��˩�`䔡]$��>��E��1b�PsÂ������R*f����@�w8� <��/g���t��(�s��3U��
L���~����$��
4��\�}q�5T7�ƲX�/�3�\>���>k�( f>�	,�ǀ����f �5"�qkW��@N./5�X��b"�|&[k�z��r���y�I���|�gm-M�4ӳ8�\r��)b�+��m�W� >�9(��˸&2�ղ)���yn��7?��9�K}�I<F^���;8lc���UA_PU�a�xF���M"��p5.+S��+�*�k�$�\�w}K�y���4�nOn��ߖ���"(}׭�`�.���:����l��ge�U�pEIó����gM�ץ�v9X7I� :<:����˵�]ݷ�l Y ~���j�P?E<�~A Y��H����V#��]��<�<����!^aO�3%�s�(��d��;&���v�¿G^Q"�bGc�rUI�D�M5��i���j��S��=���hV��%�b��
T�Kk� S@��ƈ'���ƃ�<���U��v
{�_6�$P)��;7�dx1��:���8RYN3���h)���&��(�ޗN��8�*T}��\YՋ��z<^%�{H���+�W��Ӭm_[G��5r1aW ��[�1S�ߠ�V}�	4��^�0(��&A���_~��f�1�Ǘ�֜�K�]i��{+fD���J��+���-��B�~T�r�U+(�J�l���(�T�
@
�Eؔz;b%�G�,1�����!����)�륛ӑ�o�ȗ�<�߼�l���)/����l9��p���5�8�3`��u[����,-,"TlP�M@���І�ۙ��!�(����UA�F2�c
\ѫ*E[�kF6��=�B�$��}L�J��Z�Q��}.AG�UH(7���c�En���F1���Q^V�\��f U�_u�*t��+<�7�†�]7��x��T�
�t1r��sP6�d��?�G����'���t(�ۛ����ʕ�M&��Ġ�E�U��2D�<T�N�TM�����=e�|�:�Z(c?Tk�!+�����|9V~�D�JY]"'Ga��y���D��#�2.���x�U���B#[�DD�(ZB*�!Jƕ�7\~�(�=����y�%r��U��p����JO��aX���I�O	{��*訖�h�S�'���ɓ==�m:4�mC)r2���)K��5�hc�C�\y1��r٘�ā�K*���E"�o�h
<Wa="T��K�9�z��"�R�$"�i�^C�!RR;��Q�Y&��k����4�G&�þd�w��3��&���r�1#���� ��?��'����>�Շ���K�g���XB<TF狹��&�BH`b���u�/<~��8�%�?COgV�n�r6��l�d�i�ti}�p �VO��uV6۝M�����h�|��6o���m��0�h���� zK�lч5(��^8?�����/���w�����������d��i��IDV!]f�;����~�96볳yg���99��+61_�*�ǡTv[�~��C�k�C5��h����]��H���f��tl�t"���!�A"�ł��{��T�z��'��gN����y�U#��g���P��3&�)���T�1h{�g@���5΍*�����y��+x�~�c|N+��*a�o)���ي�c�0���Ab�2�_3R*}�D���#��{ Fza!.J`};��y@Z.|P|*o;pc=��B|~
��ef@�˽��&9�n�EAP��u	���Ԭ����X�S!Bq�����%�����[�K��xc��j�/�2S��k2��qx,��t$��D���8=����\�� 5�С�i�H��<�����gʲR��Bd���1�4����x<���9LfT[o7[r�����@�ٜs�����H0*�s!����US�wZQ,���%Zw�V�@T��«�N$�#��L�w=r�� D��/�dMԷ��&�Wv8?�V�Yu4��/�ߙ ���\�7MXA&�~P��"X�=,*{%�����0J�3����4���A 0#.N��P/��U��V65v�9&!"H�u�Ϛ�}�#�j(D��YX]��⫈>+���G��<i|R��2��>߽�LC��x>��h�Y���/\��
�F2���%��#�?�ap��^�} ����"���-$�Z�E�>#�|�	 UiD�F�	�t��қm: s�E���)�g���+B���ِ����	��`Q �����s.��o�HmS�zk������	W�/�5�X�a�ga6U�jS�}��̭ד	~dnyŏ)l�F]�#CD2�Kb~$kzWC��]�K*+�7ν(��#�⬠ [�b��X7;W p�"�uк�����l�#0c�	�˴6dU 
*�S�De�j���N�Q���
W����,R�)�#�k���5��n���3���̇�{��A��&�?���{�u9z�H��Ϳ�ݓ�e�x?4�>.���eM�:z@���D�0 U��nM�Bo�.s�^�<�`;p����̴K*���&�$�m��ܖ����O���3j2�4��$��(+�B�@��|G��3C�L�bF����C$I(Ԫ�!bPF~=#ј�x�C�ї@�F6_�e-WR��_��qV��:(DZ�`T+�9Pm�AULl{�+��ͷ�?���},���i����>�w5,�X��&����.�XPn�b�p�f�"�'��VF
��0G
K��`p�8��bE�QL*)�2�S��1q&)�_�����z�*��Q��R�g��Ռ��U>8 �0�+������d��#�,s�,]n1l�(X\0�APH���/�i�U�R��/�1��ZA����#耠�bO�<'l O|�Lp��fS�/���9����%gխ]�!��s���J�^��1��;���8	�E���$�y�wU�Ň#�EV)#v\�_�]e)y�Xc��HZ`�%I-����,�t�U��M�S��F��{���0�=�6X����T�!7��CC[�0<(�.���躴!���㮫S���K꤁5��X��Qw,@s������7�#N�,k"�ϖ�\�A�n����L�8����2�w�s�-]su��>&#Q�������ٱ|���}��8C��`}�	��si�'<�3m��N�I��l�ĻV� ���'���� E�Xz��RO�w�sqcg]���<y�T�_=ӵ3%������7��Z��yX��
p,���GU6�NP�`g :%�Q0�]�9�84���7�q*��(J(kk����(������ppa�T����+���������'��!�w����*̾���يL�3��<�`���F�ɳ� 4�ٽ�v���-�h�>>�ԯ���Iٯ���.����m�NW�N	���B>���!��g��d�д ���ϊY�3q<lfܰ~�2�����2Y�(C�K�R�J������T�8���H����ʷ�	4j�e��j���H`K�����&����� �P��1��$1���4$d%�V�m�X��i�W�G9����t쀞6�yF�j�j���f�(m�]�}*���9u%��lL�=��B��� �*0��L�*k�:ѳ�X�ȵ�]9-�ƍ[rx:��L��rN�:џ�`�o]z�۬\�_���@:ݮ��,Pӣ �c@�.lD��3���vӞ�l^1��b�* �Ϗ/)���&W67$��?��?���>)��w\���կ-�~�m H>0�	*� ��F�٪�z��g��I*�Š��BQ�(�qBdS��c���1� 㦾��Ky���d�{�bD�����+�O��.<y`B5p��ނ�	�����I�US��0Q�z|�Y���C8��Ik*�XՆ�▁�k����y��ڲ�T{̂����@����>������������*s���c\��u�ʦ�>�>�$��S� `E�ͮ����d8T��&�=���7�u����R��y1�x�L�Y����\LuV�%���`]�'bdXG$v1U�g�i�Ծ4��FB��'M��,�����J轷l疬Xg/��>/�j��
la|�v���s�S�	��m C$kqtͺ&������cNqf雞Tyux)���dm{[�1��t�sP�� dp�mQQ.��Y�x^�߈�Zg�PX�=�n�PEB�̘O�g�1����"Q8#h���ﷷץ���ZH�	�>2`O~������p�Qa0GU$��GAX���ۼ�$��t��O32a N�?H�7�7� -���8�=t0��	�XX����zW�Z�DL��M�񳸙�u�j�$�i����تȼL�?C�71���e���%L���u�}�T�o��'���3��N���#uxzA����4ֱg����Hs$İ$S���+sh�QE�˓�eS(	����*Mq�J��\���E  9ܨ��*�*Ԝz
9�eFg��{Z�!��&_�;^E$[Y�=���\}�YNQ��JCea(���#^��Q�X^v�Jx��u� �6�:�������7�ܨ�� �n��x)?<;��;�䭻��ߥ���"3�%C�\+e[�T��C�w�e54c�eiu=H�+����V�؃�u�zN35�c�U���E	�̀'�S9��+v&s�fskt/JḨ6OR�Y�t���"�-���Yt>�d�0T�� F<���
����I=/02KR�@A���sV\�萒��=6��ey�O���07�5�a��7�#1L���F��
���<��git͹��ǻ�+��=99?�3 E-և�z����a��:��*L���bV�;��[��(��h	�m*��v�^<}�X���(ό�(�����m�uK�M�V��A�I��xW�h`��1�+6��O5�������8ט�|8�F<�t�j8"XcŃ���kƍ��<:���(��������+H�?'"�Л��U5� )[� 5Ax5*����Q���	Q��`�P�$���T�z;�୛��6���g|o��������A�I5 'ؼz`�d(H3����8��
��(M�v`m}[6����j����dx�������XC)�]6�-ƺB��h>�^cP� ��N���S�ۢPT��Wz.ML&j����	3&��]���E]�F�wjJ�@�Mh��!��]�+��Y }�3Jb���1+@XQٗ���b��fI�X�~�\��.�<�N�k]�Ao4c}���+b-��M&S�����=�������fj�H``_"VF7F�Z�&8��R.O�2��Sz���P E#�VYh%�T:u�X���C��eQL��Z3��/��ֲ*�ʇڣN[��d����J��UdTAzk-�S>.X%1 -�s �D/#�m�?��ba�x�^��(�3sDP��=H1{X���vԚ�s1�x;L�xj,�b4���\a8��h�S�L��g�\�j�.(���2V&r�ibB�ۉ��X�3�*��S h`��w
�1}o���������޹"[���09E�"*+���	� �z������4!(רe �p�g�>��TKf<��ՙĠ��i�9�`��׋��)pE��n�'�L���L����PБ�"I�~-M�����\��*䰯�2��C�7lN1n��Å��=w�l�w���?{�棽��{�v���0M$�H|�a�x�NG7F�-4&�i���s��?*y��b�����8G~e��`� ��Y6���p,��&��9{��l���sk'�������`y������1ī^�5�Z=ѵ�S9VSP	��J[���ˣ����|�y�1�l����_��q���P .���ļ,)Dr� ��y"��L��Ϙ����,R󏱩Wg���ܞM����g
`� ��{7���엄��z���D��X34eL�������/�>e*��F���$���Kē����q`�Sإ���d�0G�V �8�	��aSmd�։Ef,�5d��e��
�U��N�Rk$��BҦ�\��Ča2W��`Z�9@���g'�ۿ���Y�;0�@�{M~��O��ݫj7B�%���U&���*,��P�d��J[ed>K����c��Ky�����b(��H�ώ���B�[k�q�,�2ƞ`��"��[KR�}����ѣ�}�K�#ϥ+&X�K ��] vD�
#\4���K�Ҽ���h��gg ��1j`�,A�A�C7m<���t<�o?�VoM�{�����8��O4�ސ�U�1�A ��&qkp=��f���=��Q�ȭ9�$y�N�QA�**�+Z�OU��T��Xf�CԨ�r��H�2H�
 �'�����N�A8!TKо��`ö�s��w~���K=��p� Pi|��x.�M[���w��$�� ѐN�F͊.����`f��)E6�
)�+�;{n"�<�Q�e���>?ʅ��<n�sv[5����s�ļ��T��Tһ|�j ����]�~#$FH��[�o}j&��y��0f��>`h���#C��U�f�!�x7&X�I8��9����i����_ 
�GR��&����kF�,�_6hp��~$c�_���9��0J��}�9��;FqN��5W�Av1�j>�,� �碒N�M1$�SR�P�A���gg>R�i�ۓ�O�h4�k�x��)����C�B���=i�c�p��@���*���䤂�N�d�zQ�8.@1$����x\Y��/䇯�dU������ki�o蘣b�*��n��Lzg�9;��s���Mht3�yP��z& *C ��u6�g;V����-�?�N���O5a��O�w�)����L6���p�IO(R�=cø�^Dݦ���9Qf
�!)'�c
 v>��9��K6�V����*m�J@����(1.C��2��z�fL����r ��D����&�艴;��A 2џy|x ��\��G�^�tx���R�x<V;ېV�'���5@ܺ�-�7we��&ihӥUryWr|��z8���gE�:Q���E����9b=��j{0�z�I���rqv�~�&ᤩ�F�i�Ր��-����ޓV���{YY���Q���U[T44��1E��,�$� U������8g���\M�2�	����LgV�j �.�/�_kk@ޗ������]���Y0 b!AMF��P���C�Ԯ�5���"�M¹e�Rm�ԆQ/��'�@�<�N���>G�Da��"�(�_ܰ*t`����*N�
1>�� ��1�4����/���O��g6��ڢB����O>f��2����|��
t���m�bEeB0Nzf`TB����q�z�pU^#��A�c�Y��,��_}K��O5ɹ�8�[�n��kW � 1G&�b�ݒ��KQ�A�>�	9T�Ѣv�7!nz!���s$3V��3���ۜ�'4`���?�N��U��
}F/�}�"E����j��i�^%jo�z�0���N�J_̙��<%������	mhO�XS?��6@ ~��ic*�^��v���KB;V��9���"��Mds�*����ɥڤ�,4�j�bnm�=�����aG(�0�°�Q��o��H���Tj<'���s���	E�z��X�T;���9��c98<��>G��R�o7z�������"X�T�)M�,\2� �`TȒq�z�Y�z���9c'���{�R���u0�� �J�2~��/Y�S��7�a�hcʬ�� .��F�*nT����/ �!q}�	ū��b�ݐ���<x�m��|KfeƳ �X��1na�.�k���X�XPPo��0��#P���� g�&:��j��z?�Q~�w���>��<������\n޸K�I����u�J��2��<�F��� ��:��ck��b����ٹ5�3�N�PS�L҈1=a����Z��[����X4tͬ�6�n���B�	�҇3P.�*pf	u7\��P�Ø��8� t3PL?�F�̧y��s9x�G�L���;��Iad��q�3��[�po��y�]����Ƞ@�u�X�� 2E�<�hy����\>��g2��H:5Y���s��h��dĻ�ʆ�
L@e��.+P`��Mc����]��&�����bF�G�` f��5pq8W�]1����&�޸�.�q�/�ec��^����}��.|$��\��E ��(Z �AY�A�7E�ϭ����eO${1��1��G/	�z^��D�$T��TBKx�@T�{�i�
Ҙ��u�ïCI��� �:�T��!��t::�%�&���^��h��x�d ��N�Ug��˲2��\�"�̸��#i�����Rs��F��`[�	� ���2��3&�U[��D��*&�8("���:QFMť`A� ���Y����ÓK9C��L%+�Q*c�(K�s�|�$K�[��6�y匍���I$�!h�)Q^�=��Pc��)�0ƜV���qS(�͎I�DO(�6�MSN:�����N�tMe�K���~��o#?����'K�B���F��#�&���J�(��<Ԥ�`�����-��T�{�+�n[F���M}(.S��@եz�6�-W7e�'FϪT��q�R�9u�� A�#$E+'�#�щ��Lj��Cb�5Wcqzt,?~�Hj������j� F���]��a$A�E����)$sP��Q^֪G���u��yaxj����3��4U�@��NNE���\�����+*��?f�
	��(�&�J�ѮɊ�`�~0��
�t,m� +�zq��K?�ԩ����mi��#��T��?���Tv&���t p��mR9�Z�	c�K��i�E[�{]��@D@:U]�N��k�u�{�����4˽7�d0�mR�A���<A%�x:��h0`��ֽC5u���D�[�9�(I�	Ή��w:�)��/����,5),!f�A%��.����Dd�͞\�qS���ޑ��ڛf��#8��3���V.ǺG-: V>�Щ���5ȜL�
�jJ�	���Sy��Gy��w��5��$d%jʡ��f�^��mM�]�mML�Ϳ�7rm窼�D��/��_���6�����1Zef� �@��)�U&u��k\'�&��d��O������3M@��5SV)� 6.Ț&�kk�r��m�u��\�yG�iW:��>�ĪN�"V�pv[��-��x.�qj�+5�6��š�����L�݂>�O��EU
�ͬ�����X7�'��$i�#}�0N�y_ǩU��:�;�'Ky���D�g�i�����mB�/�� \ւ��SnBK8wLl#��u[6�	�ya=[ ��Nu_���`��,�Q:X��~�Dm��~��1Ȅ
,�����Zv�\���z�[]T�k�����>#x�Z��P�FP��w�HפY���4)�[bs��O�hy�M����MR����W��iP�#0�������%���H!�p�x �p=2��`���LƮ��(F/��59XW[t��M�ڹƤ����$�P*��&@V� ��3����W�`c�����B����	���~�=�x�@-P%�s����z7���P۵I{��젮	K���Pm&(�qR���l2�Y���i�m��`4���F�)�~���{O�����@����l'��MMl׺[����!�[;r��mٽy]����n��&����(l.�q �H�7,_�v5K ��H@u��`iq�N�6�����#�.�l.(�Qj559m�5�����E�P^[ߠ�w��f�9�Z<���`P/�[bN튨V�!�-�Z�@-G|cCmD��j6�8�*������l����{�{S�X��\�~�9�m�l�f�Τx�Ձ\����X��Ҁ]���7�b�Ő����o��M�~��9��Ca:�8��Fwt��٪B���*��[�.X��8�9ћ�uZ�Q�f�]���Sc�}P�L�l���h+�_���^j��DsntV�5pn���&���˰����"�D⋼��\#��&g�Lo���*�]٠-���m���,�q�̥��cT�'3���]F����f���t��A����TbL�Z@�|sEћ{z����1�N�yf��b[�nd[w�� ���������A ��`4��5	$f�o�������&����Υy �DƢ
���%,�2,����+0P����(s;pv>��4MN����������T��Ķ��ŤЅzX�F�`�w�l���Qá�MD�U�������M3S�#�	�V5�)�E�h���Bx�\�5o��@5P�����L�Z��3�fr�K�2ޠ�ύ���f,3���H'kPWk��� �@O�%�� &��h���W_p�4���|"�������V�*>�u��*A@IV7��0�a�!�5�E�W�fjֈ=�9
��Wg��Xg�)�!rC�/�@O��\�3FB�Fw$�@���u���������Z�֖�O��쩫����u��OM� 9���Q@�";p�^��Ӈ%EO@`��7<��?��s,SΛ��N����Yt��E���UZl)wp,���}�-G8֓�և�3#r1��g�BFG��Խ��lh �mm���+����?�04 ��	0��UR��"� �W�c��{\K럍#o<Om��� Q�L�e�Ay�)й��Qy EI6��Bb�6O����b�LPZ]�~t1���@�jL&@���}I&��C8���Q��M5p=��6�F[�H�&ݨ�w��1^&�{�Ψ�Ρ�l�`63�?��d�ܡ���Hz�5��M�1��I#ЦP�먡�]ov8�I-�O��a�CAu� �w���`���顟JףSo(B���#�E6[aYa_d�#M��ٻ6����p6u�ir���j�U���9o.eu��B�H�yu��ݐנ�# C��� J��WG�"����yɷW�	|��;=9���=�P5�����Ԗ�5�� a1�[
��Ź�7|uS�����M.u�r��}ٺj`�I/�5���W$%5���`q@�0��>����W���O��ُ�ɉ���{jw��� �pS@~X!��@�u9�ߖ#P������濔������O{2��H��i�$@�U;�q�q�ABa4J��~�����<����������O2=�g��`"+�oT]&��K����s9|�<x�#��W�R�]��g��S5�����+� J�S�E��H�Uk ����������^��W[�{،�l��AU���s���d�]8e�~�#��ui��Y%�Tg^��٣5Գ�JaR�e�t��=҆	���lb.[LeC�{��&"Fe`�S�?��Ʉ"ǂ&�oV��V�n}�A.���lAP�I���
��F {�=�������Kz��Ф�)�!�/X���
%�	z���Gc�|�P �ni���i��%j�uB�� �B�#�j7�n`H}D�d����cl[��v���ޡ���}1b\��HF�$K������>��?���S�{��d��j�.�Dm�[�uuW����G�AB�?��d	�� k0��^h0��q$�a�V���w����p4�G������'Mp^jR~)�&�e:f"�79ӽ~���X�l_�-Wnܑ�[w���IBU^�H��C �mHuh#� ң�@��>�77����Z//���?�/���O����Z��c�)�=WQ�R۩��wEN59x{�����\L�5��eL1Tf`�q�Q7��0�H��Y��7����g��ϭ�x0�~+?|�g9=z!���t퇬����*o[�e��^���������rU����5Q��	7����ѵ��8�f�bBkIl3�� �@OZ�6E���x�Dm��|%G�{����+u�vOק���';ׯ����lc�(˦�
-g�6��
j#�f0� dGX#��kkB{� �h8���9=��`O�&���Q���\k��ƶ\����u�c��o������� �"[�y���+�enչ� ������g�W%Y��~Vh	?�,zf�( `�М���H^<{)g����h�f"n1}h S�����ܼ���R��x����,�������$`�cBYc㈊�������O�<��S���;��rD��1`[����Ɗ ?w���mqf3+��#:�SG�1�;fL�pmA�n7�>�qm�~�
m]��^���=y���z�k1�j=U^�]z�t���ҳ��uE�����]�u}��ǌ�?9�Ū�-C��Zo�n�:'֗6|��:� ��wl@���^�/��T��8 ������c��s[��-�$�Y^�e����ʀp��)�P�5	4����!MT !w
�o���{�q(�s������+)��tcy��L�Nh,��o�KM�c&��l}`�G�� pG���0��Ɵk�'׮^��+;r��{=�/9����D����r3IA���ށ:��� %Ҙ���ܿ�M�$8�،���2S:�%f�r�諡�7�D����7�f1!��3������|�9i~�nh<փ�j�T�%Q%A�B5�9�+�L���+���X�e\䂴E��h���e�䆓)�j!��@��yЭ��Xpf�4Ȝ����3(E��[�G#�d3b�mj�����_Z��^it�0#�m��Д���(�3��S��PIW5C��v��O��N�Hc'�Mu���u�Y@auP<�zf5X�iP8����X2���D,Pi�f�D�?5H�͚&��W���h�T�^��,-
ISD���T����A��bI##�lu(�4��Rk�FpZM*�-��L�k�N�����������4��r$��Rę���w5	��ٕ+�o�q�#��i��L4��Һ�\��,���DcW4�����jfJ"yC�gq:�lt)���Єg48��>�w��	C�� ��6dcC|oS��{������&I�~+PAbW(��Ԓ���͠��.���4*zL1�L�A��م����@�T���8��� � ��7��A�����{o�֕�z�*f@�Eج�@F���P�w�k��6�g� BS��C���	���gv>����d��r��̎��Y���t}[�K-��5�@R���ف<Sg?�<���@���H��_�`�m=���eQҜ�2��z	([����f�|!�|�<��K9��Xj@!qNz:jw:4j��@Ϗ&��g3�S?�R���꿖�޹�)ϟ����P�UY��;�ViU$Q��}up�{�'��������A�{���-��H�侢� P�u#bВk7�d|��N�y��;|5p�Yݟ�+�Yv�_�Y�}0�;]�' *���zP�4	ԉ/+��r�3�%�*5�>�9�5�<?#@�����kp6"�w�ZG�d[�+ׯ�=�o=xGDnp�um���@_��	�V쵞�t|��O<L���^�F�)��F�t϶�7�^�# |!G�،.�nM |��V�t��ܼsWvo�9G"�����Z�v*w�- �ъy�P�"�+���]���<N$����22������'~??���DK�-طN�/�vo���U�P���Y�:�S���=E�hNyy��rq�YEw����pj:��V�ƞ���nD�H(v�~�k��?�$��Y�e��]��7�c98���~R�q���>kk[�5��ѡ���_��������{�=�g��B� E�X�KW��X'(8��g�J��������@���s���iB������}�'A5�B��L޺}K6�V��+Mr��TN�N�P��s���ɀ~��X ��Lr�������J�L
	)�����?�^>���9�Q��{�R����~ԥU� DJВ��B�S��z�̸����V��"X=^�ɶ��Y!F�E�� #X'�	r�p���VZ��HJ����>ߧ�O���~�H�4
f圝�{ *�znr�I{{}�1�J�sޕ���%k�zw���S��o?C��^�f[�8�� +������5M���<��+y�ݷ���Ϋߝ�}�P:�
�M}��Ֆ�޻�����������.�W�X��lIPw�4%�[R�1�FTq�0��TLȦь4����~|$�}�|�D�#2�c�����_IK}ݦ�Vh܀'�����фP���%�O#�OB�\q��Tc1 8���t�� ���ʍE�>�҄�j������F16�=Z(�>~._��<��1[4 "��~���o�v��xu���M�Ե�u����I�`����x,	P/m��1?`��ߋ2����KX����˧��/��=T{p���@�ߛ��M��ۺ.[�]�*�G�3]��ֆ�D�_=���t#Q���ބ膱s�`c=�n�H<��6���x���?����ɏ?ʾڔ��G@�&�]�|�Ά������/����Ձڧ��2ߺ���,����-h�x���f���iO��Ĝ�Djz����.����㋐t�Z���u-��Ѡc2AC�(u�m���	H�T�	V���?�k�u�6U��&C3��[��޼{Wnl��Y�I�@�>3h/-͸�'�>@$��2�� �Fv���U��%Ss�z��ݶl�*R+3��{r���v�v�k��Mn�իk���ֵ-YW����r(���ɞ���9a6U���ɬO��9.˽/�,����nD89��L8��1JٹUE�(A����V�UG�#Q"4˲y�4�8�5��h������k3n��Y�`�����EF�d"�"��6�A|h)�Y}6�$�ѧ�S���5����aCzzAgiC�f3��SI�,7�^�ȉ��IG)D*�
A�U%4ڣ��>:($r�6x�zv ��H���� �ʦ&�%��KR�Lp'�v[���� �!#���V�R_�@�Fd�y�7�v�4�F��\%�;qV@� �4�s4��D�H��?�9T����L��P/�QV+[�X����>�[���ؐ��=�L����VǨ�&N�~����JK��1�yM��r��0�����d#�P����s9x�@�����ԠU��\$�z�l5��X�4���lO����0���[���~���'8�I�����P�L�k��zT�З�QÛ40�&`�2�(��8~���P�j28SGU�/0��s65&r�6���T��&�o��{�~$��6z��E�ʤ�-��V�#,2���W#��ѕ ��J�s�/�O���\ɫ���t�	}��2��ZL��.4���u�O:���[y��]]�_k`�3uޛzw�2O�5Ω�Jz򠐬?A1U��0�0���5MV��/���/����Ͽ�NNt���҆�d��	��v{
�0�B.5�8�szS"�	��B���,����5��k|�J�J-��
K�Q���F�~Ԥ��l��C���/�៿�s=?�Ã2kE��h����p�0��P��`�k�5�K���:�KM����s{�w|6M��bL�&�|�8�U8�΀'<__��\��?����O���ZM6�-��K���}�s=��>]��H��ټd`�ޑk[�2��{Oʧ������H{sK&Pd�8�������D!�N�������\��V[�\:�rG2Bх:{sP�@R�d������{.�m�gz�Ƭ��P��Ƈ��5��[;r��B�=�}��U�76����DP�6���7��s�s+}��-�ߛ2�����.�Й�����gO��gOj��\RЖ5Lj����+�������Y�s @�Nރ����I�����y1�;�D4��m$�=�@Z���y�77(QΧO����פiON^�"�7]LH���kXC�f�/������ޗ�޹G �ǧ�9cu��%����>yi��`��=��J3����&�G�%ihP���y��;�?���E�������;��_~ I��=<�/����8�����g�����:|��U���}�srF�u��}V� ~`�a6j6a:G�z)�v[}ƾ����[��ϟ�Mޗ$p�_c���{������/�ݺ'�^�7�=��/Od��@�Vm�����g2�����~.mM>��f-���iPb���32`t�>����rzz(���?���	��5��i �R{p��u��r&^�Ő ���.Ǻ�KM���0�S�,4!��IX�61cܢ��V�� !Ȏ��Oan*� ��<�
)g�B� .4;�O5a��o�?�P�/��ޙ��&�z1n�b<�4~���ń��`Pd�Wq�!0rz1��ֽ�\۽�vA�Vh���з���&Cz~C�wk�cN�ї����oe����6�fw��QcR����ou5i���(y,MT��ߖۋB�^����@ ̫o)��oF�>�o��,Y=O����2�\������5|L�)��%7���j�і��2���������m�j����u(wߺ�k�͸rI1�G6$�������Z�2^�����+0:��.۷�C�`1	�{PE���վ|��/���>U�L��)E�x��Dw�-�㗮Y]}թ��O^����r�����l��	S����R޹��%꽟�̎+��w�^y�PU�h�gS4")3%�&ڈ�agwbwb���iwv6�Ȅ4#���Htj��4<�{_���vO��@2����B���{o�9y3�1��ra ���!iV�e�D�O����g�c��C���[M;DD4Pr�t6˂k}�=����<g�0>��`|z�\�A�&�լާ�MG���^Hb�1mRA@�+�w����/�~��ϸ&i��
ϼ\�Ե� *F��a�dL5���%^e���:�Y.�c&�n���^Y_t�#�|K�����S��;Ak�f��'�ՐxW�f�;Gf�X˕t�A,��5'Y�0���dI�lV�ƶ2j�x��%m��t�j��>�2A��[fH��L���w�a��zB�o뭘�J�I�nG�������$�:2x-���J� >Rm�����6*dj9�k�(�cV/�\^�G,El�?K�8>xyP�}����Pr��	7�C�a*&M.���[�r3��`y��D�Jn$�*����:_]n��%y�b!E���YHi���U���,�����,��=�!uː�6������K|KRA.�P��m�2���r�zo	9�t}�J��VFÕF�H����� �@�&Q���4ll�ܖ?�W�Ƨ�0:}�2R��zӘiR�(!�&c�U��j+"&�7iY1ku�i��H%�lX�8�޼$��g�%`:��@!u�%��9RzKZ�6b����"�;�+7^� ��eg��k�ae���%7*G�B=�+���f���կ:�m��{:ǽ�bR$����n�^H�ݤQ�����	Cɠ�*;"z�����$���<3����O��7�G�Fڦu�L.e�m�"���__��*�����[����R�8*_�D�� �=�8�F�d��]���h��l�20	)nj@h�ZIo�����}%�%YK�:B�ԖK�ͭDUZ�D�Q�d,��$�KY�f�Ջ��xU9�>�֗�N)�C�x���=S1�I,:��$a�kUU��j��ր��d.?�=W.\�ę��Y����(�r_�ۃܭ�
��J�E�g�䴫�m�`<qr�Õ5Dw�Q���ȑ�v�l�,�O��*�<����Q��Vr2k���kw0�F"/-35�5f~M$�f-���Y[��:{P&x��n�ӣ����3��J���on����c�\0dE؋pЊ�g	�gF��ŷ��s�=��S<��	�>^VOF���^bL+�6�=2;5�������&�~����֪`�_p"/`u�	��}���6׹����;��VLNbx�C$*U�(	�i,N�U$)�pU�/Tq��e���	��|������!�}���&���ʶ�k�e5f2� d��+bu�Iէ��3|���Ĝ`��}��&F���3F��UTչ񑴻pr� Kak?�L2����HHE̦�7�2�%�LzG����p)�����0iK� 	-�t>7Q31��V�~Y]^%�y����N5� N�eTݳ+BT3|3�v&��"����
�_��s�/�k?���V��;�c��q5�<	C5T@����x���^|�$�ʼK"v�|���_#u��w�������DS�u���E=k�N��u��.7�޸���� �/�ڪgZ��c����B�@3kEYO�3���K=����:�F�?�VVp��8Z]#1�+iYA-�v�ݛ��5�9�H����8=�"�:�yb���q�]߇Og�$�hc��p����7�^��S�{is+�&�QL�jxB�:D�[r����$���c�|�}PRA����M�
?�}�W|B��!��5���*{-O�Z�����0D�\Z(� �Ò&��|�f(z��@˰�*���͵+2qnn,��`����l�7���0��W.��Ex>X_}��ab�H�[��jU��X�����"I�.��g�ꘋ(y�e��4�yuJ߸Q��_�ԝq�`s}O�<F"~�����3x��M\>7�3�v����ߖ�v��/��<>����	b�r�y��z�]oe�l�:��x7�=oݰ%�w)����t<HN��62ץ��c��ɭ��|dIҿ��!���sm�����Y�M����z��e�}q|BB���G�V��}��t���HJ1`��3���C-9K�bBZ����{L�f:���zE��H�B!��"���1~�K��A��Q�a��9���ȱ2ҴC��F��Z�x�̼�(�5NFri����x+�W�W]�G�?�K뢒l��a����{G���=<y���'�x`�����H�+V��C�88L �|�+�P"N�Wsܥ3zFԿ�Xex�O�bE�h��ujmU���J�2j���:x�P��1��]I_)DH����1��/H�
$�ܖ*,�����h��N
Ā\˲�Ea�W&��D2�B��q��<��E���9F�t�z����f�i�[Ie۹���r/�|�/>� {ė2�/[��v���
��Nӈr�-�dҥP��Q��˔�h:HKh��U���Øi(�K�[/],��P�;�%�\Q�^[Y���O�f��zNObld����&��k�E�T<�̘?Ĥ�Ŏq����X�"i�{kvf#�v����b�~5�`�_��rΝ_����2��s�d�Ր�Ղ��j��\��E3$l�*+�ToK�F2��ii���/d�����F�8��B���ZL�`ls��R��9UT"b�lf�Jh�{n7�M_����=.�G�d>���v0�����4X���G�� Z����[ʤ��R��%�< �'q��H�L�(G]��<���֪V���ʕk\�a�8&�א�nj��g��,��p/^hL�i�0�*�*i2�QHgQHD�� �$��l�<��V�z�gH`g��by�_ǵ7�!��p���/"����XE|\��^f	�Sd��Vi�V���6��[EBl�|�x-6�y�R����@X�ƑK��GUͯ�w�& #2���2,>M�s�ڛ�����FNn�Zvóu\��ur�d PnE��J�6��.-kRٮ��ZdbQ��,!q��R�A�xL��b�t�_���i!O�|������o�&z��0 z�U��-���&4�-r�Y�jէ� ��^�:0�%-jb_)��>���!�A�d~����]�:j�j��j�VW��N�HG7qz����wp��ý�e[�L^�X�P,4f;dزe�v�<��_��e�WIg+r�"\M�V�Ŗ�f6�5r\�lb�A~��r��N	F8������]K���n]bRL��܋R�$8��(p_�~��z���]�J�S���������+�����8J���]�M�܆�=�ғϐ<�������DL� ,�K��%㳛����0`��um0Ж��Y�������(j�"uY5V�u%թ|�	����T��F2���2�It����^i��q�1�`=3>H�dA�`"��"A2X��PD�{E6~����|}��N��Q�կ���YA��W�sRF� @f�,v�'��V�n(d2�x��|M�r�$ǒ��� F�pXj���~��$��x���΢ȹ�}�6��� �s����b� �h��ݣ8�I>7������L=L����K�uU�^D��ø�$����ܹ�V�=|������\�ƆI�\M9w�2�z�._���Ԉ����o<~�Aڑ��y��c�(5q��5�'���k���x������/B'n�k��z�lю�r�Ã���v��E�WMn3�ZQ��#�%�i�LN�bgo[�����k\�|���q�Z��x<�����3�����V��˿��{o���2&L�I�X ��U��:�$�C�Aq@9]�� �R@�Wn�_�X�g~�ÝU~�"a>��c�G�l����&�N&�սa2IgA�Q�ǌ�Y���s��p�������0��_��;�Cn|,* Q(40�`>"2[\^"���>W�׬$	�x���L��d��\���1�����I_+���b�a�+OMcbn��S�DAfp�<��Q���zED�lZhLdH:�F�Ϧb���'x��K5o����Uf�ZR����,���~-]}�1�$�m�p�~�p�\�S��x��HP�K��=mW�"��6���Vµ�G��fli!Sn띘�0��IO$�3��c���UxBV8:l=ǝ�C�B�MLT�*������/��x�||�K����� ����@Ḩ-|�Fx�Ӌ��C$�^����@��6si�rI��I1���@$b��?��~H�!�k����{�5�u�2����`*��/���a��,���{7Z����́'XaR��b���y1+����ջ���	�{ͩ�>G�G���}b�.d�7^Ǜ7�cxh ~�	�:��'�X]�B�'�o���M�{�.���ȒdK�]�87
ɵ3䂇��K�*BjU>w���q�eފAr�}��u�t�m�����J�k��������\�<���K�<�~��>�;�˺�����\�t���'?���pI�-Y�L����E�g�qT:���v�t�M��jh���Y�h�����^L9�w�S|����K|��n�׮b~n�$�2�.�TU�i����pxt�}�i2���r�+:��uy���8{[�ܟ^��H������V�%�V_�D���c��xsM
h_hg�(�έWp��<z�N��.����2/m,�`qi/�7ppLRHl�;��)q�Z����g��`j<g'��vTKì8GP����ͥ�P�oui-�*��Yk���|�f�8�)ώ� ?'q-���g��0���M���nlnaqeS����&1��l�Ȭ]����]mbl������s�_3�������T����N����՗���������cg����n6����]r���ڈ�N�|E@@��f�w�O}�*!��7�c�F��u�tVZq�x��17�=��~��/K�p|����;o����&G��X��e¢�1,GL_�hq�Ę#�zQ�3U�3T�Vn�}� �&1�X�ɼ��V�k�v����/!����Ǫ�6rM/B#��ý�Uw��/z��5�-�**.#?M��DLB�gK�I۪�'@5�L"����_��>*��n 3r<p"�K�c6T������Z.
�/�Am4�K�r	W^{�CH��:s#3��TmPg��ړ��ШH{���}BZ��+�,J$���	��:�$�iy!H�:�g�uJ��]�K�mf���E:���.~��~��!$
u�/2*�!�r�/��v�Q��[.���)�A),��i���ǻH�o�\�:�(:6n^S]	��u�	�ɮꄫ�$�Y�߿��-&�^����06t ]�Eѥ������'��u�Lå0&�� �,��Ғ���&I�ҧ$G(F�Q/e�L0q�H�m��S��G��we ����;X��:�k@[K$��Yk��Fz�I���K��*0�5��JG���d��X���w�x �0�H�kIx�\f.nP��Nkr3�����毾A�zƂz�+��-��r`1����j�Q%�=o6T��"�C�����=& 99D6��bb��6��.��ܬ��ΤjU�����!��$�HUq$IM��Ŏ�ﾁ��E�Wa�k(їa���[,ݖז���6�p2*�!vK�=Ѱ���x5X%���S��d���}��M�af��b||Lq��K���Y�Ƴ��?���>N�~r��")>�}���@_��a�#�n=�W���d�M-c,
z�m��}s�)�6I,H��\3�Yf��Һlљ71� `�y�h��0�� ��jU_n,�'m�13��\�[O�0n�Ur+a8M
U��(��o�8�]���\e���c�����A4�������-�O�2���cE�`7[��(W�}�bv!?�����//\���+(��Z]%[C	��lk+�z��͡��-wQx/>�#[���p�{��~���E?��T�w��I�0~����ڋ��r��G��k+�����Ϳ��Od�w��3dsi�S+�r��d#P;���3g�]�%*p2��3�cs�`>�mM��l�>A-}���^��E����k�p��?C�L�C$Zq�T&��,�������m<y��{_~��t����cK���@�;2J@葶���k�s�r�����
�/��ߋ[W����Zğ��1�Q`����X]��_���
�"h%���:x������O�1F��?|�L!��c���u��D�*,�:*R�V!ò��퓑���OC�KZe�]14�%�E���ڰ����>���6|1�q��<^�r���#��1w���l��Z<vU�ΖJ�V��o� {b&�9�ȳ��#W�5Q�sp[�@ֶh˭�D��oauk�����_�:s�`�!|.;��=��3B�٬��W�մ�+E�F#�E�J���t>�ٸŭ
�k�Q�Ԉ���J�'�)W�U����_I�Ǐ����1��87	'����:��	���_kv4���Mz�k�iZU};��`k������)�|�٢�*6��R1�=l֫��*� K�6$`@�SCL���ܿ����G�7���ҕy�pnR��DoЅӃ��7��?��?����֭�x�Ï���/T\O�=E`���"C x���33��9�]�@((��$Q5�J�QEoOP����s��m���7޾�w޸�ى�V��&����K����q��EƋ~L����_�����ǳ�;� Y�"�8��&�f��9'�w4�T��1um�D!�)m��
���.v�6�ڝ��?�>Ξ�VmQ�v	!�W2~���~�����#�DO�o��6\��X�X�>�Q*$�1�$���I�����Z����O��M_������8�TF(DMzgw�E���;$�?���x��>�Dׁ��%������k���9|�����~��4:�:d�>M�+Ő9ق���@��X� ���p�mE��IQ�ޝ�i<��1~�9B�Q�����;o_��h?�$���3�� �&017�B,[˫�����`�X�a�>^�8��i6����� ��%�"0%���4��yO3�f�I�ޛ$�C:~��>�مq���[B	�ub<��gG�έ��⫇��ǟ��Ҧ
&�v۰��b*b>���ؽ~�C�5��5����,�2B����s˅װ�^�m��ܷ76U�Bn���W�q?�p��YL��1?3���I��2���ť1�2���C�PPΣ�5�R�1����bU�A�}Im���R-q�0d���z]�X��G4
��H�>��k�;�^ǝ;W155��0f<�����P��d�%�/!F.�H����Z�6Y�g��S����(�hv�sn����arj��n!����r�Ĳ�xCfk�4�&���.�����0s�N���&J&[�����8]%�9rQ�!^+�EX/�/����T�u�C��K>-���������ݵ�����*K�����-U����t=�:]��W�SDi�h4T�Gn<|���]��q��U�i2hH��.A�)��jx���M�o��[J*�%����
H���u��o����h���|C*[>���Io�J�w���*�-�(6j�ܰ��Uav�n����!��(�U�A����\@S(�C�E�Q�`rv=�$bY�?��~�y�7�:���F�%W�J��TWf)t����t�j�2���� z���)�q����؆�ǁ��>>BID�z�㆐qi������5������T^�p��(�J%D*M����nJ����0�l/>E&�$h)�����(�r��l����ZA����!�+�qJ���ez��Y����K�fۖj�Ő�V�"I��Bf��1U���I3D��4zr�ĸ� y���:��1�ӶIC����|����m�DZ{��$5)��e1���42x�H<d [T�d�G�HL]���t�h�M�H4�`y������2�7��r�/��ˤ�VR��1q�������PR�ɑ$g�J��%H{� %J���@G<��9���"���*�u=0�~�i�kHEMڸk=R�!�����9��$t;(�Nx�Mڲ535���������>����~��{Z����8�^.��W��$��ެ�om��3:��㹖�Ϊ�,H�4$Lڒ�K5^f/k�bG�8��!�$��&���Ї{��Ϥ+dlff���t����I6_��~�����d�1��Ĕ���I�8�� BK
,R�T�e�1�,J�2��s����2E�kXz���-庶�x��&��0��$�=~4�%�v�}ް�4��^�C,��"��!Gp�����c`v���X:����Jw�%#�m~�TY��b?�2�IU˔����a�A&�n]���׮��I{P�'s!��G>�V�c�.{B:�繗y��d®�<�f~���7�!Pq%k�]���p�������V�Q���	���0>�C�{�}|�2���Τ�\�����s��v���S�a�p�<�LR����T�k����u�Oa�̂���K��Ÿ���-����~��k�9p�5&�g��6�N0<9�w2�����In�H'���$�2k^VU�T�����������߸����K�2����|��KW	�<�-��8�IӚZdT�5!��7�4�;�u�_
m���
�}��>v��k��gh^��~�M\�8A��Ĩ�?.87H��>C�����V�Y�3^���:gN��~��)���&@
f���ﴣ�b�d�����{;[���/�����^>"X��$912!1�3>;�"�r�j�;I0�mk�ư2Ke�t���G��Y,A���s�0B"@��p�!�i��c�{���j�/]:�!�+�7a�O>a��z1:>���L����Ɠ<g�e����v��km�Z9uZ��#��5�Y%I����0(_��*4"�&u�ݖ5n�2
�u��Hҹɽ���12؋w��:޸���~?��.޿�u*㐱,D"7/���.�x�����8���G?�W_/ꌪ�{"��b��db�&�!�w���M2[���n_�m�����������7��wn0U;�׼2�|�K'���?�:�`hЇl�{?���'�η��k���������,4*���G{ڪ?==E�2���M"#�"]g����H���wv�U���\;71��t	�]}�GdvY���Z��hvvF}��>�w���}�=��G����L����p�N6S��Q�kU{4w��M���+/`�h�vlC�Bq���(��[���q�gz��˸��M������P/����|1�S���DH5 �x���������[���̄���E<y���Q�qa�eǈ�P�Z0�#.���lh;H��%E)��#!�����^-�3ocvf�ϱ�_��G����ב�a�ՠ
i� ��hܼs.�|!��fQ���rC�`V�;��B�k	��F����j���#<�m�u���2יOǹw��\~�N5�Tt�� cP��!��w��q�x��*�X�R[�|<��
}Cp���5N���h�[
,2k�>v����
]������k0s���,�L���p���8q��Y����8�������g��}̵ܫc\��r�\��q�eU��2������j�؅���΍�v*	6P������	�m`}��e?����~�Dz�$��X[y�*���X�Ź~��a�Rp�;�+�++J��a��6�hg���.!��lvG�)&�3�`v�Ǆ�ۈ祕�]j���.�B��c{s�����!q	�}�����U��yW��e�I,^SS���������D"��g �=�"�L�׶�v� ]+	�R0n������+P���]��W��ܽ��h��xr4J-���ۨ7X��'�&�,�l`�	3'3�[oTl�Gp�I�6Ak�@�Q��c��ُ��[G���Xy�DM�_�=U�I$�
R�du�n�����}���7J����Ď�I#��K����	�}f�q�=�!ܾq�c��?�H�5��bnJ+���}�JP�n�:��RH�T`T��n�`Ju��[h�K��K'Q�� ��"8��bj��3�z0=1���~d�q�H��":�)j��|�@����#�l/k��ln��OO�^�uh��_[�چ�R�hw��]�\������{*��$�\3���%�I�����o�#�%�siU����ut�K�̋��&�q	;�_+!�z\8�p^��[2�%@R�]T���7K"�r�d�2�%A�@�c�ϐO���j,V�,U�Q��c��V�|E=N��r �'+��u�q&§���%�aQʫU���d�c({vLZz�eҖiW�%	�O�U��������~r~��P��~�̥>p3\��3sڒ#���m��cǫL����;��;n�~z�<	p�6d���V�d��xQ����NC�d�TT��KfMS�c��|�[$#���Ƿ�{S�ŖV�!FҵM�S�𣟘�"$�lN��V6A��{����t3E�����(����� �+yc�Z@��a�+sz\�,o�`��m�I,,����A���\>w�.]����gJ!�_�3�[TU{{<\������=l��Vs$L{8�]� ��`ojr�k�=Nf����!�s�����
�{:��7b�s��'H�����㳏~�\6�&��!i+j˵�瞝�����qn}���>��.�S���澚��K	ʚl���K��D�Pֳ�>�5ޖ�)bQ�;���I d/�: ��z{¿�bLL��=�'!j,:�X'pumE����4^�:v���8IT��c2�S�@�o��H�� S(�ͮ�C��ēŗ��n"<ԃkf�,�=\�g�cxſH�)IDĳQ������g�����ގʜ�1�����τ<w� r�UP��<=�!�Xm�t����e��16��Of�k|��]�}��=2>=3��ko��n���I2��iRI~?c��vm؂VX{z1�?����O����p��e���A<���9�B
Uv�13��/�8�7�Wn�T5O<�ĳb�6n�I$�3Lޙ�>�0���"6�^�N068�˘�CPv���T�)mkj�+��1�QϹ�'/��i�@�@no�1ؘ�d�Q�R�#,K�G�����3D_˙K�t������L.��_cg�%c��@ʇ���qS�����X^zʵ �<�7~$%�s��	���s�˘��Mi�9i3b6v06:�p��cRaV�"�_R��6�Y<(�Jl�&�ޗ��pm�{�_��1;;�O��9��3�Ǜ��!p#�wprz�X<���}�U�3����I�TD&:n�v�����A�S^.{T�U;e���n�.�VE�����"��K�'�8R���q���NO"ĭ�E@�_���2�	Z]��^t��a!�_����rq�|�[����{��]������HHĘ���`w���
&&�:_����.Qh%A1�WH;�Ϡ��7���7߽�6��?��G��Â��0&l�o���{f(����c����o�.]���_� I���b�s$����r�8|p\�Y��
���O����^�������x�G�3�������ϭ�����1P�a�8��0��/����x�w�g��]#�Keb��>S'���%TeR|�k��
l�t쨦6���U�}��%�檢(�3��O�r��i;�G~��s�����tNcjN�4֖W�x�~���T����w�|i��b/��1ci�������ׇ��`��2G:�Z��v�����Ƴ5���,�^��x��>1��[�:.�\�ť���uF��;��[��1�	��\
�U>���5L9���݆�T=�9Dg�̆���|J�a�R⚶T��?4����.�Ub��n���W�b��}����c��֚�+NL��w��x���GX�L�D��:�� ��ha$N����:�;A�t��SӰ�0:�LS��\�`HB&�]]x6��y̥�<�g&�1=6���Z!VY|ʼ���7�*�!���K�8:M���I�5.ȍZ[�C��jē�'>Lr_tF��-h�ӵ�g�{�E�,��o�������[ߺ��������W��Tb{����}�/��O0?wK�[���a�Ա��F.�U�%��͘<�Q�dߕ��$�lX�Ʌ�(�;��roT+�Zt�ϭ�k5����u�{#�]%�Ĩ꫼��7tV�����ФM4Z�j!�Ru�2L��䊈�x�fF���-Z,��x06'�.�S	�+�Kc���d��k"(_�_���3�OTo�ķ�f�l�����5��r�I�4�N�V̒9����#�C�`j����|�6���OY<C�\�/����J�`k���rуm4+7��FPr6�_mJ��ET��h�ڗ�n�$��	(�%PK���>�K�Ӣ��!�g�'�/��Z�����Q#��m<hkK�x��3ؼ�����bGA6��z��F��<i���K�|bf�MDQ hJ��9���d�!+><������XO���Eb:5��!Y�l���w����!N����AB����J�DԢ�4���ll(���^�x��[�7���Qk�YF)sJº�f1���$0���>LE���ش�����C��2�:�~3N���cg-DP¯�!�]G�-��Ѓ�|UUf���n��t��<O��	?G�DŬ�z������qz�:+"��/҃�@#�#�s�&�X#�ُ�H�>���9����Ƶ�/��z
�vX�МLԝn&;�\��g@�@�H���-	��k4ƽ�#�%ܣ]��-��G�A�{v��GZ��Q���7~���'8{ݩ�3R���Za�fm��.�n[v�K0d�Un,ċK�3��.R1�����aܹ}�����������Ә'Hϑ�>~�H���Bp$A����p71�$�l9�ܒ��\{����"/��RV~6_p�܏]�ي��$-5�PX{]�m���90����޶nm�\�C�$� ���Q�;G`�t�Q��z�w�A`91����{U��
����R�FJr.�#qr��VB�eb�}�"s��$�y�6��|�|�����%	ldQ"�=|q�S��+W_���7����N�E��Ruơ�y�]'����&I��˺T�E�^�V�]�^W�5i�T~O�#��|�dO�� 
0���*�$-��<�����wb� �A<Db�e@��8C�-�*�b!�����0����	b�b<Ge&�ґ ��S$ e�:�Myv>���j�
����}u��0���m�bQlm"�ͪ����x�T�a��Rf��"�A �N�{edx#�8����E�B�k�z�dvC&E9�bv*��ui��6�
�W��`����w�Pf046����_���#��[��2;���T�X�����~	��0!+^�I>�(�ט����Sbk��U��6Y�)
�b͢PQn��b(,ʏz3(@��@d0�J��]2O������
J�������G�1��/�fg��En��<vV�xf$)7168�d� p�t�{Ţ�!k�OԢF��Uޓ�B�'K�x��{����U<[|����7޼���㞿��uLO ��F�c��TZ���.��(�/�U�������P�B�t��3$Lߢ�7�ߧgH���@Y|8e�+W(�m�� �MS:��������V�r	�����{ek�Γ�4�˒��s�ز4��wx�W���ɓ��ͼ>�����,<A��ط�j��}ձ$
�b*_oՍ��a�!� U�����"Z"�;77�sg�h[.�C������uYl�շ��x+�"�^;�~�?�_����%�v�"As��0Ug!z����m����򼥙g;$�N���!b%N<{�Ƴv½��������=l.=����p}I��`���o ��3r�g����sxo��:I�6�;��H�3�r�n��jkϳL�k�K.{Go�޺:�����1W�a}w����`rX�E_��\�/��O%�$�Bq���kll�����@���]�v��ϭ���:Iv���H:�oxJK!Ln�d}�*Vfm���b��!�=a��ӊ=K��H�1�s|��CB�"fg���_A4ޣ9si�1�$�ǧq���WWq�H ΜX-�`Y�g\�I;�Q�#�8e>���ݪ���+�:Ob��}sqaF���	��Ƽϸ,Bd2��c~N��I�"=����w�[ ~q0��
�?f���Q&��v ��ᙗ�h'\��:�-�D������ղ(M�4�7�ѡC<����q`qyQ	J��We��b���-��U{mcgM;�~��w�K���_ O��P�{Ml�d^�՘VA�\��M��j�ZY/)\wU���!j���5��z��H%�����w�Yn5k��v(;���y\�Y��ï�gWq�������C�AL�?��|��Y�����eV!�L*��3�a�_��Q9W2h7��$C1G�y�K�?NLkҎ�ɔܲ�1f۝��1;���$fg�P���n�l0_1��wr�$�lsq��_��{���Ϟb�کG���&2������,p��
�����M��>�)-�r��("-�VƯ��_3������z铻_�+�Q�U�a�U���Z��(V&�V���>��a�*�z;�-����WݟB��A�Z&�f����3���j�hTs��.�2Ԋ�T��@N&)�ˍt"M0�����( 2�ad,�7`7����(__�		����e�%���}d�;<�����ۇ��쎪�\�|��У��w�jm�C#	\!�(դ\:��]��17g�#A&�1�GT��� Hr!N�����\\��^@�@?b�d��+8�]ՙ���E�B����ܡ_�:����W7�";.�(�
ⳗa�IGQ��`���E�����j<ԧ�hX\p��H%�}&oqn�'�� F0�`v$�ӟ�c����ǧ`����0��,�J�� Sǐe�we�4u�Bn
dT�F�JVon�]�(�l�>?FHz'��?����� I���`sm�ϑ��4�W��Z&7r��/N2�C����ԃE�;ZE2nq�bb1��N��3�G�&J��S�8� �#k�B��I�	�NX,j��P�¹�Iܹu�I߂��cGS��l�;���]�y(���ןڥ�dl�n��77t`��@�5Hi�f(O�����4@���IM��`pp�MbF�:<F��gx ���x��=��2I>O�����A��y��+�P���Z%t�M[�¥��hMS�OHk�u���̿�:f��\�z�/�Oc0��P�a�gf��6�ʎ>֭�m�5CL��8K�-
Yn�~��;��ZL�>� NB=<�gڣm�f��춴�@��f����Y6C6v����΍��A�(i9��-�G��D�ߦ&'u~�x�{����͟]e���ވ��b$�]���*\�pw�N   @���IDAT����OPZS�N�Hqqϛ�3��tj�Z:��9�%)M�|�H�C�L(Am���pfSb�{���}�<u���3Q%
s���^���ġ'4��g��K�6Wq��Pq(ô���<��$A���Y�z����2�#*��b����r{\
!]������j ���c<��%&�LD�|�Lt̆�$�֣#�8;O�/�8�ŸTY�_A��9�*�c)g��˜��:��do?"<G5)4p�դ���U��s���Ǚ7�����>ŏ�s��C�0�̌��F�W���K��q*�U ��i�f�����%��h�yKZ!���64����h�7i�J��Cc����J�K뷇�����a��;������W_��x
�0�׫�%�|����*�w?������_�p����p%ZT�ƚ�Jk��5Q.�����
�xUPy�V׍I+zf��&-9�$��뻈D$.������{�=E:D��N�ٴ�ʥ�׭����YX�6�r!��]Tze~���=>P��e�Z t?���H����� �3���=�9���B����{Pb���-�p�O�'����E�k	��k��x���zkyz����b����N1�8����K��!�Mk����gQ, ��	��z�����\�3s�83;���W@������MTe��@������{�|��r�nC^Ɖa��v���{�QQo�t2�`��9	����l�_^��8�1�;��Zڴ%����ɉ,�(?��y*���l4�c��#0�<���C�Ykk7N�U5!Rػ����9W��=�Q���_C�1fo�X��NH|�� �K�%�2"���L�ߕN���>��Q����Z�e0��C��8<9$�@��jh���4�5�k����յm���WK���?�k��t�\�r�h�T���*�Nύ�?`�����5mYK1��H�<�L�G
L%�}����k(�?~�5f������x���>�VKR;#O��zd�m����q��涎�X
A���Y�E��-�����S=�c�|�{~�_��<�Gk�[V_���e��,�\^PK�-�����z�ƀ�J��}VU��_+���J^ ��ys���R7�X�C�jŊG�76�}i5@�S��t��z���yr�E}�����Ux*�M��~�ɒ��.0g�J���j2�R�Jө ���/��X�U���*���;ۇ��a(l�ى+�Z��"���i����A�^/lQ��*b�?� ��Y���(>��A\�x����/�P��Q̥����!&Kgj���B���*4u���(���H�o�slVB����f�`Q��T�'���D�Q&�H����� Kk/��z|b�g'��'�c~f7.����s�jף�+*�خWy�`�'v�9�
?��P�T�s�����*��)�.\���̏�	���m���Yȶ'��1��_0�o�c~�^|Xl�K��Xg�E�:eƜ׿�����@������K�aq�z���2�/
�bW����F>�!��vlos=�/��q��?���Y���ß���<6vcC�xD}���]�n����"����DI��P�F���_�x��m��Pm�sh�to����d�+����vPZ�n\��P�A֦^��py����_��/�]�� �b���K38�0��Mܿ{O�^S��G�u�R9��f�����8*M�������ί���Н����[ek����3���*�U�A	`�I�#*ic=�xn���v~����TH������vv0;3�E���
f�16>�/,�����F&�鵮-�1����1*o�d�����82L,�2:9���Ȱ�}�6J�C��G�56D�'բ"=���K*����Q�y���Բ#���M�����7����sm����eSȟ��`׾G��zƈ!g5���r�ɪ�/AW��8�}LV����eU�! �I�=�aR�S��ܨrM�#�<`��������gS�՞ʭ�+��"�cb��$3�F[)�e��``�T���;��������+�@	��w�����pf&ϐl1���x
�	�>�\���TyT��͡�W�I�R��Li/��nI�L,�Ҩ7
��v
��;��U�������")�ְz����)���҂���@�)\����	���DE���ސ"<b5L����q;(�Z�KޙT�D�Y��$��.]r�rI�rd�w0���	�m5����a��+W��� Я3���c� #E�P�Go<>^~��g��d��IPxP��'�%�ꌶ�#��9�F���׳h�V���A!�P!��^נ��~�[�;���Q|���x��v�'�����b�?B�Q�E4�$z.I����3�Y��c<)e�
&��#%=��7�R���#��e@��f���$���2i���N	N��(��2'�r}�_�"���u�|����E����/��q���z~����n.>Sϯ[+D���5o�"��"�ْD	�0Ji�MbT.)���V'&,	v��d!���!Vq��������E�����Ko`����uY�X�?�x��g�����#��⣏������dR+�W�w�}����ںZ�HRH�ln��j�'�h�r�$r�YOHKS��"b�)TFZ*�B6�G�����EMJ�"f�Ը�&m�)���f	.���M"h�v��$Q;�喾m(J;<j-����!�N�
�LO�q���'�X�ŕ����(���=��V��8I6`q���9�%�!��a>����P�Y
Z �#9c��d���*Q���j�jR�1@px��ϔ�9��1�����?���76ћ�2cf�����%7An�H�����c�����gIT;8<N!�or�:w)?_�D�\=T��g��Bl �>��clԄI��ܸ�)��~����O��"y��|�n��s��E�����֙���8�_�:��b�K{���^F=w�ý���c����*�c�\�^��մU\��O����ޗ�y���p����n${�����
�	I-z���k�D������|��le��f\oa�d̅6	���En��'t��;Z��Q�\��_(w���󖑟UG@LΉ7�^"����W���e���=1:F�eaLt0t�M:�dnK�F,v7�i~"����q,-m �9P뛲�Uf�Fۜ�Y��6�m�Ce��d&c�F��&�H3�ģ��A)�ܸv�"�z{Uu{o_��(Ia��Zn���,Y�Zǅ˯�ʵ+���"�~Q}ڄ����2>��MꘈQu�П����̝����n&��j;�����
��y�&GpnfL=v��u���s�7�p�����A���ވ�-�s&?U���z���ܩ]/Ƽ��\��b1&�pZW�^} �[A��S��ܜ���pء��k��)������۷n��R��"	�tQx�h������6��^"20J�RU=)4��e�p��ƴ��K��؀��6�g�QϞ�h2�8�^��"���|�<I��Ξ<s��ף�If�ŢC�����>���o���T-�V�gBT=e�����H�Ұ��h�1+�>���x�r�H���toP����>c�2�놊�x�N�.�1|B�3,N0b�%b�X6�@0���<f�&K��u]o>#6�*�G[ým-r��̎���D�D��i J�����z���6[�3��b�������
�vR����PkUq��5��9�!�$W������l^г0aި������u���6�f"���}A}O�,���Q%Ϊ�j��v2Hq�=Ƙ������w�"�J��1���R=�&y���^,?S�iǎ�Cp�������?D�Τ>�Rx9Md���,�~��])]x�bQ5+��l�-�gm�xς���p|t���s�OY*e�54����c������"&	gM�Z���\�%�uQ��(W�SD��pjs��SWF;@UЬ�Qx���6�n�ݛ@%��"�Ο���é�M�|y� f$E6G"�M&�r�ZNF� M��x~oܺ�`�K���Uɒ�z��,��n�>'IVP��K���^��pzH�t|@��C2iR ]W�<��;���p�����V�Z��P$`���r~��	��2���^y�[Fz�|�>�<G#���8�3Z�n��O���t�g#��ֶbH�����u��!zn�V1� G�6�n��u&%Ֆj$1���?{��"� #�7�0��T��T%2N�P�N�8|�'�1���A\:;�X�)/�\������`JuC�[������b�*`Rn
�ʢT'7�n�B=�|b���~�L�ĸ����2Nc[$�Y��9��c5R�+k?GM@��"�1:T#��NL[Y�o6ۼ�n��_�e�Ah)&Hz�d!jG�t�dBd{��Z&��>n���A�R��Ag���b��r��������!*_|�KI��tğ1����(�-m����1s~�IF<�l��*�͢�y��X*˱�c��3L��&mm�2|�H�z��p��``x�]0igdJ$L}��06�a�X�%��nVɐ�7[F�O�e�WD�Կ�{暵������ԭⴵ%�E  $����;��^�	3�IP.��p���W���KU=6�nU�:��B*KL��R��p�i�W�u/6�ծ��f�9i��|�oJ��3蔋=c��.���-����?3�T,��aT�w�DF�k2�.�^�O$��e��i�ONp��0	�(���.�Pb��������(�I`�J=�NYf�ۆ�j�XP$IN�Wom��F&Siiau��["��al��D3@�b�3��7n�P��ŗ�d����J���`o@=��h],����F�)��Y?��˖n�����;�%�g�m�J)�+�܈?�إ�o���?��Y���	�M͐pT"��,�$�{'G8��cmm~��G��w~��_�?���/V��P��	(z�ݤcN&F?�1��"n��:�
yH�+��x�b+n]�R)��M����ת����D�m~a����Q����C<�dB]VSq�Ů
�%��Yv�*;K���0�H�����85g�[�Ig%$v��M �����R��'�*I���F�����k�p�
��������Ξ�Q����g��w�Uf}l�Ը\˼���
!�"_�%!��f]0���YL}�fi�)!�h��ZGo��g'�5�T♩��Vi���`� ���Ob���6�I$;܏O��Y��7����	I���:y)��#�+��P�.Q���X-6v�S}�(j�7���y�r��	6�.�88��/>�m�i�|��ļ�f���pae�9y��B�p�<|��́)Z����*�1u��C*�R����y�Z������D��r*�7����s�����'4��b��E�3n�yn
<�n�s0Ƚ���ʜ%.bvj�9��ݽsLY-��Y���9���іB����n���e�;��YQ���uEFD\IZ[c$2^�/��/�>���cc�:β����pP�]"�A����!�v����EF��/cb��Vk��3f���ߢl�a�-JW�D�;�\G��(U+�}��;�b�H^����:��Q�y0^�pQ[�SQIvbqq^�/H��%���Α�������ҙ�!���e̶x����_v�����yw$�>�M����.NON���;;5�K�.jLL�c��#���
ZOO���<�>�򸊞��X;�/,dOZ���T
�&C�NnjD�O�全��tȜ�H	n�^�0n����!">�*�����"}!������ �i��#�����`��}�u�8��{����D��x�J[(2?�Vͩr;i����r�dQ�j)\�*&��	��E𿲲��aΝ�F���0V�}���Ke=7��+�������k�p��9<_|���>b@��������&���	W�rA�x��c'�t]G$F�-��*c��n|���t��>�2�	���*#��{-�Ⱦ��Q�P��S��Ë5k�"��}5�Ȗ��H0�Gn,�l�1'�k�S�|�����A��ו�y9��/uι'� ` @� )R)�$K�7ت���u����v�]ko��WkI�(����Ca�`r�����s���߀�.�jjݯ���/�{��yк��*�q�
ٲ4��l��c�<�r�'�(�����>m9�O쐨'�G�U"��������$q*4P)�n�c�1e�ʬ�Ȉ�~��1M<Totӭ8���$�~��
�i�w�gB�Y�O�?�����ɬS)�7J*�"-"�R�{E"����p��=>JK��L�@l"#�D������21�L�%w��Ȝfڭb��-	"�u��ql-L������z�q��%�~���bg���.�H%�[Ek�m/��lW{@��5�E[�.Vt䞿ŉ����y2[��n99��o�a���\����Hыl���3�j9�ِ���f8����jς��HuA��2rB�Jb�BBQ�%���G2(��Ƽ��5�>�O�C�wBF`�,��7�N���Eb(����6.�yct��]����dI`̖�J�+�UA);�94"#d�Z���"����4zoO+�C�Y���+D�inzN^07�W��A�V����Y糧˪"�A"s��tZ�|�y�w��V��@��ZM�D���ʌ:��;�xy<�4E--N�,��E�bhp��E�o�2���0��.
<�"Đ'�Z'0���d-Z�Q������^���	���ep���\̚	4F>�|���I�MSò�F���l�']��Dn���JN@o'Ν�˗N��&�`L��3=~pK�_[4�6�K�ŉ2�G�TSTI~2��m��IGy�3�`��g�t�Dc$�fYo�?���h�`�L������4d(;A��YA{{+�D�JM[�>��n�m��l&���{�z�/�]�#��77�ꂪ���;�3Ё��M:���X_�P�	�m��؍Y�"��s#`9+~vQ@k�;IH����j}���i���A�&��%�{;I�;2������:J�Y$�7���̟���vqm.7 }������'��&F�Z�@P�i���R��U1�(K��4�K�A�$��=L��^�-~n)��Y�A�3�1>��A��"��2V)��p�7xֲ5\����>U>ȆH��j��U�D#�k	�^�H�e]��+Gk��^H��ZCJ�l$�~_ܾ���5�"wv��G��$������١s�=��O	��h�l%�7��+��X
[<K��t��}8����ծ��f�3��hdEe��L��~������?{���Do�ɥ�v�3/\ֲ�ͭe������#6܏�'�$q%�U���N�F��):�8K�����f�Z"�T�A5����#��D9�'=5ü�lN>�����D�F�� S�?F;�WU���n�#�?�V�!�9����<����o���ҷhi?�>:�>$K���Cc{[2*E�հ��i�ns][�����9�o��!�lV�rką�O�y]<�Q�T5H��]8��GN�����(���� A��nђM�ť�]�1U)�uA$܊�~:��F��2ɒ�F@E��Q&;�����c$�$�l���?���Z�7�23��KϠ��6�ۣ6uc3�#*��>Cb%sO��<�\���$.�o~� �ى�bhfJ2�>�G�7���:��! p���d	N�2@�{,v�J +�:~��RI�Ř�o����&��~���!E�!�"��	ʂA7b	�f��-��ّ�!�m��[JUKNW�]m���a�𘝝%X$xu�	2chtIdz"AXyܼ�>V�g4�褍�C8w�W�5B��" �����9�R%��x�hmm��D,���\�C��\Z˸�$�.O ]=�&�j��fvkk�
D����FtD��=�Ǐ�{����6�O�(���h�۰&8~	���yy��g�09��w���W�I)X*�2�EH��(f�Έ���j	�T!7��ҷHu��iV.��J��?������`&�M?Ӡm����s��N#J��ծY߀�(Ah�	�q��iܺ{��<ѳ{��Q<�����I�*��硰�{�o3��-$y5=�r�ed�T��h��<}�^Xw��W,omb��^��q�dz�D4�Hi�@GW�~T�G�c�0���Y�����{－��u�Y�]�?B��4!Z"�#�oB4��Gz'�lK�aW�w�쥓�'_���˭����+׾�^U�M��t�S��SK��R�.��!��Wז�ic����*�dVD��w�M��e�-�Vb�T��4����{I����5>$���.�Gpx���SBGȍͥI-�n������,I�-��M���o��#��4t$N�v�u�0�#C[���b�|�-���"ΐu��8(��� Y��6�l�r��- ��HB����w��k�[����k_��U��7LA��R��{#���CC���C���rڸA����"T��L&c\C��U��6��-�E����)ޙ-�w��������SH�<�j/�!dIW7H>h|>'�y��B"���ߡj�tl	��@2j�����_7I߼�MHF��4D~�7K�@M;J��Sz�qPnh10����܋������'�hu����G�=�$1]Et+�3v3��h��,qA>]C�צɕ�L��'_+�T_6x�K�Xf����}��%	5VM&�re�]@��;����\�#[����C��e]���F#J����=u��F�Ϛ�'���?���QB�uҖ��f-�I9�f�KG�H]��_<W��o�|SqL�_�2F&F�mMr�b��դ����iީ�_����U�}��A:WAa'��R��i_ۋ�T���IY����̩<�o�`�'I�槃������3F��QoEg�C�l��Se�$A��^ ���rGgn���T�!rn�S�c�{����Kc�S�+NW��KTK���P�xȅdnmmhL.���7�2��,w �֎M狓g&�(���'�(屣c��� �F+z[( 3�w5��i8�N4��ڏ$Y�y�w���]���02<HCsO�rE��&m�ժ*_�<996:�����.�����I�_%a%�*u璡����Z%�_����i�H�D���gE)���z��-��4�U�A �`�f���*A����uɥ�Չ�l7�eӹgk*�zp�G|�88�$���H�hl�\��b/I7�^J��`��쩌��@K�O���$��
b$FIdqDRo.k(�Z">$e&Rv%e���)kY�����a���k�C����et��Y�ҥ!�E��ý�j�@� !���Y]���������q�N�m�h����	Us�]ƴ{�7��I�"FK�8��u�2�� �碑������|�$��&�d�������Lh\�DQ��yi�Nc3����A~�2Ax�4����g�wI�c���8��"I�5�[��\ה��AɆ�Ϋ�D2#!�R� �qx�և�����q:��왓$��:[�|P�F`�I@���^��/~ż����9����R���)�G���7$�U��(5U]�� M���_��.cd ��g#�`��<��|�Z��hwsK�I��T��ni/c"�����C�J���U��IϬd�����g	���rQV��l��%v�|JFǡM�f��p���F�����Z2�<�~qn�D���x�̥c$ ��8E�a���=pt"F��1��7��1)i�gi�eΓdV�q�[�d>��+�lA����g1��Vf&un^�P.����E��4;��ｺ��{�@W� Ə�@�i�ݻ�yFC��v%��`��G{�eޟ�E�C������R[����?���=4KvS�`/�OGN]���XX�ŷ��m<�������:h�m�?�!�):�*��\舶�ؑ�:�=%��/���
g���}�B���"R��̤I��ѝ�bd����0;?�/}��HJ����<��vj����T�O�LO�ke���0;�-m�viO쓙i:�X�$��|�"�s��-BD;'=ժF�u���J��J��2��a��˹��p�S�1һ��v
/���9	I3�8s��m��nW7�iI	�������8ږ��'�ZZ&����;�[XYOk�uttG�������.�Zk2���vJ)W��_�ǅSG����B$��$i=�'�m�lo�c��#�+گ����8��\�h�bi "S�'���������f�I%�&%��s�>�y�e�ח��uN��
���!f�I�����|�D~"���������{|��Etutb}v��'�G�F������Tk�^zy'\|^!��X,�=�
)=�V		��-��,=�R�(���TM�j^}�26�<�_��o��AgW�`�Y�7�Al�ddK*��O��`ye����ڗ�F\с�����T�H Hθ�_�k&ݿ����{/ 	�#�ta{g��ތ�xo���91���"�5��."|���@$��ƺ�V��(��|6��!=�U�R!�����A���>/��OJ�-Zx#q��t��@��w?SC(��~����淳�t��/��$pf����h��ۇR�BbjS�tVs�ʆ�CW�yO�x��X���]#�����>i1�&pPګ����0f+�!���Z�&$����/YqBG���ّ��e��|M�E��D�b�3ڐ�T����ݳsO����Zb��?�g���(�n:u��dS2�[�kԠ�(o
��ZhK}ĕ,s��KK���ä��V�T�g�U$b;�w)��0�z�w�A|\Ѳx)׭�ƥYI��[)�dM|߲1�; �Q��~/�� �����+܇T����hqx�!�[�뤼��qh%�����u�Ա��Dl2��<�k.Bh͆b(W��R���uU�D]��$�A�ԓ?MŚŽڧ�H��]I�V��$�ii �'y���nC{��:�v�bk{�w���YQ���?���u� �� &g?��2�,��}v�U������G}?Q���]B�dl�9j��� b$��S������}�}=u�·3���>��R�\��Q�j�̠��
��������I�rR��W�"�JU+���s%XH.��.�*;�j� ��ף#զC�=��I Gq��M��鲈G�e�X��l:���	u!��V�%��r�L:g�Z�"�@_�A���i%��H X�A)�1���y�q�j��n(?	��!�h���z�*�g��!���Z*���͓�^�!ۻ:�ۿ��i���u���.Y�?�BE:��.��c[�*�>|t_ko催� ��l	�TJ\{h��:܀������|b��k"�l:��A�����ݍ��,����,)qn�U��P�� 	����څC��D}��L@#dB"Xe|��!�R�D��bT
Z'��:��O$��Ԇ����D�V�S��|�d�įA����	��Q��y��ϑ(�ol���j
����w������F	��(�Y�~[�OKE�4>Q��R��-%-���JW�N:��$8i1�w��E��=�Й��n��2�4�A�.7əDI�tz�X�R�+٨T���`2�I�X�y<~=�@R��(0z�W��Ħ�3����$���$�5�L�69�Ū��k�R�4^���7�H��;_[�vI��+$�.$U�'L౺��u���2Qc iSɜ�ƢA�m��0�0X��.^l)Q�Hӯߣ��pmu�j"=-�� 9�o�:σ�<��ge��b"�,i�^�M���3�jO��&���f�tXz�vA3H`������w!�bHE�C�TGk^�%{U%��|�r	~ߎ��Gx��;Z.j�L���ۉ#G'�n���x4��XϜ��?��?���o��g�]X֙]V���Ưjf�_�,��H�f�fp�_�/܈������n�}t:� �Si�-��k�Z�w���6�gx?�!�������C�2�+;��lų\;�\� �R"C����5��	��$Ilm�0E�k �Ϛ 8�f���a��g|p�C�v�b�z_��=-� |<���$��]G���$4�����n�`q)FP�Pp �1~f��7�u7��dq�LH�(���w#�;��Y�`���&��-8}�4�f����o<�Ž>'&F���?z�w�Gg�3T� G[p��Qޯ���`pd�}�ݿ?9�u:���=m���%D�!}�e*n����$/��v�_�:&xO��N"�ss$���Jn�pV<��\��ܸ�?��bk/����h#��Оmn�b���W�*���~<���V�����t�;|
.o��� �^���AR��K�00JPrǏ�x��&�G�����o����#W��=��w�����
ڢa��Y�=B8�O�N����|��DVF6�,�2*58<�%vņ7\;)��r��_���F �f22�Z�ͽ����r�w}��J�E���nm��q��c�s��ool�f����G��^2�m!�y��R��)��r�O�ybN�x���~��dx���u��g�ǩ�H���'�`%���f��1<<L`߅͍����9�9t�]��X-�v�M��@�S`��l����2�2픓�@U�2Z:�Pȝ��Q�,����|�-��9�1g#0���<�D:�àKr�\<y
'���~>�*�ٍ2^�a�P�9!�!�һC�A���>P�R���@�������2�V�눓$���zV�����\����Vje�!�8B���I��;G{�7���-\|�y|������A\�zwN��$�%�W�E�d;�m�.�J\]W�ǧv_JN�{���2���Vb�n�$�\���/��hw2�n�M�5����(��n��-`�w��	(P���Kʾ3-E�I��> E+�^>�sjUe��LE%��M)�o"D��3~;�8�����ѧ<�N�<�*څZA+��M�#}�����o:�Sb�'���ޚЗH�3���c�N�I:�p�Z�����>F噖_��]7f\KK�dZ�|�"=����W����)��Oyĸ&E�ir�m'1հb��S��CP���:�fgiGK8s)��B�ص��̰��-��}���I�j�f�)j2��\3b���|^�����\5�g�ͽ?4��mtvuk��۰�zHҢT�a�M��d���DL+�)ѧ5��TS;f����y�~�$�N<Uй�6~)}��JâmY&��w��ͥu�����=�ǈ�3��ѣ�!q���H�wՄ��e�by=���^-����R]�v��{b>H��� cw�uC�� �M����Y?�d�ju�;��"<Y,��Q�`)�<G;��݅��!�����Kɵ�����+��V!1���Zј]T�����IP�L|�;*I��e��T��0I�#?���j)?{����RJG���_o }ݽp��;H&vx_R��������׬Y$9�yG�u����q�V��d�wκ���3�f֌�e��+�q�r���DBj�[�D������~��(�ݭ�����Ņ�UU��C.O�{k!��bk+ɳ*�b�1S��$�vj JX�֬6��,�&��b:������A?R��j���H�M�Ƨ��B��;	 eV�
Qh2)�l�BV�N^�_�fe@�d#ֶ�q��a�Z���F�E%���3as'�}�H� ��n��5��n�dHI}R)�0I�E(����lz�f�yUXt�ZHh0L��c�@�����_�]�������6r^x�3� �����1^��Y��� 5�Y���IǠ��=_+���t*�hj�����Z?�(���Z����\'�o/�&�G��/ҁ�Te�Crz��i��NР�Xm�s�I`�A0��u�#�M�XZ^�S:�����dd4�o�4�Ϋ��D'T2]r�&��ަ�'�*��������胃?�xzk^.QԔ����ۯm��|��G�l'r:�<S�jTD���Q�f�W"iru �8M���D)3�!�b�u�	���B���k���'�.U't�X^���� �x��$�����ڂ�L�Q\{0
�Y���C�?�!��&R�A)Y�
��d��0BTJ��<�.>���;�����;��\�و���#��8v�8"m8�DVZT#U��54rGd	����*j$6:S!����I	�����1�GJ�q��&_�9h|��NT�Ϧ@�^�9pV�U�٤�BT��I:F'�ߧ�T�8��ϧʶ.�D��H~�zN�Z�������������i�7!f�jtI�1ʺHp��gS��=t�!Z�={��?�ξQ�B�� �y�_V����]\�t���ϥ�3���������I`/��e�cGI|�y���t�\S��+�e�F�N����w��ե��<?������)Q�i�����Ȫ�$Wx�vv�^�#�P�%^�["�n�=��tv�~�y{�e�}�c��Ll-Q�s@���]���d��%�"�o&ᶩ#�eH2�)z��	g�q�l�01v7�A���?��N��BHE���W_���!�S��y��|�7���;������A��s�4�^q�}�:v%N�CK4��E�4t>$�MB��$f���r����@+G�b��v~9���8�f��-�_�׿�:.��y��^^�"0�����cue]ˈG��"H�/�Rv6v�$��]���Gh�)�� ��sS6ʝ�o{SBpP� ���F(�^l������'�'xp�C�'�����Ͽ���*I��^��Y�R:���ȉ�<�%��=M��o�#����:���t�&*f�А�	��R�&#�$RUaT¨ ��n�u�3j%"Y��(2���V���\ƾH�P>���zڢ�+=W��~��ξEIy�j/��h�TȔVꅸ����C:V������][��%h��Z�V������w���)��2v��L?���H�LJ{޻��2~)�U?Q-џ��oa���٧�$�_�����IД��"2$���Gl���Xf�
9�0�%�9�f��"�!�����'�O����h���@߀���"��}~V��mC�v�8��
D��.k�=�����������8�/2֨^7��[�;S	C-SGL�R����Uc��delǜۋR��E����q���x殺�KO�����I`m�7��o�(GQ��8�x�������XH$\���7\/����Q "�&�j!�e�W��X��}d�m$wK����h��\�yϜ;�K�O`�dau]�ED�d��,��ӹ�XZYU��II6Є?|�5�I�H��'[�B�${�v����u�2_���gMz����Ұ"�я�v{Q�|�R&����GGp�����5\����s]������C|bՌ�=ݭ��Z����&��J&�[�kiEg���F���ZR&/�KH���rU{��>ϚbȺs�M�A�3�ݿ�6;��'��60�/~��:�V��f�f5k'�T���V�3�{	�I>S�ꦝ��әeܺ��vl��Č~b�tp��r���2����l��R}Q��Z��I���?���v�C�9\%��=\gi�X]F�>J���<�����qLFBf<�K��T�����7�ގ`ȫˤ���>;�_\�1X��dPy�j&�[�q-��������#��9��^��*�JSI]1_A��KE��},�����m'mɷ��Lf�ݤ���-��!�w���A�'Xר.� ��c5��@C49�����f�����a�d���J���\/K*��/c7�4��g����o�o�?��e��n�e%�->�$qu;��CJn%3i�S�C��|UK��v������@oO�v�G�Hα���UxB~U4pv7�H��yߞ*��|�E�9ys�WP���ň9�q�.�ЧT�!͎B!;����JY�`Q��F\�L���-bV���	\~��kg���W��abo	���ư0��ǓS�>��;�=~��x4�@>���N��_��<�+��+Z� '�*���Q�j�`����&�Q1h��X�}I}���|Z"jT *��� �2�V�7��^��D��|о��l`D
�"I��B�;���`��tb��C�u�(�9�N���J����@H� 6 J[)��Ի��E�[�Q�$�$�BfL	��F�b�>)�1�P��`4���>�cI�B�����*��G���¦�@�� �-���j�����5�	�ף�[�K+j�j&J�;y6��؝.b)%9�,a�`F�Tlo���N @�O��%�(��/���G����?��I)��֎��A:L����,/M��2���k�>
#��{��F���l4�6Dn�@���Fx4��7O$w������ z��5�n��3���"�^�HLO7��P%����j�T#����׎/v����w]�64�
�&:t������t����Y�w;���jN���(���x�}^��y�up�?>���C�mo�B�(M�kUE3���7�5Uߨ�=hL*u)�ijS��}A��k�\�A#V0!e�R�)ec�=�jk��:(TJ�Jt��h��؇��n�N�"�����$�u�gZ[�1�9���H��_�A���x0���2�CH�(5+95��%:j����E��4��d&��RјK��H���=�-��'O����]_�n��S3�u��Y�T�,.+I������O�����mʹ�P���y�+BT�Phh9�D�<��LE�F����4͵�"�׬m����8}b_����=Ŀ������?��o�ț���� �I����4$����8v�8��Zqgj�k��/�4"j�A��|�#	:I������r9cC�|] �z��©�'O��lŕ_E�aA.����;����Q)���t�j���<�<F�Oj��;��ŭ�3Hg�hl#��t�i�M	ԙ�F��D�D����3�"AI�@�[3��+�tStx��8r�Y|��O�dqW�i枬�j^{� NT�������/�g��>����V���G�7��ҍ"����'��Xi7��'�׀���I��C��9rR"F�'H$�;���3˒u_WQ�j���x�H�:�(Ϟ�$�|+KHƥ��u|�����h� �.�ُ��/h�8ϑ���<?��:]^�S��%��n!����;q��y:�5l�i�o��ގ������}���q�dOF�|�o����t�[��{||��������$�����X%ȗYhb#��vj&�P�l�M�A�~K�SlX�T� b�a�$�kU��T '_���"U{g��D�L�o�����l�����tvW.]�^C)����ՠ�dUЌiFP2^7n�Fd5N@HR#��Q�vH�_"I�@�f�z��k��(Uf�n�;D{�h�@\�2�q*���	��/������~��w�b7���;wH܇����
b;{$]y,���|�����Z�*j��./	����Kt_�rE��R,h9���ed�o}q��G~�	���<7{���2[(d�H�&x�lJ*\�7A�P�8X�]��z(
[W�u^�U�2$UӲF�dP�K�aTѻ\�ڢ��}�"j֓f:hm�Κ�H�W"���H+"�}�Z����E��v��>z]�-��rZڷB�j���2�;uڞrÌ��Mڟ,�m��.�[��E���P�1$���c��_���.H#)e�Ã����7��և,�����H��I�./"�I�����_ZXо̯~���T|o?ŵ���������b�wSzs�n�����Y�V*�,*���@�YK���}�2��/�m%dsc`�_��?���y���3ܣ�ڨ��U��h�t�U��v�̆f�V6v�G��������qoV�U#���կ���d�J�T��r�F�T$�[��&��WX$!�9�	ֹCx����BtG5��m�b��S%T�Ua ){��C��y��9���,:{G���K;����o5�d����>tu��=��{o�਴�H��$#�l�LO��0�`	b�sb{I��,1�O3Hwn��~���*�d㥪���#|�MLNNcqi��"��M��)���Ɇ�H�`���L^;�S�\��}DLL�'�р����A<'�$�-h�9�Lbva޽��l���"���U�O
�X�����w��������]�h	�����x��n�"Z*�YS\+YD���>�dP��\B��8I����|ܺ��J�.��3g���{�{����sv��c?�#~H ���}t��ً��-�>��Y��>�m��@w�,!n���[�U�#@�#�V�(��Ke���蚈(f�}�cd6wI��ڂ3vh��8J��F�cv��k�̳��O����.X�����A�g��Uul�YD(=Z���=ed����ʺ1�F��+���	a��W�M�X�����zt��18��d����Fp�3���K����_��6g�g�I_&dϮ��U䕵mx�5�Y���>���ǅ���b�M#Y�	<�{�O�
��O�������¡J5���3+�mZ.�v��i�[���Y5[0�b$Tm1E ��n	��A&{��q��/�	��1���]�pE�L�nkӨ�^lWk��bL 3sLH%s�G,F*>����B�!�q�옞#!u���^�(�H6�~0�W?��F�L\L��[)G��������J��4�N2��%,�(�Ul���cN!mR�!e-^�����>������)�8^�$SH�bt��LT��3t ^�Ú1�9-��Kx��Q��0�����������)�ӱ�Kp0'C%뚴h*�(��ZB���4�kd4�l�h܆&ۺ��Ew':�>�������΢��[�����J$P�\�6t��N��E%y%:����̞�r�؇�	ɖ�.i����i�\Z~!3)�=�lS�V�D0��+�����Cw2��LJ�1$���U��E��I��sJpy����"���8t �F�EiPz'��n,��4Id��-�Ice~���^������������{{��MH���8=nTx6��l�(���X�����&?	�;����5�?��@́�|@;���1�A�'�E���!LR�v`o桖:����!��i��G�XZ��r�W������Etw����T(�Rn�|,�m؍����>dH*�����F�L�u#���&��m��t�G�74���74:��eΗL4L�\�<�\>����g_y��?�9����8u����u���>6�71��{���ŋ8r�$jVf��:g3�p}C07�9���`�����I�&Kb*�ڶ�^$�4*W�5���\�p_��7�i�q���k�����7q��Q:`AU;tΑ�~:�a�ĲJ�w�<#~�B����w;˻d��Z�I�G�7)/��ڦp �=�I�<�$��}�s��0�_~�g�ɛ^L>|���|ɬ�L|��m�<��������S�x���M�|t"�#�a�������9���a��Q���$ę�>�l�Iz��p�Dη�w��ժeoo%v�Dg��׍p�O�#w<����l�h��V���嗾�׿�e�=����xB�(�]����Ȗ~�Ͻ�-:1�\���S'�t����;��:II���6F�ae�(��s|x�~�߇�_���������˿Ck(���sȕ���7>1�7^����&0�����.l�T{���#8r���]X�Ki@H���wR.��HMEɺ8m�!��ie��%�V���T�b��)�x�=��S�t�y
�������[��Z$9~ ������-��iՁ�#�ݣJ�3�K�3��iyq�g���:r���a�x�M����J&���0���.����R'x���/B\)�n��N��\�q|�;�Q��XL����s��Nݨ`n~g/<��_{7o=&��L����$����i�3X����?��ͩ��5�����6�	L>}�sgc��!�l/�J�"	m���)l�m�����W�H촳��J��! �s�����p�jf�V%y��k�d%� f����ɤ�\TJ�EXB���!�ͮ��P�'>b�:����gq�ɲ���l��ԙg�$�kT���b����'?F�dZ6q?��)]X���GO�e���65�����th:�>�
�a���	�~Z�m2�NgW�vUPdx`�S����!����Vw��as����&����Źy\�t���%�q~.���il�ƭIܺ��4I��X>��S
�؋������u�2i��XQa%�"�촑��,%�fI���b	����IO��/H����$��x������;|(�M|�����mJ�����x<� �����xf�$�Fo����I�I�״�P2�R�p�T�D�CL5c�d��{��Ml���$x�һ+8Gs�� �ޠb5"��H���c'I/ax���Mm�� ���:��p�o�M�D�(�N�J�j�!ئL;!v����r��=�W���^ڟt�`v֫-L}��f�C!�m����5Ivڥ�%ϝ�����^MϮq��H��ٜ:J�����*��TF�E�+�y�Q"'�B��� ����6zs/�`k�k	K�܇��i�h�h��qX�:���C:�������,���Gfn��a�1M->7}�nI�Hֶj��ZLFE��3�7)*��q�3VUQi�bH��,N5�u�[��������^����]{S�SX]�D�x@2���Z�����/`�����Ǫ]-��o�hshS�5����h4��@��'��D�*Av�h��Q��d������
q�U��d�aaq�Dq��RS	��z�>�>r��� �o�۷>�Y����׭��[}2�#�'��p�*2��x�w�-T��2tE\$���	�Jh#y^۲��� ˫�Z�S��=z����M>�q�ݸ�2�W��:D?�6���:��|�x]��4��9T��̽�$����9�Ox�2����̳�!@�e{=�R�%7�aB��B"K2��H����s)ܒH*�DI$�Ӥ���į�b~n�F���eiq�]a�(&-|�CkߗW���g$�q��`�w����Ӛ�}u�� S!%R6'����=wنfSJ"�o�)�ݍ��;Z��O�G@t��}<��t"GB`�	˥$����o�����h��&A�4H���'%a��R�e�Hfr�F�p��Z�*��0�0?���c��u?a�oޛ!�N��	�{B���"D�&����~��ѐ�5�{���<�~�T�$%���3X�g�d�$��Q��5����8M�X:ǡC�=�V�i#! �t����$�$��|ϏtO��p]?��� ֽXBK_�$:c�V�ˉ#th����0�	�!<7"_, Jj�e���jIR��2����Ԗr%���٩Q�Z�Br�LP�k�HT��tR���RA�I�4r��Ew��U�vS<���D�NH$FjR�#�v5dE�$.����!��������^/��.un�=��i	���{�_^�c����)-A.5��%��86�{چ��y/�K)���C�$�!��Jc����[�F�L���j<��[Jl�|"t!)~5�,�DgO+�ұlN���ocu}�������I�2�ah���8���M }�$�f�]���}U�"�\!P��=2��Qs]�kY���5�ʛ�f%�9��Hg��ݏ@w��bm3N���ǁ�=8�<��Ch!��R�۷���4ZA��=ܹ� K4~U:��.>�a:�YJ`[��>�h������
�.�N%�.�Gm������tk����M����W�C��9��Po;N?{�����΢�_K��<�y�Q-������4��<ׅ�y`l��ċ,_'B��O�(϶X�趔�J���]�E
ۥ��,�,�ini�S#x�3������T K3�vx�z����;W�~���\����$W�KG�Q��$7vg �|�&~��k�L�5zGN=K[�����@0�[t�$�,7RŐ&���2�Hs�� ������o���Ο>�����C�(��=WW�&T4�'�%�>��:&)���/�/��n�$���m�üGRN�U��f�Nܐ�l��:l�7�G�#��7��w�ҥ	��	�7����UX�=����,
��!_���7�8~�e\�r	�GFU<I��]t�GO���7����8u�溘��&	�ͦB$�OF�����kߠэs��ǧ��K����p�s`�+Ӵ�I��5t\Q�P@�@\�:nݾ���4�w�NO#J$�C�p��$
5;q�I�w���W�k&�K�8L*�UB �\��1�(
�ZQ-�b��XY���N�]A��w�?���G��>��W��%��{�[;���Y��7�E��3'��{�*Tt��C�Ϣ7	HEI���<�e��b^+7�\ۦX���L�@��$ahEO� V������.|��c��c�L��~=$R�ۋc���\uwu�*mW��obgOiS��JJ�S�kR���Ӌv�V��8�r�\;�7��*v]�"�K�q� ى�� [@����A+	�ѳ��:����L�8~�̣�-�W^����O�P����O1��z/�xEV���W���ױ�*Ӟ�ۊ��f;�����(q���%�+i�Z+����R���⳺�ϔP��q��i�nnbeu�!7����Dy��7��?���I����Dp��� ǉ�DJ�F������}�-,�� Yh���бSh��
�z�h��Q.RudKeQ�Y�$�*)y�>����:�>�ߤ�?I�l�����aFZ���;� }Y:S���G;�E_���A[�E?1G���I޿��	�=�Y�q3�S2�r�įI��̋lj/vC���L8eD}R�w;H���%ɴGI�XXIh���|+��h�6xf��DpЁ3�!�D� ~ai]G�s�v�s<�n��F��J���T�Y��c�{X���I֫XΫ�]ww7&&ƹm�X��Ո�n���isΜ��#������[z�����h�3�=sW�~�%��rSE�|�v����h��X2qms�7�@���W����L�0"�f����Ȣ3jG'�^6����[QMӟxE�>*@�whl���R/�|f��#pMo�h�g�Uḇ���qJ9��-��R����rI��Ș,���14F�^I�4�(�����&�����nޞA?���3�ܟK��_��vL����/�3ϿD�|�k��Teu��d	[I�q�g�s��3G��m�B��`�������d6��d�ҥ8f����_]z��p�*\v��ǘ����5kY���jgw^gk+;Z�j���SZ\<_^w�6��`�V��G[5�])64�,ju� �s��(�T$(J�R�.o�цYql��g�y$�c��z�6R��g�w��h?�����f�Clɼd٥u�U��с�!L��YQ��d��E�>('�į%��_�Ц~vC�W��J&�i�=~2oP��eΙ��5�5CMH�fd��(��/�G,ڛ��K���3g���F���%��yn�S�LO����Y��,�.�cw{����F�?j��n���B0ԯ��bɤfO������t�+E$�9�;�2����%x˔iY��ׇ��M<�y��U�V/?C�>�y+NzQ�i�U���t��D���Í��IW:��#ܔ 2�0��U@C!�vbD=d�`A��=����"N��cz D��C�LI�i2�/]	�T�Fx&���GI&��z�'�ؕ�-�(ZzG�pIIQI}E.�5�?�t��FF������_/z����"1�93��)S�U��*��ia�r%�̐ϑ��'s(@9=�Ǐ���������|����ƦF�A /ٷd:I �5�s2���V�J�f[K .��Y��yy�>�����-:�Ӱ{�H��!��� _��5k���Ӆ�'�4�&� �4�D�D��@=Z��r҅�-~�:�UR9�k����	 �gx�+M$?!��4��H����[Wq��M�[��9b�t8}!E"D�L'��5�ӯ%�R"� *�Ū��럒A�+�¥��&��Xun�E��[��8����p�ݟ��?�%���i��hY�^����8}�8z{:T���҆���_s�Ӵ):�:� R|�*?{�N�AB���t�*�aFɈn�.I3h9_��m����{5+p��|����%'��R�}Z�r��#ܹ��$g�xt���s�\�?�g�[tܳ++t�#�9�����k?���/j�0�s4�R�%#m�v%�U�B�}�ɼ(�B��S��ޣ�1��X]�VuQ���F�Ӊ�x'&�11ԉ ���L9x�a?�E�@�MC���m��`FK2r�N_��!�Q�K�@CC���J?�
��, ŵl:��-�*͆����/�<�8޹~/��g�h������2~y���/��sW�p�·����`re�O���(m@�0>����sb~uK%t���o|�gË���hF�MЬBVN�UYˁ�n�LS�xxCR��W�z[{��?�r��U��o}�5F�e�_��$��4O�㽮9�`z	U��>�[�K�˷���j��\��h��F%K���p��A̕�1�H�.�˩�VO���p�ŗ��{�����>�Ug�܅Ӹ�����03����ܼ�C�Oaze�kk\�#����y��a�X�|�@�wQK--6�M�a-��.���G�����a���k��Y�N~��D5+��s�]��{���il/�px(��o�R���O~�����⚶?�:s��_�K$��q�?��������Ρq�����M2C�vB��D����rV39҂ _�\��s�-�?���]x�D�	�y����y|��������>wt`o��X"��4[�I`:����/����]<�Z��y�V���FoAg_�!L��8��L�
L
j*:緦k*�Z���\��xb�H��}+��^Ɵ��E��1Ν:�H4��~:����_�ڵkH��E���^UU�|��?��b�N����}���ȡZ^��dUA���_D�H�
=.'ϔK������9v-#�(ME�9�ӆ��#<	�?Aw0��f�~�����C|����3$��y�ۉM��-�Y\���5G�jqEP����V�" �s��y�]X��W�u�����Oi9��T��]^���<Kr~�7��lq�/B!a��Nm��X_����q��m,le��� ��Ǐ�A��#I:t��<s�H;�BI��Rޫ��V��S�mr?��b���C��>!H]�3��di'�Ƴ/��}⦶p'��I��&�w����_���{%d�-�U�<�<�{���6$�;�s�:����Ⱦɝ05A'��*���**'�Bj*JX�̞���zې%����Im���&��<�����%ĶWP7�VA��������l���d�������#|]������*���0�0���C9R��Il��QU%�Ү��OT�ͧ��z{w�d�g7��_����7-V���{s�k(��ߎ�����1��*D4Й�����V�Ň6��C%�nb�*mY,SĽ�y�Ώ#�R+hO��#��^��ŉ3�FR�����S+��{$���<gØ�Oj�����GxFu�HY���Op��#\�B(
���ZNu�BO*�ʢQu�Ќ����y�ϝQ���{�@L�B��S2����>E�ߟ��*<������y�����	Leg��w����!CkwJ�����p��j �+s�@;C�XR�O�W��ϗ �/�:?�lUݐ�g�au�d���dz����fnv����c*D�K��
��j%~��O$�]�=����=-�f��DH�C8����a2�=��V4�	��<vxw{�B���|8��u-͵�|Ȑ���~K�z����R��B��Gz����RW���u�FuY��GFɔ�
JU����F]�!+r�e��1%���j�1U2$cDHd��&1~�Z5�,��-��Y�a�R��+{���dۛ	I�	u�*����FWw?��D'ju� zcAUE�@�R$;^���a^�,�k��>JgdC�@B2+փ��
 Q���i�?H������F��� �a�
�d���[�*t�����|�t��obz�)���N�^�gH:�M����ar�V�k�@�����$�ј�x��zz��ׇ]�Ƚ��\EZ��^B�	���+��d:�4�޻�G������ё1�xP�Ö�,/�#��"CC��j��s �K��̴�2��Ը۬F�RS��A(�ZlM��ZhX�K�H��� ��Kh���||w��\'��"jE�nŭ;5�*����]8�w.��h%�W)�F��-A��)r��ͫ"�C2K"�!3�"Q�n�w�Qji����^\���~�ͯU�9q
�/>�K�?��o#�(�߉m��q��a�����bq��#7	t��!.�]3�2���0���ҿhsZy�*�M������#�lΣ$��vv^ވ߉f�ik�_���/�B�ԡ������I-a/��,4�Y)c��$8]O�`�v�kx�Gա�6��ש$����A�0��Dm��SoȦ��b��FF�NJm�	���5����K 6���Ho5�1@����In��oQ��o����)I��s��?8��D7�ro��.��cϠ����SQ��2>����hdZV$�&R:�NK�z�������0��O���{5��,�k��8�"��4?��/㷿�~��.����	���<��`��x�կ𞍪�eHf�����������9i[�z	B��pv��o|�#Y_��iJD�ĳ�{i����A�N��m�^%�x�W�B2*�xu+���5��tU�����ǎk�G,���xXdn����y/D���ؤ,W�jJ����H2����Wz,zw�Jx��S���㙗~�|��ɻ����'<{�$Ν9��9v�� �]ھ��n̤���$b�	,�niڡ�����q��n$�`=� ��BRbQ!,�	(��V)h)v;m�����8�BZ\�U�/�
+����w����=���k8�1��cg�������N�jDU�?�������s��6*$;<�"I.$"��k�_z��)�Le�*i.b*B�¡N�kY��Q���|�Oq��?ţ�Y���`f%�S���˿����r�����~p�h�?� ҆����T} ��]A�����2AZ���MU��$2S,[L�����:��Y-�@�Y���#K_e�z�V��f2���|�Ò��ë?��ˋ��|�m<�=��$����������������m�~��?킯�|�Cى���=\��-��a�?|�;�!����PY�Y�U�Ţ��2�B�/Ɍ�K���������wn⏾�%<s���j�S�����[��mG~;+q7�S�`������ѧl�	�7h�
�����������a��`+}��j���i���&�?�C چ��8�H�cc�~t������^͕�W��>�\o��2�}eyG];�=3mbB3z҃�С?�'E(B/3!)��VO���m��5�b˻�������h��)��r�{����k���?��G����w�����g���}b%��瞻f����7������ߴ��O�����;��-��q��1K6:�[uJ�<�g0�*j�|{�К�2��P��5.�*h�^�z��s┈�3O���?�د�xv�N��Uٍ֟[w���[�{ު�����g�}bO�ص�/��h��}a���������F��CKm��>o�Ͻ�R�5�'R�x��J��hܔ'���AU���4&��=�F�������G�ٿ���VF`W?����͖u�	��lm_c�H�٫�W����r���+o�+���e����?�ǽb�Q)����A�5؃v�#��^��aS��\�=����~`?��mtS�"����q[9qAJ����nn<�������������+N۹Kg�"��d~Dl���:�Iv}��@l�Y1L9R+O�"��Ƈh0r��I_I���TK����:,oYn�3����W�%x`�^�����׈�xX�{?��c���B`�<MѠl��y�p��=7��ǨR38�/-6N��<��eDs-W���|�&$�W��]��U��>�uWc���v����63�bDɟ|q���얭�l�PA�̩3v��6�x\b@��f��9�\#$��)c��c�
#6{�[޴��x�����!��){�U�S�匏1`���ɔUt={�!u�<������/޹aɑ%[>s�fOCO[�Y���kϨ��w�&"��A�L�è��¬
*�8c>)���c�
,���;e�O�؍��v�ԜeKfT?�G����ʣg���}��C:?��}ۢ�*�PT^X8i�O ��e���$#����PH@�c�)h)q0���=ܩ�l�=�{�<;a��t͎���o��ݺ��-;f/��������U9�{[�dk�z���36:7g�3�6�0cS�;�l�	qzT�'͹�3�IY,�HnȆ`3��-�M;�{�V҅����q������R��v� ���;�� m�ߊ=}V��y���%�6,��W����+���0x�H���D���^���$�	�.�T����l��j�����˜2�f鳯���ߨt��[6�u~�6>����z�p�7�)D�����~h�O�ٻ?����_����� س:�����4�M�����7��DZd��>K�	�"��j�Y*N� �Mb!Wm��;�A��\�1b�t��ܽi'�q��o���_����So�Di�zK!Ҿ��0�K�N�v���;O-5vLU�d���4𡴫�j�	`��:X�E|���W����l�� ^OUM��"Q�|y��AR��=s�~�w%{�W�Z��8�n�4 ��ի��mT$����[Ł�!B`�&�"��䴋2�;)`	� p'������G��i����g֭Te�wvk69ֆC(e,S���1�˖Do����7�c�������~�<۳������?�Ⱥɂ�/��x	�/�r(��؇�B ��ţ00�A*�UKAM����zWt��ZǦN*���V�9�t��M��sh�S������f'��7���}�ۯ����y۫�-]8���2D���YE���C*�M���/������{�sx�~����g�� �P����^�|k3��l�_���@	��N�3
Rڥ��.�D0�'�#� P�_��)Tdo��̾����d=]BW���gs7�)" ��*��"9���P���6TLۅ�@�[���C߰��J~�[�yî _��M��< ������{`K^���sp�ܡT@���ؿ�"�x�Z��SrT����I{�������i&�	gg��V����G�C{�Woۧ}d_x͚0o}y�>��=�,�N�o�[�M��cx�c�͇3o�8wӇ�5�MN���5ša����[8 M�o��O������5܉u2����s�4����G�6�^���\��N��H'����}�`v˞n7 6����6�|R��Hub�-�3�M����O�Y,&�ً�C��l}eRE[��1ӌ���՝]�<�ѡ��޿�c���b_}�k�������v��q[:��cٱ18���!����g�ٯ_�E�?3�[� Ga��^%�ù�]f(��OK�Gf�Y���8�@�c���{���c���}�'��_~l�~��c6�;G�Z�g`EhNtA��;�y}�����՗���tc듰B�diΧ⌹��� D�E�C�-�� �s
�-������-8�%��?��)����������ݱ�Cv��j����zt��o��&WN�G�ۇ��[qd�R�Y�)����֩w$\B`EБ�-9�J�g��p�3�#e��*��qm���������M�(�֧_����_�]������J��_�X�Q;�/S36�3��F���_��K+#X�2%���7l��9U2��Ф �r���n�UKHo�n��Tl~iʾ�{d������Oޱ��W�_�џYu��v����\��=�)����,'��&���l5|�~�	��7�4�J��ɳօ�iPtg�����k��K�Ɩ�l:{S�{�؄{���}���ͳ'�Yir�����ō[���vg���k����$@�ړ'��ɚ-�<i/����O��]���g�$l~ �K�;�0�~X�VS]�J��Q'f�D����>v$��c�6�u	�<�k����O ��w�����/�ַ7��$�:�zV��z�]���z�����|����	��f��o|�^y�{��b/S�>P2(��K��sNI��r�9`�N�-�A;@�O�ә�^�z���-��]�#��߳ �������w-?zx�z���o���M�5����������� �J�+XH�9)
����	�1����Z*�2hu3�=����{�!�����wn�Ww6��҄�����O����>6�P��([fx�Nc�N���s�{@��G���	4��>�sj:�'���5`�O��$�:Bq�TBX4�akB��J�J�>[���oX-lٽ���޵�q`��8ޱ'A�u`�;��mك;O��9{�2|�U�����
 ��a��ɢ�(�\�B�����q�y�2��V�j���7n|�}߷��|Q�V�\�V��������[���Z�>��ݹ�w�j$������ߵ��]��Y��,�rC�ݼ���Gh|�����('�7s�UF|l�}�؆3�9���'G������i�����~lO�a�N��&�������{�߷�g��MF�k��`;������>s�~\V
R�N�XR��Y���@����6��//�cc�8#��?�Z�.��y�l����X1?n{��́�֏֘�y`k�����MN���	�����l8�3��^λfH�jc� T5��J�kų�Ӻ��8�A�d��k�&�K8gbf�~�'j��o���lX��m���m���=�Ӛ��G2�K6s��-�Rs�&9�x���Q��LS��I����!u��D7��GzM)�'���h�Ɨ���t�=.w�ޝ���ͧ8�;v߿� �E��c�v���z�*��	m� ~.$t^�R�M��$�W��H��f?%}[�n?��=�NE���S��xx��5����&3cj.J�} �@���z6�6�#X+k��u�3U�٩a��T���g,@�ό����=�uN�6qr���a��޵/�j6�zղ�sVa��Hp��D/А���[&�������჻5�%�?0l$1c�F@��7��&�V��?��J/���mK{ �36� ��՗R�+ײ�p��,� v
O��sA.!'����a�f:�6��bg�{����T��!�g�!+����l������;���!H3/'Y�j��rh�;-;��>u�wF3qʕ����-�+��%�L1'���iVV_�Ι):�1�ML� ���U�`����{`�yI/Ϗ�%�'e�!��^���|ϖΝ��W^�-^��˻��Ѧ�A��ֶ�ؙ�vlfقܰu�2�9 �<���E�r�tV�1 ��c ���mW��^�pm�2���T���+[x�=\�3��xQ��,J39�s�B@��uط�<��,�H��x/R ��<;.~ΙԌ�ʾm�men�^~�{�:صOn?�u{�V�a�\��� ����GR�d0��s119�* e�}㐶��O��*�Nr�yII�����%�\�{�5I����ܟ�����T��[��ר�S��r��Ol��s7o=��ȕk�mt~U�%����?�Ԋp9�w���n޾o_�� ���h� �S�7���}V(��'[ {���x��oz)�Ί��Ρ�89io S���Ϩ�yGA���3v��I[]^��[ �{뇢R���;���&�1�11�@lǪ���'���K/Jmkk�&����7s��l�_�!*ki���o��J+����������gO =��\�x�N,� ��d�j���^��p���B@z�Yٞ������^��M.���p#O��֚U	�����������0s� 1�P��	�����e�I+�=)$T*d����xÖ��ͯ4D�\�۳o# �$oQ¤�tt���I��J 4����Ğ}�K�� ^x��`��R����}C��1@�����aF�h����v�����G���KĬI��s� l���aמ{�ff��ރ={�s��#��b�i&e� ,�g��/�2�Q���`ICd�q|r�^}�[v�䪭=~`�~��� s�:lI��܄���ݸ�k����w�iq�׼eq�͞����q�4w���1���[��+�Q��1cR�{BD�}��8��:{cv���a;a۰;'�_��偽�ˏl��5�awpF�������̂e�v��{�}iOH�=f�������e��p�֢�T
�)f�_9犙[>7{C8�'��(}!�v�e_|���[�� @���޲��O٭O~e����@�V�v�G�3Ӳ03�ܷ��������pl�.^{ݮ������.11�⼹��.Lt�C(������ѣu[==ko��]����OoY�ܰ��/����k�߰�� �u{�x�|��,@J>Ù�E;��ݻO*R��\��o����� ��x�\μ��ks@]��T&Ś�+���C7�ԾdRI����`���䇕b�_��������[��;��/>�H৙$ 0��l���]y�Km$1f���{���^�;y�9�|�o��El��a��省�s�U&��!#�Ps����=����Z�bƷ��5�#`����qo��'�Ώ�W���(�˳��>waզf�������#��3��I�#Tླ_��v��X����8�$�E=bV���9[X\����wlwo�������|/��,�z���*w_��6���gI&�x��*�O�������0���Jw�	+iʘ�ύC�7;��XlT �I=�K{<\��)  �۰���������f���Z�}q����FKSvqa�V���,��(iG*�$Ē�� � ��XM��&Ai�)�Ȇ"��~k���H�l��ؗͶ!�~:|��>��M{�����Bq̖/��xә��Dk����\ ��$Ģ�Y%Z:�W�g��A�e�엑)+���zj�+[VȆ�0=���i����9ڱ��u��Ï�Ν����|�`��M۵W�k/�Ί򤒞�ZGE�d2���b�t�B�Z�'��,�t�"
��]88�a->}��vHQ���GgaO�d�nc�#�x|��ǆ�þ��/!��gX�5�u��	5�n9`RXO�� 5��a�#��nG*&1}�J�-G����L�2�Ĺ��dvq��x��ʎݸ_����,���������w����۷�>S2�8�`�V/�깫8��b��9kr��u���Lv�[��U��5D�f����C�jv1.��~ӞnmY��g;;n�a�p�"����Q��z��8"c��4:�\ �=�����X�NmP��*a�ǀ��D1Y����k4aG��G��1-�(���2�a���w��H�2 �l�����[)7dS�ê�mDl�ڳ�D&M1*m-���F�b�p�g��G�f_ ��q����%�`(���'3�}���I��U��x�d�;�:
R�#���⌹~�������Wݶ����a�m����6
�Cё3}��bEmtB3��p�;Ъ�Z���}|뎭�\E�tقt���CQ�X�s��U�P�U9|�����i���+��Y�O��'{��m����V���Ɓz7�������lbfC�K���L2�p��p����W�a@X��l��: ��o�f��~4���}�Q��R��@0	�w��Kk_|d;0
� =��:w���������اg�dl8�⃛k l�  �F��֡"8�=i�{�>�q�FU���*��֤e,���$q!8�� 0�@jŢn��.��)��}�n�\�����ܲ��#0�K���o^�B�*� �_�޶��]{�����ؕް��9�ꌄFLjx���T�E��|6�WE�t�����+���������g�ڇv���v���u+��s�w���c�;?����MLN!��k��~�0m3��qi�Ì3#�L�_<=�j��HD�jGe{�xY��囙� d9X��P��tNB&lBOa�.>����?|�������O��  ~F�L�� =j7�lỚJ
ܺu[J��E	�ʰG�����4	�TV�=Tl%3��y_%��K{����m��������4���#�^�M��w�����s��ہ����4|w��;��ŕ�[>#��2ޏY-�F�J���uS�0���qK&�~�m��;�07i�/��q�z�g�v�����ش��M �!���P�����M��a���6� ��*���Hg���W�)�H�����}G�J ���PIi�=A�f�r#�P�+�<=���O&��@����}��]��������Uh��iJ�k4C��(��F�,�mF�ۧ�N�a���s��KE��uM��v���p^�rU�d�-����l3�܌=��R��Zw4��v�3�x��\�V����FWp��Ĕ�)
t����L��贬]�i|�A�bI��E�$�S�Z���} J�Y�ř������"�]Z�����PV��i�� |(���[֨��v,����]��)]�% �׳u���=u�׀l7.��;�^K�N�=@ 1=E�J�����;Aq���/�O;�/�����;������kZ��������/x��&/<o�^zÞ���=H�>c2&�����!+Ұ��/$���,>��l�+��f�ӳ��Ol���k;�2k��Gv��e;ur�*��i�Ӷ���mԞ�ͻO���u� 6�<~��_y��_��Ә�Z8�I ���)/R ZlǢ��K�_{�k��&�������;������Ϟ^�ܰ��	�Olc퉽�B�~�`|����g?�_����/�+o���_{g��;u ��b�W-�/.4���T����{�R8~�˴�=Q �H/��A�3OS�����i{�ͷltjVJ���[0kc]7�������e�=o���|��g�������'��e�ã���I���KU��u�$�������>>���E�_�)" ���F9;��s� w�P��ٕq+�s6��شl �uH]�<P��e�þ��rm?}�%]���Ja��� �v
O
���� �S�.Xufު������.�Kq��C#�%<9;����#���x^+�i|6������O�<&�l�����Lfqؼ��ci~��b���?�0��J�|a��$���>��m͊� $C#�����q�)WO������3!ƣ�����H[��-騘<3j�a?1���@��@	d�˓��'V/�� �l{o��=���y ��}��5*��&���%[Y=mS��HLc���AqUL�Ji�s�����1{d���� 6���cQ�l���i���!�5I����S�#��6�����:|G�̳��E�z�]����1ظ��������yŤf�$���X��W0���k���@�I�0V��":�<�wl���Q�G��>ܲ֍=�_�r�y<wM���a�6��lkm�*�g2��+�p��%����%�G�>r,Fw]�V�QPIF��쑡�R6�&f����9�SE����p�v6���D�=�:�Z6U�ٙ���I`ϳ��zN#d2'I��Q��I�Il�S���}l��Lٙ,�Y%(���[��trX�Z��~��Ow�m���΂I�ӳ��q_X�E�K+�U��PI��vm{dB�	=R��*8Dq*�����������2������Fu?�b�mO�@��b�� ��1L$r��fǦ��ŗ^��q9�ܐ�����M/��|���ێ�W��@�kdɆ2e&n?��gUmf鬝8���3����B��x�	�25�"�+��p`��^�j�����(_����y��M=��x���! �} �5JncA�m�퐙�Q~��2=\ߵ�Z������Y��_�X� ��CG	߈=��ni�:8��[���,O۫��=U��~��~�����K����-��m�{���>s j��=�G����l(�<{�9;��([���"���Ѯ��و�D��5���Q�(rͤ��=�Ԥǀ���lpx`��m�S�4���9�W�������v ��ИM�D.����mc���珟W���)$��Aj�L(b1�D�{r����J�a˳#v��e������q�v6H>��:��S:��bN�FJC�\Y��}��d;��1;}�%��
�Rp���}@:Ϸ�`�������Z�Y�!@Є�=}�E����wm���	C���-�\��/aߊʲ��a+��"���&@Ηw���c�r�.���`f ��lz4����L��1�fS�"T���UC�q��a�r/��82n���{�n�pxӋ��&�r��U)r����_Y�ƹ�
3|98����vl�M��9*�6!|'+O%^1����k�JH�8��pA���0�:d�Omgcvn��\y�&f�	�?��߿�3^,|�=+�Ɛ!�&c�c��i9,%8
��	\f�%\��1cK�`:JR��xaP�@�C�wRĞn�KY���i������g��;?��' �͊l�ҥMI����av�ߵKϿa{�lW,SLYS����&P�+xv)��x���@)99�(��*���f�C'���f��1��E8����cU׬�@��#���᱾_S�L���8SջSmO�&��=��4�(*�� �j�^�NP��"bVN>�jF�Iȡ�ꡕa�j��H��іqv�E��-D�fV {�m�{k�{弋�b�k	?�V92�Y*��?�L ��+Lw�~�$TU��nH8�f���:����͎�Yj�'�˪.3:�Q �TBAI�e,�U�j1׾/�¤Î�r�#�mv8eø#����0��=�>�N�8`O��n��M��A�okO6l��V��Ƿ7��K�?��ϕf5�������m
����K����61������
N�L.���~��fo�2@��{w�����.�,eL}��6� ��_�鼽�ۻ�c;O���nZ~ҷ�g ��-������>�ge`��U���u[>yѦ新�y[ۮ��ˊ�8l�o%͏tgf�Ն�=!)�=����g8�;fپ��?���9���O����Ǟf�������߆{P��>��vD/?c����۱�+���D�]�`j�p�D(�K���4>0�=h��2y��Kk��p)0��� 0!g�����-��)u�lf�T���^�>��p�*k)�e�����s��1(UF��E�Ĺ��V2�Xͤ�o6a1h��Y`�+r	I<�|	���)�#�X�	{��?t�>+��t���@�b8� ��@�
.�8*P8��ﬔ��3)���
��� (� ?��V@"E��1��E����M�d�7�W�'v�������|�D�
Xh�S"�tB���1�+�N��*���6/�]�)�
q�Hxc/;����|��̲����օ]',d�� *-<��d��T~W@�����dtIl�HW����+��!�%�Y�V'C��$0���V����#�_*;?��=��I������ވD�F��`�"�˺5Y}GS�2T /�^���v�E|��@�A\�5��E��I��#ӓ�1{�t�1���yo�B�9�<��Sv���-,.[id띵�jK=�����ɹ���٬���p����3;b4��S	��q�ɸ��79������Nq�I�H�Z�F��-���З�?\����1��E%Fǧ�4<�w-��z
�
�U�RU,��s#���D	���Q���a<�i?pUt�c<_�/Z��`��y��Y.(�������Fq&�{�����aR��f�� -4׺�)��$&Ĩ̺�
A�-�W(�X�X�&�g����A�)'Îp�ci�d�S�VW�W��mj��R���������F�/.�$�o�G���W0� �`T����:��VOJ�T��A��1��,�|�(!�������ܵ�ʒ]�zE���K`O߰_��	�q{��e����+�8ұ%[��S����e�2vzi�&�����Z�iPw&�j�'	��r<�	gc����b�/EF�;� %�����]_��^��8���,n��P-@�1iM��W�2���r�609�|�k� gm7K�0�5 
cI�T�e��o�é��K�ڷ��1g���mb��߲m�T+���G<8����n�����an�l��6{�9[<{�ңs�[����yO앣�ʥ.����ų��]�,3/�b}��ƶ�`% ���EK�{�������𼵑!Q2ַl��LYq�������wm�3sѷ��eU�F�7:���i��� =�N���`4����./gM��q���]��wĻܸ��ݍ{�_��W_=����^������_�_�K��C{�g�,/���u+M.�A�(��E���9N@(u���
ST���e���z�>~Z�F�c��N�v��M{���W޴�{���s٢��E��=`���-S�.���j(�F��9��醢`1ۯ��I�v�ř&:f#kp�b^����l��*� �k϶��9>>j箾 s�>x�y�̶�f (9t�B��:�dV�6i�칥�F����N����2 (�oPU�ad%�	�GŬ,ĥ�q����30�Ż�8�Μ�j�J�6מh�uϑ+��$_�ll>���v}G�d�O��DZ�j:� *� K��H`��0��6x"³������QK�Ӷ�y�n�sSv���vr�4���G �~�z2o���R������/Zh ��VY�-R8��bډk!G�mSe.R��t_3�|U���D	�w]ҁc7r��qꌔh����:�=�BQ�X9 ��!hl7B��t:���Uf��"F$M�N���o��L����+p��V�Y�$
���^���d��� u�0�p76PD�$ٷ�
���l}@t`ss�8�3�'�r��~2��W���I��.���|�|�OR��LV2�dQ�C�>Pڥ6�F_4�1�Z�f-��>��nP<9�Z�{�hg8�7 ����p��0R�c�,,�@pd��#����u�Y��t?�5q���|R�&&.�)$�(�5��. )��8;o�Οh.�'w��q�*��[[��/��sg.��  ��v�T��B�JT)�j ���Yx�|��P�O��3�{�z���<`5�ە��������/�l�|�|ڈ��@�[�l���J[��d��%��o;�z�F'�P��3�]������>�^����J@����/_ XHGI��ɉi��s���ß=��v|��}���������uj�y*��4��5#���n �\���Z���c�W�X�Ƥ�6�;�\Ӗ�qV�VG�EV��̉T8@3�����2M�̈� ���`�io����W�ށw���'�����ԲDI�c���A��y��H�P�q�X~�=h��
�'���W^��ѣ�~�I˻�¹`�GY�DN	� ;��F��T�{�E` ���Ŏ��v��^/�}/��;|6�M��1�g+|ܥ�W�20����6m�4�����1$�.)��.�g=�̿����g)	2�����k��;�k���m�J\+�1Y\�>��5�	��n8e��A�(p �s6Cͽ��P���4������Y�w��p/Sz� �j�V��p+nwJ��IґDG2�ر������6�k�}&.(R�kp�)�J�^7;�c��l2;�JEI��Nj�KF����w��]��923�,1�^7V��8�=%���[7�)�W˳:���;mCCv|%/z`����T �x�<�r�N\+b����!�8�`�;P��3����Rr��4�H�I?<'�qX�Q5Ø9�(���j5p�lx"��@~� [�DⰨ�T��grbA���M'#��}���>�"q�@��SP��b;K���|Vχ-½��w������x�P>(��:2� U��\X��S��#�K
�p|4��&���O�@I���{��=B��l.�q"
LaS��"ˉXo��+j%b�a�x�,b��$�drJKǤ��&Ld�5�>RA��Y��,���i��}G����1AE�ۢ�0D��2���kt��8��v����ƏG��iT3�܀GR���!k�ͻ�;1g��]�S��>��}�����Olc���X�ֲ��lrZ�C��a\��V�8:�,�ak �,�\���,�3�c�I�,)�:rO�ƎN����8oϽ�"����ܳO�nٙS�$||�����- {��aq�[�q������)��:����r�� Rb=��g���L�����0<iy;hn>شّ	���V��A��Ȟܻkw�l�C���c�K����ϙw���^:�5Y�:�>.B�=���]�.8�4l46��l	�gfO�9Hp�	*��hV�Jep������c%����5')Wi�3����'�����d��U�mfjޖV�{T��-��āW������T�ՕT��D=`�0��q��2�Ŵ�<u٦f�?��k�m{� ~��=8�=Q����6�@G�6����,;r���,x'�3 V]?��"bu���܌&8� �T���hC"+s�v���0��O(>�b�}�g��0�F�\���({����:x�����K���_���,س�!�
`ϱ�d𕆁#K�x΀F�'�eV7��;ƙ�;��َ��(`01�b�+g���=u��������HQ�3���j�(m�܍�O�F����h&	4��K��	Du�w�ML��MqҐ����%�*�ͫؗ�r`E�Y�C����.�B��(5GC�ߣ�F]���@�{Wzx�����X
�2!������]��;�w�a�&�l��[�l�vP����0T�5N��h	��K626a��@w̉�t��Ṗ��X��S��Tz�$R�S�4sʅ�p���t��G `�xת-%�D����Fq�[�Vs�|���]:3�	�,h&eZT4���&pII)j85{�X��-VM�T��$�l��H{�_Y9��9fr�'�ܷLA�|N����r�P^��M��<w��:��֟m�8��a������J
�Z����eU�a�7<LA&��v�d����l"�@�4 �i3I���w�*p���9���}�N��j6���:T���C���T�����%"a����}Qo���"6�M�E�b���i5�1E��{s��"9g�{CUk�PR�藆9���v�Zv���zj���g��B�5yLt�v��ρ�<1���'{�|՚=�Gtp_5�#W�́�z��wm����i���� ���h�b��'��|�[9���O�[�3�z	��:����ĢXy*���j�7H|�:
B�h�<Ҡ�1z �ҙe��gjck�Z�Ź1{�7��ً8��؃�5�fqW���!gÆ�W&�h��lm[�`xtʊ ����qO�%|=���^�n̶�j�3C��A�
��̥�l:_��st,�τI�1���6��8�Dg.��bD{��*�� ��-{����Uq�8��Cƻ�j���Q��0:��{�X)�����jW��+�J�D����H����DM� |�>l*P�=�0��}�@|� Qt�PH�m|Ld�d3Gud�'[ם8Ğ��I@�k��
\�����.R��8-�6��x��b�D2'�n�s�$�OP	��9Z�N�D#�VGJí�c�X̒QO�lf*��v0A�PmKL����wged �ǻR�}t���?�CV��L4�_Vy�)���ه'WO��҂|2�=�`ONNȆs�_"�ջX�{D��#j t�5�c1���5�a��_��(�L�j��� �CLl����g�Ϭ�B諺Աɑ1�op%��)���R�zј`h��d��J4�nixF!71"��D�Ԉ1�}�)���w�Q�oƑV|V���I�/Uvi+�
t5�-$Q�X�T�V0�i���"s=�db�ļ\c�5���J��L$�A��������$�DSU��:�`^���:�[��=�4k/����H���^�'H��<��M�Ԭ���<���}�޳DW�вT�\�7�I�EC���8[wxg�NLzƶ&��㈪e���)�}b߄����M�\1���l��[B~�ᾁ��mU���a*�'9�j�k!p���lJBS��gS�.I
������@�M����	 �{C��F^>��|?�eה�ľ��".��1c�Q感��"[�͔��������I{ul�&�lk�}zk��pe����Y�_�)���l��t�ڃ�x���z\F���s��a\�RD��T��u�2򾩄��}�ː���KL�ح�������A`^nc�����IfK'pA�V�%d�x�;aOY��vp�:Ӕ��t�9���p�G����x��!�l�[9c'Ϝ�����۶���,��FG3�������Y��V8*)�50�de�M� s�KS|?(�����J���R���S@����6�r�N~jn�&�'N�S��g�����Х��&��\�f�� <&��������N &���l�|�Z4v|f�H���B�Li�L�ڴ�� �F�<��b�[k�A�0��ݜoE���Z�D���D~>��~)�@y�sR7X5���63V�_Ѓ}xj��SF�^Q&0���D3e��GP��^9e��c�h5���N��<��UȚ�x� ֝tDf��(���ʵ�3\+�������Ô������L�MΈR�E�!�Y���Qe:�_��.W�Znx�ؗ��� -���/ �0X`����\�/��e�`�/-Yvu ���+)��GuR��)k���U����TV��kO��A%���-2 � f~/ג�{f�YY�"Jh�+�m�秧��/*`�٥,:��[~�)[5�+>�8>)#X�޶�/o��E� ������a3�	��a9���Dp�OX?<�!�(J�'�b.���!-1)�\ZZ�!бs��Җ�U� �+k����(�L�_.��*(��f�j�}�������'���jG�a�uہ2���u4w5�1 �@��L��p�8�cs9�T���Տ�8Xu�ڙ�[�s�Şo���F�0S93S�ђ�>��~ �w:��
��GLq*6�|RI5'8�w��~�i]��%+��Pb���}Fg��ǻ&�3��f�j�$筈{=1���n��g�`
�+�}b�F�t��L��nP ұ.��y+3�V�SS�B&�Ѝ���*�c���@Ξ�����$��@��k��S�(qx���&�Wn����-%^H��ESO��p��&0��o�L��ډ3'����P�y�z�<�tj��j�� n�ŪS�~�ާ�_k�#x�dƔ(�մ���x�U'ܐM�s5^��e�~��C �Rd�}f�}T��S�����=�����YIǽJ{V>� ��)�15;��Bڵ20pK��3yZ��ު��4�C�+$_�j�z=\*�M��9��\!�5�ߩ����dc����	4l�%G�ق�f�6t�Ω�܍X�c?]ڪ�])���������<�������ä�����fh{۪b���'¬�3`�����LA�[�8K-ҢSI��^��Yy�؄��qv9�,>���wkzo	�$]��nqfmGw-)%�@}SIUD|<7�vSj�|�z�TmZ���j
 wt<%��v��J8זg����K�����S�~ Jb���Y5lr4P�-ToL8a=&~ؗG�� ��lJ���:�@��)�����UR&m��p��I��H�2��� A$_��P Þ,�]�K+�K��S=R,��R�j^<v�HX#t
����{��UO����o{{�8`���<�@AaWl:U ۱�BT��|H�Dᬤ�Y���/&qq�c&�H"�ߧS��P<�3s369Q��P Q�f���j�_�U7�8.�/ׅv��~����>�1�\�@��̢P+`s=f��T�H�d��(�(4���f0����2�KIp�_��9�V&���DoH�&=���T��qU=��H瓘�g�B{�׬ɷv$Y-�>�u��=�������I� V�b�#�_%4�-���5�0eՕ����t��դ��uKڊ���!I	��9x?�K�E�ebie%nc	t�񺰛R_���`���k'\D�]�!���xmD���tj����Ou�
�
/�/��b�@�nLI��[�#�#�h�	f�y�Z�Ӆ��$�U���j�P���yI�(p���{=8'�k�r�Ah�Q�7mmk/H:�Y+͞ Pݷ:@=a��6%e<fnTM�L3���T��O��D�Ǘ���Pa�D��qA�yaoT��CIɋW��0欅`��a[�nd�e&ϫ7����K�i�W�Ȉp(&3	�䐘_�i{�*�1���L	d��0�`�4����D��5ܯו��ܫ�M-ع���Wkq�3!c�K�=Ul���|�[�S�L�f��U�V�_ԙ^��=
��q�'����$\5L�;p�n͏I��*�D[{{�h+��ͯ��œ�4�r(��0�4��h6Y
`P�
���hY�j18�i�޻�ՄSy����p-U`�0��촥�����c�zp��pX�ZC���1�p�V��X>˹3��MTo:��10�9 10aK��4�&\��e�6AJ	 +B�ǀ@�W0�0���m��I�!�#ݫ8��&v�ΨҘ�sd��6��
�I�J(B�D������L���W�jz����w�]S�zJ��]VW�4`p���r��St&����#8�gD�z��J�	�q6��àc�!Nbmi�������N(���;*Γ�S9�s��A䞑Ƌ����Zd@�} 
�'�����A��%5�+Ȉ3��L>�%3�i�IRÓ�h_}3�˼��,�8e��e~�o-QE��(W�q�!�g;�RR��= e���@�� �N��w(7��UԒ1� }�΅	�	���˗
]2A�;Po��ʛ�ϓ�tsێ�X�?���~`kϪ���pR{ŉ'�h,�+=Y|!AC�홨�;A�Dv��tQ�Cp��`�> �(�({=q�����.�^��I�W�o���f�Xp�4������>%R!�G�V]�ڭ���4Q�!�S
"��87�i�I���=�z�x גn�����"*x�+H���$9�o��E��#ڃ,�]}�<�Ion��
��!pi��V�%�U�Eu4� �fG 9J�2L�$��U�Cy[\:`ճg_~"a�~��5�W�+��&�f<����5�s0�`������KR�w�a;p�F̌���&�\�_�R��(i�|r���a�ϝ]��Vի��_����5���P�0�|c�Ul���YJӲ5]��|��UT�kԱw�+�w��e(L�7޹AK�7��\��枽��[��o|Í�a�ۊ��V�u��3�Hߌs��} ���ÖE|<�:+�� �(TE��t�:�)G��T4�E	�}G��}``D117[)%�Ha$Y��r/�l�O���IV������-���	=%��	�����9*e�8.�@{��K�����h��sQP�j���K ��� �}WK>��C�9#�k�zˠ
��5�[8�\�GiU֌�J23���.'54����3��ƞ��T��w?��TA�_=R|�������`�J� ���W5��%9��#��C>_��!N Α��oq�	F����%
z��kh�L��E�?Ѱ�b,m`�����wBٻ�K5J����� ��&p=n���� W���a��Z�BWo� ���t� )J]1��l:����1r�W�g�ɾ�\2�c������Y$�F2�)8g� ����Rҿ3y�6P� �"MM�����rؿP���\���{����ƴ�|"��r
�\������4xNE������\��v�������ya�m3�B�O�i&�Tg
C7ϖc�ݘ��P*�L|t��/�=�Q�j��![TR�7��&�+{�k�Q��S_����'�Ҟ��r���Zk�J�%��%En�߿�;�W�1-�����3�]`���c.PB1Ĺ%c�C?��a�Z?a���<߃�c�P,�K� ]l���;@�֑ꪧ ��p���=7΍�
��4�Lrr�� �J�ݲ��L����L�`��z�����}�3�=۔�Z	y�4ߌ���������v�,,׫�j��]fTA6��Tfŋ��sR��A=�ne P���Z�8#�By���S�R���c��/�>UG6���s(=4bcǎ[4:��E����2����wLV��fm4��tVt�i*4b��g�<d����N�Z<E�����p:E�ΐ���41�d�ǭš�83��4o��@C�}�L�e�i�����fE�ſ��)c� ��04�x7}�Ո�`�����>�.��� ��Z��������	���pCDY�����e��á�\�&�C6F��0���:�/�\�n��B߉,$C�����l�`+��Zw��`(��GGD�m�8hJ2�=S���D 簱�*����)��w<Y
^d;p�m��n!��+ �T�% ����79YR6����)G�	G�`�����Uo�;y2$) fYu����a��	RPS�.��*s�l�ve�B���w�G�.IE����ʪYv Yf_CzIy`�e�R��x�"O]-�;��;	�����Eg�\� ��w�f%�ߓ����֖T�/���N +D����&Z}U�B���{��rA��#�;�p��=vX���K�	>�+=)p��̑F�`����\`cqv�d�76���bm_7V����l�/ ���{���g�0s�6'��/�o28{N('Tv��1��M��X�HLg ���9��yɞ���U�q�U��Ƌ�b¨��rp,��ޅ�'%fA��~,5 J���Z��(`�p��ؤ݄���T1+��~;̄>��HU��H@����`$꒯�t.|,���u��,��`k]�B�`<��L�<r�������K��;��T�8�F���m��_�8�U�U�D'�$Ar�����rܰZy��w LR�F4�)��Y%����������Lѝ�Fy������q|^�r�Ȇ��63w�v�v����*A���`)�;�jg��V_L�{�� E4|���^g�꽌X��ӿ!�O8j�$�e�}�A�rE��{n�Щ�23/s��Ĕ�A�c$V����~@
����ѫR�X���^��L�˱^ ����X%Tq�N��)B����.�^'և�sg�H*.>�\���AV���/�G�����gG�ܾ�t����y7t�`���9>�I��������+����=k2�3���\��U䋏*��d)���H��y�Ѿ��A9���ؤ�:���^�qH��XR�Q���=��q���`���VaxY�S�6n��{�\�$j5�Th�ڣfT[�.��K�Q	x��Um�-��Ş�6I��ؾ��\��_X�c���� �dr����Y�g�ߧ4���US%�h6=�-�JM�K͞6���f:�"�V��S��oׁ�$2�s%3bQ�w���� x]О�,����gϱho��X}I��g��SU��l��(Y�����N�����I�u1��s�_JJ�ΎHYԢ������v'R ��P�l�3���6>�B��P�"��{�����ۏ�Y����;�5��|BB;�]�~s	F�;:��'�z�J>1�Ƅv��	Kp}I��CI����4�J���WG���'Y��6�̽���Kw2�zF<o-�p�5z^_-8��>�ִ�=��R���Y��X/QdG�/-L�X��޸r�	{���b&�'�zM��ƎN�R��0�/%X�s��SB-����ئ�>�n�K&�g��}q��*�u\B*�f��x]#W%�Ӵ+�9?H�^���P�4|%���օ�(2}5�h:� &"��S�A�{9�o���FsQ���dy�����q�tj��l�xD�<�w�K:걋�Be
��e92
M�٨H�t�4j�WW�ViZ�0��}*7��K�rH'�����jep�a�-BT�n�7�CI�a�K�9�gfuqϔ�+����e&��cf6e��EW��p�Y�2i��k�r��zI�D��2ʬP�����?v4t�0H���ǹ&9����=.:/o�d��乫6=:f�Z�jͶ円�G`��I��8V�XAm��2�YmjB��z�U�yV�b�w8
.3٬�*B�tϣK �}�����n��f�n�c�����_���ʄ�Ym��*E*UPƗ���+���ll���ji�I_t.e�w)�C�nnO��*���W�Y��y �Z�'U&t/}w����K�����ڝ�a�ܴ�b^�L���9�)�w��!x�J\�� R��0�g���p� @���ǧ� ���q �TXe�h=��c��L(�2�7�R����e������2#�P /�Av��,:�ޢ��G
���yGy̎-�D԰=�c�q ��{5q�mo����:�v4Ү���"Gn-� ��w@��g`Ƒ�?��p2���X?�>���2��uX��ߍ{<�\s�@�����/�Z(@F���RF���TXTQ�ܻ(��K8����%FusCM�s��!q
}x�bB��І�{��*~߃H��=7Re�b)f7�����o~ݓw�I��י��ز炁4E*=ɏ��ۢ��twv�J��O6��e�����Q�Í�@��g�cc�R�f� ��H��l�*kF+3��f͂�劣�s�P:V���](��k��e'PO��F�L��Ah?���Ùd}��:$�}�lV���v�AJ�Ј*�@�Xc R :��+��"x�zV�0N��R���o�!�Cu�K�3�M���OXe�Z;���y��W<�cs��	��������{��r��� b쿫�m'���̈�S���d�P����I��j*9�^M��9����(��*��5�!vd���	 } �p�.`_w�ر7F��
L	�`�g����� �����#[�3��Oa�oG����1אv��B�_O�ų0YM��%�\��(Z�\��+^�WJz1Q8�#e��x����;�����^t��KP����괃��R�7�]>�cG$j��S@��JY�/����h��J��mmZ�ܶf�W�X}N=W�P��}\�5�3
�e����`U��,�
K�����'ǘt���\=?�
RB�\���0(��mb��R˱��LU�r�s��=j��(�((�G�[ ���R�
�1S��+����jG�%U5U�	��_�U,��GA�������&�&�����	�~�{������R��6ܽ|iVs=C?��x?rþ)�tTh�v��� ��B�ޮW��!ksD���N�����+l�dU���LA�1�e޷~[6:C!����ǳm[�`�хI}��DaBBr��\�h�����V�����o1,�c���h���S\2���g>�I�ϭ��Ӡ��*��0TT���h��\l ӊ������ N�%��)5ͤB�w3g���름�I��p}؉"�9��V^w�W���L��gHk��{Ͼ��<{�䨃ȱ����"�#5=��������זּ���Ҋ��l{���OT-c�,��}?�
&�<�+dm�#<�*�#��f}ϸ�g����j29��~k�d��8���Ë���Z��Hy����	�H}�I鸰ĞA�����%�H�/���Y���`gK�M���fqv>����9���$�Vr[���o��Q�SIZSPxt�-�qs	$ى�qo:��ɹ������?�D�`��1+���0 <�|~%���!+/��G��ܔ����ʃT�>�跋�SE�gM8��h8Z�_#]6VWVV��W߰k�U!��V�n�� wJj�(QY��g�֓A
�@	�E��FO�sK��/p��&���w�.�@\�S0Ѵ�#i��N�2?d	�8�����\*Z�=.{@�gLy�K�V�.�͠ �b'O*!�IJd��(��^��(��G��j�bYN����Ξ�8�m[]�<_{ �[k����D	\��tNRE)O���	x���ծ߅΅mԋ�ik�s��/>iQ\Xub?ʊF.����P�l�q6����LdS�����|"��
RYJ�g�hب�(��� �9�:��)�O��(�L1c��P����L���xp��PVޫ���� R}��u��w �@=\�Y��xx�� '�����爱:�J������1R��naL�8a�d
�s9Ufq���زWPTf�H�$=�%{�9��*��sK��;:��ҳ/ɂ�yi���U������V��P���
Ez�[�#Y�e��L�������E���4��� �` ��|��H�!�2$����KeV���M�U�k�}̽���nv��s��b��*j�g��I9�9'�P��&Ⱥ�����4�^l(����\Ę�-RǱT�ϳ�\*ٰ�O D�e
fT$ƚ���� i���A�#TP�� �v%� eL�8��(B�ɮ@%���P�Ƽ0�0[E����ߓ�^����:.�W~oV�:@�f�k(��$����e����H�7�8y�	&~8��v���<aݳ�z���^��k� Oi5Q�>C��b܎�� X.xL{�8lȝ�J�z���Gv��3�zE��!'9�1�R�L�UB���a�T:�	��-��vH�5f��i��Fˡ|��񃝞���_�{����9�D�Eb�8R查�m*X���5� �3��iw�f�8ъ�A�����46���o���/��"h���~H^~F~�d�1hBt�x3��5��2I��i=�����a7�����/_�����^��|��_l���	=�!2;zf����(^�,�Q���C���LZ��N=	a⠫3��4
5�zޗ�G_&hw�"P�*?�x�}�o����t�h] X��o�忁+<],艇��nU�UܳB����Q�DⅆNH�1����#Vc��c;&�t��*t
��9��5'C%��wD|�Sa/VS�$�x�}�>�Q �0�W���<�<��GB��%�E\F63v^l���}�ioVkӕ�ɣx5���,�p��^{���ꃿ�=�:˻[;���B=�5v;\Ȇy���Y$���q��ò�{���P޲�+��!x��Z��JP�Eon�������4<��yG�q�I"&｠��\��f�l[����A�:K�z�4��ʴ|+L,
4����}k����]����Dy+�[���
YzQ��GAt�����'C�-�����f+�v�g�^��B<�v���=>�����{��c��7�z"O]5�ⲳ18�~��-��2I�`��gZE����#~�l�b��C�\�J��2���9���lnm����c%������>�56 ��"`�F.�4	x^]Ŝ�b�y�Pb3lE�ȸv!R�S}�w(���ָ������_�5�^��S���;�{�.��VF;	� ��|l�~�a}g��`�apD<�l'���{���ݝ�;�����^���/�m,=r!�*����y!t�������av�������Dt��K�>�!�\�o	���W��x�:={�*i15��9�Ǧ۷�s�DCf2�>;{����&'�Op�ȳ;5X
NT�\�/=�:�W��+�H�� 2RQ�����������}=������׾M�l���e>!ϹZ��M�����]����7lA�E�� 4;��L8k��(�7~�~��+����c?��O�/g������O�o�_~o�sac�k$4#��k��Jqq�-1�[t��3�_��b�o��H�Լ�t7��E�n (`4�8��YBL]K��!�O�ߢӘ�T�B��cˎ��my,M'>
�2Gr[�@߰LXj�zn���K		r�(��a��*�ȁe߃���� q��ΰ�/J�;�#y���B@:)�aC�؅�%���J��G@^����(�1�F2�ia�ϔXcg)~TÒ�f�(D:���x�Y���ja�����kw�d\�Q	M��}��N*p��%(|�A@��F�s��"̈� K?����}����7_Ӡt�x�b��Ohg���ڇvw���.B�9�/KJ!7TnDÂwS����F�掝����=
����w�\�<��(1�`�ٺ�}PQ�E���>D'��=�}c�ɓ�￿���hD~��O��(����],Ȩg�?���Ϟ:Oi�J���p��{ޏ���=��L6=�����j?� �Ӑ7��.0Gf�� �b��uc���~�� �..ձ^�Ci��{}��՛'Q�lM!|3�´�G��~]�c�� `�0�؏�S��G:�Z��@�@�����SBۛO$;_?�����K�Cp0��8���I��oxH Rn���-m%�u���W�p2,�bc��v��S�)��vKn��!��e� ���\�K����UXCȡj��=yLR��u��	-��X]${���Y�!!��T�H>�J���Al��{:*m�rv��]�z���/NZ��׀Nß
�:���#�l�ȓ�T/D�͎��.Rb�������
��̯ǃ�M��'�y�V^�y��8'�1�G�=�^O>^�&��#OH�0m�@I�������ھ��?ڻ��������cg�5�Ō:
B��`<��ô�ʡ��ɳч�싋�X9<�a=<�Z�Q���_'�nj�YL'
�>'L���K[5�T�wr@[{��`=!�}��EM�k���6:�o���),r�!�H���D�=s*Ėz�E�ޕ�qt��gF���CN�+�DP����(��>�w��������߄65'���AS���<�y������ld?��gl"-.^0�,3!"������Tg�6���f��� S�����T����\���c��׼_oѭ�/�w^��f0�)�*��M�er��������Q�� ̜���j�+�?�ب�?0�x�a����ך��:$� � &]��L�]��>�WLS�>b:�� ͣah����`f���S�I.�~4Qq��g�p��{O��(Es��$��$s:�(sO )a�9s
�	hZSJ��D+k�����%���똫��WD�$|���"Q�{�4.)�`7�^���*���B�Y��|f(�Fcڥ�g��,Vy,�Ȑ��PiA���3x�\^k�Q8X�u��p�j��痾N������t�8��l��hc�D��q�?"]�`l㵅F�]��i��Q���A�5�-���!
�3�ww^H�����f�b#n�ß�e�mao������+N����h67p&��M�f����-���-o��߰�S6Di��@�&���ج��Vyr<�̓�z�����u�����v��/~~~��~�F��ҿ�����95�(�HW默��[4[�4GJͳ���@lBk��0���Ε�?����_����_� 얭�V���NbO���&d�V�>8s�LrK�p��X�G����w%X�{�����(�����|g;�'|}�L<gF3�:�r�1hd��p|n��S��W>?��$A���|�c$���^�A�Ҷ��?�_��_���?�Ovzve���om�E���7�^�
�h:�v��BU�la���m��f�΃ʃφ�0H����kA)ƴ"��#ZH��%gEn�옌W<�r���(b�LɄ��Ӏ�~�GFG�@�د�C���l0�F����;v�t�2f4�U�,�ЋMy�B�����PVT"�L׆�Z����$�XA�E_'%�~_�DAlv$�3:� -م�)�nкY�"ظ�)a?џ�z��wo�X1>aOE(<�\��9�;��fF����������k����[R��@�^=(�q�eR�"�SL/����o4a!X(Ŷ��^C�(�WQM	]GO�62��ϼ�����{��M�ˏ�`gg_��P)��e=8��lJ�����=CU��G%�Ԯ%�1#r�&Y�g�3������77���@E.�3��\Q�����V8w$����#���Z�.����k�L6�����̮���x��7�<�Y�	d	�Cb��0��C?
��n	S`�P��7�,�w��a�T(�}=��pp�
����6��f򆃄4���`�y�yL���M�����L]J�=�o�~����d��"���U�S[��b�\��$H��~���s����!�d�O�8Wm�f!f�g$�o�����_<q��G�I�H�6�|e�į���E���:��S����AP�dn:��ړZ�A��eo��a�1m���Z%�<W7��NJk�ICL�*v�����\����Mܫ6uM�@(��������'��<$�����x�7���cpa���v0N n��N.
�G~|�"�]��1��kYQT�A ��������̩J+���P�a�?�+�hX���=9��Vμ��$��%��,���&�m% TDn\AN-�ݙh~_���n09s<�i�z,�okzu�+���Iw�fME�S`c�k���&K�d���]g��G6��X�gM�{XhZ�d~�⨦NO/ �-�N�LϹ�3�}oo���ɣ�n4Ӽ ݩ)�՘ݣ�X\z��^pۇ���ċ�qK ]72Y���j ��J�'q3nW�ti��Y���㷞h=0�_y·<[��ek�~��P����f��u�
����֋"�#��_^z�|��?����F��ϭ�vmC(�b�k���YĂ�W��Ѕ��
�@B<�{2��V��;��wH�,�[FD'�D}z�H�x�I�&j��`�yV?��J���\@���]Lwj쯤��xX'�%��r~QH�uBsy�0�y���3Y���{����M��:��������͌B�B�~���i���w&���v�����@c�Dޓo4�v8^���4R��t�`�Bh��&!?Ã�M�K���z�|�l�z]�]m�fx�a��!��s\�O�2ˎ�;���^��3}v��u,:ω{{�<������t���1�(��&yi�3���T��b0�%K��QM�k�Xy	���LWW Q��}������7V/�H��,����>|���ŌM��R��(\���H�L�񓓁���׶~�';,��:@SpK����خ��2��5�~$�o�m�r���"o���=z!�������@���"�a(k������t����VQ�����⋍;��8[t��ӥm��xs����x�"��>��,�aI3:���?cY��D_�b^�=E��V��2�5Z y�g֧���@��F:�x����wo�p��s�G5J�s�'��q�KX���FKBk+�{fhLmq�d����Zt=i:��W�;�9}l�>�Y������^��~�k{x��w�������G�������{Z/@%��@���v�鰿Ȟ�P}����ɒG��0K]�_r�DR������B��<����!r�b�Xܝ��`@#�$v��k@�������eAL�� 3v(��F����b�(!�_Ql1&���┝,0(,�{:`!C�p�c�)�5�
pHf��v��Ԅ��u�@ �ET���ɇC1XtШ,�zrq��b`糊Ip����k蔍�_G|���G�^-mb^&�l*@nj� ��E�D���� 䡕�a(*�4i��$��O�H�H^y !I�]�%3yd��ܜ�-��1q8���ݝ"�$��V$�>b��|��םJJ��렠H���*��t���GSԎ\G@G�G��0*��BЯ�$al�ʋ��Ī���ƚ�G/���@�y���bY����v��t��+�+1i�h����{'�l�s4�q/NxT1i	 ���+$�0�Qҏ���z?hač�I-�6�-�3x�����k�������K�A7�SE�`�
Zrm�J,�ˀ�pQ1qFP�c�P���{!��(��~�����N�f/N�ME?-�'�$���X4�0����sijg� ��"3����{��(L&nebT�
�*�	�`�+t��&�h~��Jsۖ	c*(Y�W�	>�a�)s>dr�,3�_�������� Ai;I�HĎ=�\�"�My9�g�o�	���n$�Ls��RpώJz5���"_˘J��7�~~����H��`��C�N��cЫW���^Xm�8��O��B*BC�_(��5�,i��d��9A�4A�z��⨕1��Z�`����`R��x�{�"��؋�8�,�k3����w���'��� | �_������Z��������ʅh\M��S���sT��!��m�3T�ۃ�%�����Ap��'��|N�7���B �I	(��ӹ�ܔ=aٽ
|S1؅@r�E����y`B{th"�g��!��K�xӚ~~c�?c�ka�����JȂ�{��,5:7����g11ꙸ�	A�����as���-S��~�����f��/	�����#�x�I#Φ��zCQ?��N�����)ݡ�i"�ӹ�$�'Z���Be!�U��W���(�5��셕����}��E$y��ʺ���L��_��b�&S!�5E�i*ff]�oy���[
�E���UN1M�[=iއ���$l!p��bA�$GZ��4���$(�\����pDщ)sI�3�>��'�ͨ�i�P�쓑�
*#�+��]�)Z����iK����hC�>E��("B{��	{�=y��y	r��+{�0���ywĂ��H�?}iZg؊qi�[��K=�����q@�^�����m�C�~>���h1�n��68n��j���J�BId����"�!
J?r5o2�W@#l��#��/�6s��$>x~��b�E���ݚȁ��n!���h$������)f炗��E�}�*PxG���I(�rY}�c
���T����������wl����&ϏB@�r���BV#j,J1TTM���>1^�0���B��Ԫ�]$X%���M��P��_�'ei���G�䂒Z����-��ظ룩�J�b���s���dȄ��2�;x�3P|��\����7�m�w�V��}d��+����ω��N(Fr�!�@��N���MO?T<�"�}�dB����E?I¾UG�<�5��g�8�����]?�������blo��G/�>��@P����XKT��0�~��AP�z􇾺�ak���;?�画��&�����G#�g V�'E��qT�J]oM{��h=ע�o�zz2)l�|g���BX�~;bQۗ3���M�Ph�	E���,"x�X8��P�ɕ�T��$�.�G�ɫ �!}�`|�Ҷﾲ>r4�)l��`z�	�)	�]�Nql,�+��d%V�r��>��9p �[ !��=�Fs�ȱ��d�ʋ9UŐЭ�k�9�a��7c&�l�a������6 y�gM>�F�﬋�_xwܿ�W礐Xg}Tv�)B()���`d�pu�`C/��#�Q�A�O�Zɥ�b�xVxϪ��hw&a �О%'F�8
��bڀ�D�FÁЇL�3
�d:�-�X�0����E����N�	�{v�0�̐�KR*�B1��=�.����$Et߱ %jѷ����F�S�A3�䦠�-�))&�����2�<���*���+YN��*<Ӱ6�"� �,�U&4О
Xky�Uٔ]�W�ܢ{j�֋����)zRmE`Ϥ�1r��Ɣ��7�(��i�?��r<���P�x��BW��))e(����L(s6/ �)�	5pb}_̦�m���ö���n��É���,:{�ˎk�{kX�4�~����)��`�&LtE57�ē�Y�L���S�Y�HYC����UQ0���Qw�PZ�#�[Z���z�������+���i0�8���1Ś��bn�N&˼^]Krh;��M�$'k�EqMei�UUER4\[%c,!0�"tf�5<���G�E>� �N��R�0�s���q.�jN���bdw�_���6�%D��u�L�N��
��=��jX��K4$��4[y\��5T���<Q�w�Wh*�\��	
c�<��zQw�	��Jй�	3J	}ON6�ZR,<9-�R4)�: �o!�^����g��	��?��喈��,&L��tſ7��!�$>�:���=r�hT,h�,6^���d�����A�2�i3Ւյ�P�Dc�K�n���cz2?��d��dxl^__Sh��0W/ZY4a�Ĝ����.�ӖIU��@XA`��Js ���V�mI�Ċ8!�S�ӊ=��b�i ��dP��>%�9'�L �^L���C�Q��vL���ɀMꚚ9'��?:�c�EY���ў�Qt<kb�%H���E9B�_�����S���D/�3;�����������a�7
�S������56�Td�����۠%X�����2U��5
p
�I��H�D�J�������q}��K��Zυ`
4�>��՜��gp�H����d� ��Y��r����z�#j�J$j��k>�E���aEy�u�JU=S~���v�Q*Rs3�#���Y�RM)�l��� ��\MX�r�b썜��8@�n^/T�Ì�
��C:�մ:�\Bo�k�?�%�@�P��vGUk `����y(����ײ��w�[���! ���N�\p��i���E9K�h�j��Ů�G��i��$�t�^$��xBd�#lT#_A�����ԳQJ1E
ݍ��\)�㚢��؏B*��[���Ф��F�k�P��NM?���5,^��/_[�P|uXw�h�uT�2��8�^^؋W3���i�>
�,�6�2�#��hm���ݖ�\��twwO�����������m~~�7fb�?ۯ~����_zγ���\��:-)����(�	x�2����gw=��b��[u��J/~(�.�]��'�����7ZcX,��+m����[�r/+�'O.��*/J�w��lt�qӠ�k�a�`���S퍤�":MmOP�'SAAx]#U�.�?���i�@�<�����Ձ�AIy�㊐Q�7	+Rϭ��UObq����%baHy�T
C������BV��D��8}C�(M3���v����]/����ˡ���g�}q��p�$��]F�#x����ϳ<��W�T�����s�D m��f�FG�ނ29�e����:	�+��(�*��F��/��`0����t<���lz:&�� �c(����� �U�k8�p]�t�!�k�VDa���ЅߊE ���?]�؝?����e�/@�*	e��=�%Qov�����vqvb7���I�x�7;�����Y8&?�֮&�O����u)�����<�ҝ'e�ܡ�Y۰���Ը0��}5���ڄy*���7�h�����Ϣ�"\q�"rq�Dg�nd�� <H��M��'�.y*j!����řݯK=�є��(�|LL�B�������8o�>�A�4S*!���h �������௽9�:e}o���&�%!ݔǏi<�!��ۑh����+Ov{�޿n��ϯ>��<���
�$��%O�B�ԁ���ZHœ�)���9-��ho��0��¤1]�n�O���_�+�����7�\�dv�r �*$mط����V��$g�{۳�J$%u��Da͐o1	����~�V^d���ا�d?����<´����6,[���|�\J<#p�������{�L,�?��{|�������.�L��7��^�	:*@�$��k����m����a"����Kv�%����Y�?U!{򵏘�Ǡ	�ɕuS�����R�e4G���f��^����R�:�.x*88�Ͻ�����Ѵ�I���fg+/r;?�:��;ԑ�.P��u�DRSȂ�H�
~XGH:����@ޥӐ�d��5��:�_/�$h
�QL�pb�p6�����V�@ܿ>8��h�I;T�`��vi��Ɗ�9u�4�W#o����y{�`�`�uQ;L"�,��0��/h�}`�1�����la��ؚ/0�nx���+�R$�J��ĩ�XLk$bl��NA�&gt���/�2J�w�6�\,xq�WL�׾o�<7����ғ��	떯��[�c�l��e��h�?,N{��2Q��6�D��i�PN�/��� �����ƶ*���ǧV�_X]�dk�	89��������;�ϴ��/�������u��ڮQ�x0)x��x��'���Y�^��Gĳf܏8�m<�S�bi�fBC���s/N��)����1�J�>Q
�����IB@G��QĢpBá�?&�]\��S(M�=g�}m[q*�\����Ǘ~=/=�R��Sʦ�|1�sY��$I�A9m�HЩ�sj����4���*%������_Ά~��� ^cD����?���	s{"�!���Jw�6Γ��}1�b��x��$iLB�G�)��P/�G3�D�̥
R��V>�}�#$XSe���Jv��'@��c)��ɹ-.>�5���o�=בl�hX��.��)	�Y�b�8���r�����@��k��A4�˕?�K������s�n�{��L�^/�W��D	�T8�"��O�
�C��������P۟�xi�����5��͇�����-5GF�J�}_׈��S�x֢�q�4QL�v:	L&�G�*Yt&��A�]����G��o�`?�������#�䇟ۃ?�/~���g?���_�l�u�LPq���A紘x�SQY�OF�@	��I"Uu��������8�F��/M���7���,R�)nP�	E%�2�4���s����F�R��-�m:�4���h�S��!c�%��aCR7�O�Ux(Ux���^�L��@��0�q:�E�����Vpp����"+�T$gENO�-ԝ��{���o�h�I�R܏�fӉu�����ʉ ~0w���IPcjC�UQ'7�x�<�,�������9hi��n��7�1���p�~Ϯ=p>��ͨ�N�)��]{j������K����n`����O#���d�G06���aVy��k�n�1.n�� 1&�>�$Z�{�� ĬmBN{� 
0��ܸ�����%~t��<��F���=\3�����/l���-�NM;�J��s��i+h���~�_E{F���m���f��О]`v�' �ًO~`�ו=�^s�sw�E� �����R�;`@��\l��s��+!-��X�zn����!HK��2Z)���+;�:����*��P�þC�~$5٤L��OJB��PS��� nR*~���=}A�͒��&#��"7��."�,d}R�)��G\�|��UW�}f���x���{�P��?_E��b��!�!ȯ���/o��o� �|��	=�FQ��*�!T!�����Oe��7�UBAM�= ]�vk�2��C �#"�����O�)>���!���fds�4�@��W_��ى]]]�痯�ߋۻ;���������)�+�E�[cr��/'�H0F��֞߳٤��������_��?���[3�{��S{��_���<��l��	g�hhm+¸�U��5��=n�fS���V��k��?�O=yQ`�I<隆���4�v�l��J ���}���T܊ �'ݔ,��u͸��>�t���<�Hk6�
L� ��g��m!\D�^�C��Sc������g�`S���(��ψ>��D�j���a�g6;�z��g6-�^jO�0���_/��˵b.����'̔�{+�ԭh���3��(�Fe��V6"4�
/$�]����*�9��P.�og�g�y~h��?��O-���ِU��F�¤0h(��D��u��{��@K�b��:�x<G����!n~�=6?��h�AA5�݀6R�Mhӄ����,=#%�@��<p�^������ ��)�eUB�;��|4E���1���J��C<��U�~FF�}�IĪ�¿꥚�\}��w_[��U+�:�
 # ����3:��b[�/�l�G dP	/?�¶�?綴W���{=�\�DFt���1��(��\�x�qА�b���e?Gp�1$iؐ36#�Hw��}J�+�����&�:P���r6�N�/|�}m?�7_/�/��W3���z@N�Uxh�k�9z���_�'�G�m�\�-��̆��|����O�p�ӳ��>��&>��D� 2����?�!Ŕ���}�bb����ܱ�9�������;�n��_��T`*�fnD�t�X��}�(���r�%��x͈����.`��x��kj�:�U�LPm���B^	FDe�e���\��"�~{�=��X{�>{qa/����V76���݄ڶ)�ٷj��1-�]G����"��}c�P�]�L�1��W���z?n����	��V�Oy]L�Rps4�y����W4�\���b�wwP쭙/�G[���<��E�}��ӎ�����r��J�jo�{c�����9������[����������.N?�˗WV����"�*y�DPVg�y��^��p�T��L�B��}5�a=����E!�{����_I�)?f8�h�W&�4t�J�w�%�;X�T9��m�Ҷ�0��U����(0�YJd���ԕ;��'@U�ݓd�s�b�8C���ɔf�ؔ�1�,.ʶ���ۏ��>�'�b��ܼH�0�94:�������ۇ��0�x_���	';�"��T�� � ��_�XD��h�ô�����P�̢K�d�Ȍp�̉�rT������p3NS�	t���^~��no��z��A�C�c:qX�TN���F~�>�IR��?�;���FN��3�w40���6!H�ř��'Ï�x���׶���P+	B2T�^pA���0�:,=9=�%
�v`���V���M(ZA�� UV
�v�q A�.8�}���e�΃�#9���^ڣ�����hJ�d�@��ʙ]J�U$�	�F���Hv�S�#��TD��R��uK_) ��&�?�m~�oW���~`w��:L��1�(����'v�:{B�?��yE[��?c�����yb�'��û7v�BI! ��'BK��W=�aҁɎ�e���_��N #����5���8]�1텗�.C|L�Vh��uN2�g�ͣ}�k���6�r.�� t(��]�Z����؊�]�:A-�PF�x� u@�U�gM�et޵�\���aknk�}���d�E��V�G��\F����J�з�������k��L����"F���Q��Y��Z�<�d4��;{������xV��')���F�\��o<��A���B�$�askh��od��yO�g$ih�ї�8��	�j� �g$c'`iG��r���R7ģ?������E���SN�i��d���|D���(1��Fܳ���X��$��b9S,GIk{ �p������'��}���x�PѾf4=��G�]u��eH��]L_zf�uJ�]����w�1�w��&Xx�m&˖������\}�N|�g3*��n}���������ĴF�J{����QE塛y�Fτj����(�sy�A���b���#�#������H��D�a��m�(��o�-;<�g���l1�<&G)Ϡayu���8�"=���U�?*a-hk!���BfF..��=�n~ݯ쓏?����l�Z��0��Z)ZM�� �Ĵ~�g���&_F/V�;�哵!�h4v��T������v_�y����S�0xLT�ؔ0�Z�2��#I������jx��=��Ί�Rc͐��7�0�&�n��j%�� ��-�k���:99�eFhL�wh��E W���>ζV��T\6�&^Y���F�0'u�J�Ҷhj��#� �@�b���h�.�}/6���򊴐6 	�H�#�2~^n7k�x!����+���$6t��%��J�~6Ҭ�ʋ˓���>���"Y'����F�N�@�(�ū
���,f�oP�mB�M�%X2�I���� ��<J@q�{�(e\��?f/�[$��DQ�p����'?������mm o�ld@��|��H��#�D#,�^���l;�����d>����9dl�Q��@���cGn׷�l`-�D�e�I4K�,-�0 )B�6=�g��4�4 <6 �J�d���1���Wv�{~8_���;��|�tTJ���H8<Kh����y>2� ���eéo'�����T1!�g��e��d����h:Bb[�o�'��^�,l���~�[=��?��f6��{"L�+�Y`w{��{�R�
��'M���_xһ�%$�a�E"�l�4zV֗�D��mk�nn��|�}z��Qn��k�!� ��7ʖ�Qs�)�<�M\�D5��-t�b�c@���:ة��ap���c���=�G�������x(���a�������n;�Z�4�,����Ϥ��(
Eh�]�������|����^s�t�>Ii��Z-�l��m�[�;4��>�  ��IDATZ�}�x�����JO�^tI�ƞ��]L��'����2%��" @��w�iP���;���w_{B5���>��Օ]��ǻ���g�_�$:��A���q�gO��b+��M�����Tr����k���kN*��~kO���9�\v$���)H�_��0���vg�H��a[�@}�޶����B���2av�`�,k������cꐁ��������}���4�n�.�I
 ��M�kc�BQVOEp���[��ڞ�P
��N�b(�Qɱ�)��[��x:G�qd'����'ȁV�l/2�a��4=�T|��f
��擦�y�d��BK(�� ���>��d:����h1@�OQ�;��������=/�)���mɃ���,�}m\ۻ�_��{�59�_��f����)J���l����gJ6��A� ��v���|�ז09��Z�4Xxz�ܲ�B��؛e!�ء. 'Xm�yY(f�,tK�L��'ɚ�e��G�yc8x����1�<��R�M�\ڏ��m���B�'���ib�f��P��*��?������v�B_@�`(��ɩ}��5��w�~K�D��(��]������������o����϶�����0R�(t���^��?�c]��U.��x����I��wP�,�Ls���-��vW;�W�!Q̀�ͩ*ws}l�G���4�C�V�6%�K�#�"F�w�mq������l�ޱ�=�~��=x� �7x���ė�e�=�1�u�U���$Z�􈡅2&4� �.�H�����'� L�f������0���D�Oꛃ'��Xw��py4����K�{|g�͵]^�l�fBS����)�c�,^��������'}(���:= 71d8*ig�()�	a�E3��k�&��%%Wź�M�$�#DE*y.Ba �D+�\ϼ�k�����Ӵ�NQoyXٷ�o�H�"B�'�-c7D���EB[UU4�2;��[9�<� �Ehz&{'���b0�	�`dj����_�L)
A�"$���P��cagc���5͕�Q�G&�g��Xj��lP;�Xx��`����h��s��y^��ŠL�%>�快!��E�F,i.�.`zO��%�VY����5ǾB�ԯi�nxφr%����2��i�)�6� ���cn�T��3βN$��������P�g��ۆ��x��rb�]Q����ݣ}�?���?���������ST�4�S��E6o{٢������~c����Я�ٗC�q��!�@�D�_����n<w�t8��n�;NAw��熟���m��c�5T:�~�ښ��k�"@mB�=�����,�����yR��4l���`�S�T����_����n����@����x�1Un����Tȗ���3;�?�*��ú��@�b"��|�|dM�vܻݎp.曜۱�WRI�}�"��^.�啕�5�Ʉ� �D���+�}�(�I�{/`t��,S����q�s��{�C>m�D���~i���L�:�_��K[L_�d��nO��oX\�q�a��U��T�\���^S.���+�q��mʤГn�p���:��(�H�eռL�8/ \R)ɓ�զ�����#������T����B�/S�V���e���L3��R�}l�.��R�1!�`����jVx��p6�h )���@r�4�E�@��:E<z;N���C'ܧ�8@�C&s[_u���C�7����It��z��2�>�f��~HM�6<;������f!���Z�S!g�+&�I�IG��d��;�����5��Hސ8>3�����Ɠ�������^M��	cY���(�٪PM�{�4+�v��s
���"";VO�C��X��f�s/n�f69��|<�@���jO�>��y<J�3���=1aE7|���&����[���Ͼ�����?�{k�|_���`4ZI�9��yZ�:��"<�kN�n�˷�OY��K	Q=�����٫ H�$%8��㽉��G�j*�9�Ԁ�d/��#���6��p5M�mb��ӁX7 �Α�ν��ϕ�tm�A�=�ӌ�� kO��W��������{X�����T�DS$��?l(�̈́����.��vu������{�>~g��_rr{��s��Oi���P�-	WN�,�T���p�`cj-���5u��u�|>)�ᰭ*��OG�JA��S̢CO]z�	���A�d���#+�'])R�ԓ+ <d~����.=5ZR+�gr��h��j+�1^{@�jF��F�1��i��x�Y.��o��E�h4b�zr2�]�ۋ�*�>/� �c�	9���������/K{�~��Άp,���������fm+cS��A��I�G��v�s�l�f���xE����>M�q�!a,���C�i�hf'DM��Yj��L&�ӏS��=�^��8CB�=*��)��>�'�/�~�a���Q�{���tQ�x�|[_C�]�j*�����ώ}�,
�Q������M�8.1�9�,����S�}\����זX�\xl�z�{��gA@�E	��r2;�1zqc�p��i�������7�����~l?�����g'����w�������N[�,\6��+����
�?;��;K�<��� ��B	����[!�A��x����T!,�cc��`Ҿ����q�-45<#[&�0zG|�q����mµ�D5$�	�ӳ@���D o��%yJ�k��gMt4���B�����a#�;>w+�<=AqYx/Z60	��	
N�� ��cڄ�ZQy��׸�s��?m�׷R-dq��)� T�?�����KBw[M�P��'��"|߃�*��1�Zfqy)F%���j�xm�ٺ&���r]�]#�B���DN�7��)���?�$�	^�(�aoyk�ZgR�%�P���6��q1�sM��)��Bl� BK��wUg�fC�-���ǔ��=5��Z��=�9Q�e��i���t�9����~o������z�USa�8�/'���_�g_���on�o�{�%,vD9��2��n�Ⱥcޱ89#M<X����z�O�b�x�U���=�X%�צI���1��o/
p�bE���^F4=a�����4-�ª
k�a��BGJ܈�w��V�=��i5��1ތF�ӽ�G���^G������(<�E��Y�g��7�2��`�
Uy�ؽ�O ��a���`�< ��dx�h)��-S�I�ͮ��g۪�>-�0�ond�2�`�m�n��]��CE��n�"�F1�G"���B�d�w~h��
��E��mM�o1&Z/1������|~S�K�;��8s�SG &	��4�1Q��鞂W~蜽����ؚc{(L�ߥ�A�61
Wg"un�M�p����>]�s8:$�geLe�
ލm#��lz6��š� ��D�xb\��߈\+oe֌`��I�ct>�st�M�2=�M-���2sS��?R	�te��b�N���hX�է�S��0�zH���v���$,u��JY��{��I�+5-����A�\���/8�|d�6����f�s+�u�A{����3mr�]$8<��c�;>�[���%U��1y�_�� ���R\���Zn��s;�Y-w�
f٘S/t� ݥ�7�|c
Y�����'��|/,ٹ뚱��͋�͝�{�y"7Y��3���t#���xypQ�0��V���� G�ȃyOO�5�l1��1�^�l*5j#�J�(��tԱL�v��י���]Ҍ�Mx��3�t5��LYq�=9.FS�Ⱦ�"���9��Q|�[���HG�p<�,&]�qm'^Z�N~P�j�8�����b�E��]�1Ms���@��9�
~Zn�����?���������vy����[�|�d�I�lvj�ug_}�[��ri����4��<O'�O+�j�̰)��	�&�)�_S�����#0M��ʩ�������`|.���7��o7�c���D�:O��"�@��Y!�x:b)A�\qҤ(�i#� GS�){���t��Jx{.���+u�1�� [��L�K�^�0_Y���R�h�!IC2��ϑ�ܰ܁����j1�W�?���K[��w����MY�6��~����o����NTC�����c氂7��*��~/jO���Fe����[��� Ñ���di���h�܅j�nR�k����x�05� O
O����V �\m{xHz�M���{�+���-im���<�K_PጢQ1{O��?/ê�i�5+5��igR��dj	x`8��7G���j�%dt2��)��dtvvFX>ٰN'H@����(*Sz!~y9������~Ej�� j��^�UӁ���ҋ͉_ρI>]A�y{�W�mw?��`�7��TWj��DZ̄j������@��Aڱ �8q4�D�l{<yuya�_�l���t�b����p�
�I2���r�֡g��?3�:
;"�!� )�H9����.TK5Q@Z���{���0�ؑh�,"�:E&ZC��'>.�$��iBl��]�����U����,����9��"+���ݯ���q�YA$�}f�����]���u#��z�`#��C=�aU\��y������>&ME4�_�v#��I��4�����ϟ���M�2&h}�E��n�؁���E���(�ŭ�b�{^�yqg�y��[/+����� I�	�vw`�H�NbEs?�ıH4�c����=��X4��s
|y�>��U嵭Vk�t0������/>��������՗o��[�����1ܐg�ٖ�#��ů����Х�wx��A����l�������>�Ob,O*�ϋ��%��ʺ��epQ�G�%���Ē�Y8s=G~^�ZD��	�L�c�uZ:�B�k�9�
"O��Q��,�s}��~]��<rn�6�}x�})�O�|�O2���ЛQ��X3T�F���f��^p�|4���mw{�УQ"p�K��$�=8�ۦ�4vۭ}����}G�{�F^��Y�BP��r�����W�׀��T���I2wZ$�S�X�cO�Zʊ�H�>lR�k� Y#�TX���艿���'��B��kN׌$�V�x�^��y�'IR1U�?���_N��e-�8��`!��u����d�����&7�s�$a�5��S�z��<Ԟك������Ob�x�_�(Q��AA�+�$c��d�!�j��3� �X��B���Cէ�.덂~��剱?�JH����1���4�c�~l$��p�7��&,:7�=��#}��l&�'=!�!�\4����U2��Y{i	;��&Zϻ�؜�g�xkv� ����kz��2�d�b/5=��r
�/��~�}�����`o������޽���l��<�D���K����������ALU�)�I���*tk�m�������]�`����7%l���!����H��J��>A4i���{*�@��aX2:ȃ!���B=��C�r����e����u��_�y55������.?:�ġvl�rZd1�T1���a����
ׁ{6�Y�[|��<r20P�`� * ����?�����_���{�>�>byqp9�>�wwk6kf�/�[k�%�\��%���$ �0&M8�{>N�pϡ�����ޠV��%����P� �;[y!����6��R�P6��)=���Z���'���F�G�|�B�L���[��-@ZL/ؕ4l=9h���y�CD'��u(g�n��X����=��B$���(zN\�!��|a'�'�;"��θ'g��V�i_�[�O�����۵�\�x!{a���	2�v��>���}9����~�{��&
?�;x�bG�$p;���3�P��{��X��vp/�.�z�^�Q@�2uNo�\q���Kj�a�C
8���<;W
S��n�&��Kؒ��s4^xB-7��VA^�)�$����<Bi��8Z����;2�Q%oQK}��F1X@��WB�2�7↲xh-��DT O-AŨ$��
�c��֟^s1��g6�(7�;�߮�~�6ڬ)z�{�E 8:�x���i��@��i���>ڛ���奝,�����u>�7��5Tjm�����5����:8�]nEh�Ф8�gڅ��]2?��z}�M�#{����'�є�k����ϐ-e��Yg�F��s�|�\G��#L�?�F���3���ov:�5	E�1',��.���
�$T����)�z�*/a�yL�� ?^C�Y�+'C|�x�d��Y�5���A^��|~b�Ō�v�^s�S{b���tfs/����?s~zb/�NE�=Ш��Ka����"�	�
X�	����S_X��(�ނ�$Tu�\�@m4�g34���<>��^K��P�f�������+���>O�tMec��%�P��ҙ��ȹ\�SC�_%�y#�� ��;E!�rؘ�$eR�p�`3+�h�8p��	:fP�_.�&���g��>P��Ο��O_د���z�����ۛo�rğ�&/>ʳ���o~n?��O�� Wt�Z�r$H�,�g���G}��"򧦓�
!"��s%A<)j�Y��㙹�M2�W��!W9�2��t��R�[#_ￚ�@��Ǝ~�$���!�E˘8Р��܇e��Y]��%��e���Ѓ�;�*L.w�T���!L8�Ԃ'��P��Ж�&�Xܸ@����u#_r�)��E�d~�q2I��F� gǖ��7�ɘ>/"�P�`�Yy�f�ɶM�	@^h2��<1�Ѩ�tP�K�b̟����nz߆hJ��E0b'o�8N9yLn$l�G����+�_����Ź�������#}�L�f������Z�^�!�wt�.ĎU�r�@�8D:/, �ô����H.���m}wO\3&�L\�a�R���酝]�����:$�0 �1��v�Ô��x&� �u���b!�O�>��c �����d��S������_�����;�
<��.�w1�65����Qr��@n����?e���r�kE31�P���k$��i濡��:��a��W;�G��Tf=�á6�k~@Rr9����+;�u���v��Ɵ�b� �q����k�C�����{����C��W�����M8�f��m����җEA��Xr��N#L���x(�mxU5-m38�-5��f�$�"~�'�n}<(�2��[j~����ľ�~��J*c������f��	��p/��z�*<Ѭ`�a]�"�6S�����Iq��O�5e\��.�q�3y�����n�F�a�m�͆�r��Ec n5����-�(�<��qy��~����w��j}oo���8g�t«fRG�	��W����>���%.�N"l|81�y���ǜB�7!�D1�NPN�2D��}�� ����OP��Z����n��!�@�'E�4��59A�Sa}x��pK�p��1�A�a�)HS����fm�e��h-�ɂ����1���Sɯ���n/� ��M��d�g���=�b��3aä�������?����w_{R��jװ�b���Ҧ�)�T��ﭮ�F_����4&� �}�B�?4Ʈ��/� �R��ݣ�>>�t�^��H��F�ZM���^j
���p���$�D��� ��s2-O���@!�بZ��D��I)�x��y�5�Ċc��1��ށ��7�y&RD�BB�t����J6��D��(�T�<
�q3S��<�P�b��k��٨9�/�� ��F��~����7�����Ƴ�mQ8��2D�v-� �����nn�[�0��8���K�ﬡM!Su�B9�
�g<��͔ޞ8yuğčo�gO�@$�l���k����9i3w+��7ol�\����Ly�$6H ���+��e�$�<��h�����	�F�CS����P9�-.�,�x��Rh�Д��AǄ�;��"��lDÎJ#�c^vTZ��2F+2xɦ󦄀
^�>�f�h��5���k��+(>3���nc޽�{_�3/?�:�S/�g�6	e�f�*����(ĭ�&�i@&�C*� ﺙ���q�؆�4�:���K��T|.ؤm)�U�Y<����0T��MU��RMA�DSQ㵖�.��j��l����"���[��|����c��Z�5[�C�>fZ���Cǜ��\�LĶ-YQy�)> ���מ?����~�����@3M��0���6�� zB�F�&x�߽}��N#��j�]���l-�l*��y��\$�l�9O:7����蘳�O
�]�r����� ���r��iI~�Yhlh�%]^4�9Y~V�X�81�-��ҹ����8�_��R�8q��l�HHOC�r�45x�D$����ո 9� ��n�V�)pz�@�����>�Ѫ������A/���{ЭDGp�ʓ�҃Ɂ��5;:]�}��3�B�$Q;r>���n�C��2'0�6�̳�g#�D�ˋ�"��*�*�����wv����a�Mń�Rу/ 2ب�cwu�L	�ݒ��g19J�����E�"���VXGF�h�
�U˃<l}�є��?�bE�Պ�b��h�����������������^dH���6u��|������e�
�A;>?e�̯�h����Y�)� �Ԟ$S&�`�� *���`drtN<����{��A<����<�b���b�W�����HΐGV�)D�1 �w���>o)O�;��B��P^B��#ttwx�s;��v}t�br�W�`���SC}��4���i���6y��Īl���	�$�<T������P��g��9D1�S+fS�"X�����z��\^Zy�]�^[447Q~0�B�E����a:�r��pt�{U�AL<轈iyxu!bR������KDၩ������e��	�!�H�I��4�ǞK��IoB-(X	Mh���Ѐ(Q$*O���� ���ZcU��$?��g���>K�x�a�y,"7g �j�!��T#�s�����EEC_T$H+O���^n>X1������|��ۥe�@I��'�v(��>"ēnn &ހ��{-�hD�n3
���@��5|ؠH�DB�,�LO��(�G���2q�R��~���0����0qG�x�k���&<�B�8�i��u����a1���yq!�A%�
u;���b>\s�P���j�Ŀ�" n�l����.>��E(��=���s�+� =��z@�
R�8'5��暰@�����[*�y1���?S�8�{�����0�nC����G�<�Ĕ����������?������}X�w�^��ݝm�� Q�{0ʦl`�=��m��
~X?0��GL�/�x�H�%�s'C���T�+�:C�r⹟�P�}�f�8R3��{q���ٰP�OO��$��d�Ks��!do;(�\�:ZX4LN�x6�D����eDO?@�, ���W�P�Ϣy�E2>j��aC��;;Bё���7F�ӌ6�P_3�;�W��(�'=�_m�woEY �'�3�f�D�T~�!Ʋڡɺ�iBPI�ty�~O��w������9��k�>�U��"K8���M�4y���.�X�i(����3��|�y���͇;_�+�9�B��=��_����߳)/�%�W4�����Շ򡖪�%�2h]�����q��Q�lD�Tފ�#���b%����>� &�ɂ��^L52����C�?mJ^-���?�n��_�um���-����ĽC���<x�F�ZCܻ���L�@c��}�������lw�2�l	�}BX��-�v*v�b�&+i:��`*�
�gbjE�y�����Ο���{K�E�<#��M�Y(VDGǽ�Y�(����P�*���,�!I{�I<��h4`��z���Ŏk8�'�+��2�������X�ħ2i4l&E��i6��{O�Z6q���3�Hf�N��ۮ􅆅˞'#/�W��غ���y5�b�|���N�Ϲ*$�H[�(��Z��,�&�;j4�N�~BxI�\k�ç<���/Y�SSj	IQ��US���&�;����b�}!���Nv l�g��C~���j��E�F��ܞ�Ϟ�@��wH��)���<�"�W|W
�����
l(���"�Y�R-Ƕ��gӅ����
s
�ך��2Ԑ�T<��#U*bUZ����� �`�sF4?�ka���\�H�o�8Y��r\: �7M�,;&)jB��� VL�V'�E�"��f�aـ���q������P�HT�W���OjF�=B��px $<sl�>-HO+���=����q�S
Xä'ԥ����y��#��=����:°�@��!��CL��? X������;H!kO.&�()���Z�F0
�RP��K���2ֆ\���NuL���g�8��M�a��W�]~@���t�Q�S��4A���_�r��#g-:��I���D��K���?zl���ژ*��������C�G�2:G��i��S��T/��>�����֨sUI^R�����MS{�A
�k���'���y���qu���7�:���K���'^���oZ��*���o<H�5��m�4��b{�G+�:�ç�j@���%!��[N7Dk���sk����t���1�����%N�Ś��[Y�WéN���
���S�W"'~o|-"!���V(����GUA�h���e��.����a����FN:��{<�Z2�i�x�1�ϱ���=zO��*WFp�ꐰ��6;�����W֯n�������6��|����7I�{�~�5��� _j��|�0��Ǟ�Pu4qMq��xH��c5+J6�z>���k�]K�[C��8�hC ����h:~w��R�6,i��L�Uj8D��+�A$I���� �Z�j �^�I5x=�^P �y���G�LJ�XDG|�|�FBL��7ͭ�1��!Ꮓ���?a���wvՀ{��H|GL���Ch���<l������xk���F?���K����Z��=��o�,{��;����F���^\��{����?����ަ�ON���V�	����J�Q �0�_?z���G�t6�>�XÖȇ�*ܘ�o��</ �ljN�Q�A/���s'�=$w�U#/�����/{L��7��8�;[�V����Y�IR�PH<{:˚H�%2�m�j����F0f B�^�nł�q���QNU+踦iI�)��M��������6��G�����ʾ��ol�ڊ7�{y�� ��{���ڴz�
�D#�#I������ ��a���m�h�Ы��xY�Y�?�8������.��c��eK���D�u�*q�A�Jl��ņ�֚\�����[z�z��h�F>��fs��%a�g(���sX���V��T��r���<�N�0H&����������U$���L,��*��>��C΢~,�D�{/ں����~��<�Ͻ�ySU���.�� R$E�H���Ўf66b~�4�F�FL���H��J�-@4��\W������n���V�����zu��e��<yNM�$Mʫ�gl��WJ���h���M*ƒ����6�t��1D�C���?���/��ζ�_�uu����n�w�ӂ����6�R�ÞSC�p�B+�吰f���P��x�����.?<�#�O{F��4:�ˎ1�"+��1G�Q^��!�c��8����cu�`;* 9OYj'p-#��ۤ�T�g�1��c��$�|������a�Wk��Efpb�ҳ�)T��U̧Q=CS�d�&��37��Vju�$�&2��+�2��a�N�f�Sɶ?�]k[g���v���$�c�x�]n�h�Qϋ�&����0v]Rr�BV����L���$��nPf�7e!��J�#�/p��͛��}�s��ȉ+��\۾|��g\Kܰ��Ʃ�N~���p���E��b��ք��x*"E�g6���~��PH+4H��p��^o�yzZ��	Spb@%BvW�R
�z�צ-M�]���V�L6:���uR9�	O虒�*�\uH�-LAPi"�.5���������u�y�����JS��TF��t2�&��Ҁ�M�@�ͪ����"��y� ��!��ny.q���r�����{J�w��5������i�C��y��%�dMA!��Ln��=)I@�<�I	�E��R��N��|�ʧ�7�rz�� U���"A�%b��&i��KG_0�X��-�h:�35e�"Vw���]����b�gF1س��	��%,��X�o';������b��gE��a��E�^8�^�N10N����;~W�1�_�{���j``��(��������x��\�'��<�OHѕ��$��1����ؤ�h�J�9!㊦T����-#
T�O�v�v���h�	-@�b�Ϥ��~�v��;���T�v��n�Z���v*i�i��1wv�h_��L
#���k��I5�6F���nu�l�� �-KJM� F*:'��ZZ z:�`L
�n�͂?�)�o���)G>������2q�ƺ��p�xՔ�"���h�@�&������pKi(Qe��]���P K�i�<��|��|��$�������T-����qzq���ֽ~�*;�:5N+��l`�9I��,�~Kca�lށ�g��v#L�i'���;M)F�@��I
���.�@��}fu�HZ�'�pU��fx�-��yҮuĩRV��;�ؔGA$�zrbA� ��Q��wިT�4�����/�`}����]���ю\�*pE`OM�{�5�K����6���Y�R(h#�{�i�,ŌJ��c0`�o]ȇ��G�#|�~���s���F����������Pӝvr��}��W��a����542�SF_�P������1.ꎬ��Ja��XӉ"l�x�$���7��G
!�
c[��W�!�RJT��%`H�x�+Տ�@� ζĀI��h�)	۽bs*��ܕ8r���T�RAW�v�bu9+�t�i\�`���3���@˨ظ���ی�m�
�P����� kQ��{��3f���F�&Z��w�E��T��Jh2J)e�q� �wzlR��!�g���3�>4##�u�W������M��ך�(8aGZOBv3�����<���M�˓~L5N�'���JA�����+�gT=V���a���Ǯ�?[��ka>z	�X~�Ղ�O��@�N+�g�=x��tmB��[NETc�|N��8NXAk��7�2�{�(�� l�Q���v&=�J�F�g�M�R��r���vxۨ�1Gw&/UV#���JE�m��Ӡ�N���l�Ԗj�Q� �[K+պ):#�=�^e��F�7N�hEA�?2:t����,؎������]Ԯ��0n����r�o�+Sxf��KVZ�)2�N4�����D0��ޓP��N�g����c��~7��em�R���KRԉxg_=��J0G����i��c�Нf�\��^�M�m~Ɗ�qѯM�M���V_=�@�\*"�q�^�����qO=0�*����y<�㵊^�jE��8{�۾w׷]NZ�Ȼ�n@�⌱�~�*���5�Sz��`X!~�ڜjY��=�c�p��s0�bLhq��T
�0���E�����t7p'�]��&$[��I�V%$N����"K�SN�\Œ��KٝPv}[����y��.�a.��'L1KQ��%��X���ߩ�<7Mu_�=;��
��(�b�EOR-#F:-v�^��ϝҩxA��w��(	]7�n+�$o�'=�سi��1y�+�x�|\Ϧ^�X�g2�Aʗ���Eo?\��|g�O��qr������l;Z�6b'��[�k1�K�:��ʙf�P���tZ�织JP��3�v�4e�����9SK6~�n$z�몈� кvj�G�_h�{iP�`��p�����+���]C�U���'��Γ�����)'u$\�CbOS�e������%����J�3��Z<��n:H(=A;���ƺ._Ǚ�k7�A�S]�=O�O�P=�u-q1�)��wW���P�N$�:A���Aଐ�7��;��z��zN|ĒU��W�(����$�n"�_]�T�ߞ+L \�	{�	Ğ�֥�\�@�y$����w��ɷ��}R�GRE"+aY�Am"����BD�Ĵ��PB�T��Y�v���T7k�}�ĥ��1��
F9OlhuU,J��r�9q
�{��;I٤���94��d1�|�U֊�.��I�LQ�b��&�Y�J�)V�)e&�jVBߥy�ٮ��B����_���j��má�.W{�B�R�,Vy_��^�㎎���➇�,��r���5�H��p�P`BIB~����)�)fR/�Pc�ﵔ���FLO�PK�'�W����=�T��sT��v6##��.���,;����~p7�.�hZ�H>�����~IQ�]]
	��}q
�LY7���AP)����#_��LD���&�P�?�ѷ�$�0���+rۺ����(�}Y�D֤@<:���5���r�܇��=� ��,.tm��b|t�k�����Ѧ��ͫ�*�4�N^,���w��3E0���L��RjTm2��og��`q�:�ݿ�F~h'�|W}J?,�9�Ь��B��� ��lF�z{�{:ef���jT@��<<���%����X�XƝ�TZ'��r�/�`�T#��[�w�mW4?�����#��=�����/�\4G��|��ج�mg�,���kg4��_HbevK���;א׾{x����H���Tv@�}=����&�&�zA&l7���ܳ;�ԡ����%LaѨ�.�龓���\��sM �ﮋ���jϔp	�i��v��K�nۨ��=� �4��)���qM�U��l��Ӡ����R��GUaNн�i�z�y�u�a�
�$��ךzs�ꕆ ܮ2��H�'m�MgNk�<�ٔR#�����k�b���{�^d�:}��K�8Y1��ռ��ɉ��	�^�Yj�ڼ�8���i����tJ;�l'��aMa�Q�X�æ��zI�~�Q��pX�C��z���R�k�s$m��P_Ѥ�8F
Xi��T�m��y���pJ�|f��jiϦ��E��&��pA�e���/��s��L�O�8�)^2��g��ic�"�̽,��u�J�w��z��Dr|��d�܋a�N�����pb�p�D�L�n��0П��8��|^h��No�������	�MF1��ڄU�6�t�7�����齌�"��������ۘ&��5iz�����=?xDS\�`��\�F�1i6"�:	��#��C�e�P.��8d�lR-X9��@[=7(�a���vvM���\�h���S�CC�^�x�X@���քτ�G��f�d~����O����vI]m��،P\)��k�)�ٿh�V�.5���>k��W���'�KFl@'��T4��x�0��%n��R�͗�b��M��%L���+�CH�JH�:%�_J hj�(��~=����!�}��+��U��{.qP��k6�Р�ϵ!4�zӻF�"�&B� ����0��w�����ox�p� �M}
Ǆm�ҳ�lu�S�н<9kg����;J�W�7�4Z�>�KE�(F5F�2|j`j���*��d
�(�+�cD���߰E�T�fRe��EjwTu��B�r��ڐ��Є��B�SZe������@ޓD���g^rah^;A¦�=4h�h��>�i=���J����C���L�<:�_Y�il�u/)!)ҹ�^� �}�n�{���VENza{\4?�M=����e�WH�� 8p�ӏb����x�%(��B,�U"�ch�J8Q ۴�����q�W���j绎R�]Ύ,84!��^SDU�ޱL��%yE�^9�Ϩ�U�S�l����_�@����|>kS3��&Rְ�ɨ��lN~]�H&�wH�
�R����Z<j�cQZ�4I����@��Ĺ�v�U�\������q���)��l0|m4�*�f��|[�'''�fĕH9�}:�@���G�D����ņ��.L�!��P��׋A�k��ZZ�<o`]B��=�����w<ӆ�S�K���3A� ���N�
+q�$R�N'��fF�`��/�ZY�FU�|W��Ϥ�jmU����t���C)
�8?/���X��sbV���e7�4���,-�`���O�@0:!@b��9:R "@ݿ�0A�1�ϫ��(�ڵ�x�r�e*2VH�����;����oSR��$�z��C�)�w{	�o�b|���=��z�8/����>Y����@~�~M�5Nr��e��K�~ܑ�c7�5:p�SF?4�e�3�:J���_ڐsv':���	:jX�^��'�ͯ�W�^�s�������d�D
�!�G��Ө�J�[>���&'��$ymm�J�]\Tp�z�.�8NH�0�?��~Z�*Ώ�u�N	u|pOoa����l>�%�S��Q;E�u�$��s-��wobb��B󢌢�'Ү�:�b1@�G׳�L_� ﱎ�����ޘ�;�W0;�A1����P̺uc�/���ź��{�C�uڱ6b�x�������Vp���7@����`�(�\!�E;0�R-�h� �xǲ
�v<� :EsuU������3)pT�+CVA[�;����I�N鮬��d��M�MR�z���^��4�Hg��+dհ�&��m��B'|��w�6%c��l]�*�5�X{R�t:e)����ɹ��U���f�ї֢�g\�]nr뛛��KJuh/Ns����d���u�oڞz��ܣ���1z�MOct(c{���G5���T�I�M/���̀5s]�p�ڋ��h^��-[��%�L $t@4�b� u�iX� ��`��t\�挡�<ll�P���
�ׂO頎=�T;b'�	��KnKI���������|~ }ŢZf��oKa�4ZB����A{�rk�3�U;l�5��B�LW�E?&%�R����5y��lAsy�K���s2?59�Ô���a����/�h��p8��+ڮ.%�#�|�$���035�k�m��w�v_�����ƙ䔬����O��h����,2�e�2����f���^���.�K��}-�Z�����oj�=5��E̤soV��d����ulf%}e��>�C��:�{<��!�;���^�օ�xҥ��;�S-ɵ�8���kF$�ל�2��������{�s`bO�����֝F����h�~i�����g~�gB�Z:iV��Q��@뀤6����������?��]s z'�[\�0��Ⱜҗ<v�LV�j��_�M�o�7|,IdN v9��Չ����'bq�^h���	z�)A���s�1��F�\Ç�%svmg*aR�^�3cS��۠�S�l/�8�I{pN�Z;Q��p�=\v������"��R5����{/I�^�#A>#�;�;_i9 �v&�A���!�W-��?���{eq�����¸	���n�q��_.vMY6B���ꌷV�VH��b�������ʽ0PP?��fS���`��]�0�&t2+$;Lr4�']�1k���i����j�:��sO��(�ϩ��p�}8&%R]xlTm�ǽ�@͔Ζ��/�C���r<�C�֐���&���C�T*�눼���S����e��/Ke@���x�q!��&�o�wR�c�ñ�*��X8&�����׭~��ƮS���玿��8��C��]S�R��@"���r#�������u �NF'8P�,9�A�W'X�v]9�l�H�3��l�D}�l2�����v,"�pg�c~y��-��(��8��஥N���H��9L�7��'(l�P@!���F�����e�����1;��$[��att����w�ϰ�{,�Ĺ&�D�OB�O��cpW��u�4�a�O�zWk�:��x��S�\O�o��h6e�X��$7u��s��è��ʗ��9OȁlԊ�󵴩Ro�%���`N����r�g&��{W����֛6�^>���ƿ��.f��:98=i����x�l\gѶ�į�	$��ݐs?2��Յ���!��x�����#)JXyQ���Uz����0�}i�x�|'U�$j&L��v
�iu-69�{��#���7��;7�\����_aowKl'''q��q��9�����_b��)�� ��.�GR)
�!�o�G�����0�vm5	枎�v}}��$w�l��B_�_q�G}f=�'1��UKg�J���Ma�d�ӓ�q�>��V�',����;� Y�M('�/05V����������G�bb����?�V7�_���ç��?@Aޛ*��Y�(���TxOB� �ّR�������+��F�19uCK3j�w90���X+r�2�L>�����ע���(�NV���i�ώѫ�cee?��5Lg������/��u(@�(?��-��Jå����x��/=l^�ng5r섞�d��%��*��<�����\���	N�:��>'��%i��MO���y���.��GG�D��BM��T;��l�rٔB�yq����!l��%΅B��鵍��m�nU�wM�g]�_�n�b~iB
�.���+-�����1�����;T�=�_�\��e\4�`�Nbea����^�A 1��"k�ƅ����N#�p�g�~�\H�m�	v�bhh1L	
�,
�y�	@/�ք���חqe��a9�Yٟ�2R����!�v��B����0�FW��5��,��z=���fFo^3#�
�+�����95�<���p�޾5t����'��D�Ԝ)\�P6V-f1FJMr����)��ϫW�1?S��;���z���+��X�:�j�d2픊X_�B��T���䩉�ڐ�NY;��an�_�ն�پ��_�K\+bz|@�I��,j���&������[ċ�}��t��W=7	J:Q���&K�ե�A*��w椨ќr��/E�
K���cL>����Y`}k��)�S�+%�sy��VoBeg񌨷b�5?�i��%�"r�]�wc�>�ݏ�%���;�n���l�@ϴ!R,��� Sj]qd��ӦX�Y�T:yd�]��N�d.�EG�ףz-kxw�[��n:���Lw�Y|R�]�����3e39���:7iǪ��i~TO�^JY�9�DV'H��c�.�V�Q +a��4�5�F^�OmFh�Kk��T�����Zk)k�MWՒP�D���RPW�� n"�*�x2���fwN'�Z��#|U�?/��y���E���r��=$�,�wwl�U!�,�}AM�к���E�k���G[܎Y����y�L�GU �VܙQ.���rr���emA�\Ԅ����`�E\!��Ӝx|���M%b�ť�Mr8�r�J�Y��IB�H�K��.�.���k�$KSY�v#<0T��s�0W "z[�^�t�E7�*��F�uE�@4�C�ƼJ���0��M*�]>��iඎ�FNv4��R�QS��(�'����Z�Qr��2oE�۹$�̭��@�r���PzV:�M�t
N�n�_ki�S��+yJ9K<<=�C-��؏&�J������l(qhd}y�6ZJS  Pc����"'�^\];;~6�a�&0.�mA�ݕ9�l}I���j��T��q"aGG���l��V�EF��� �/�&:a�M�//+��"g��c��$X�˱��h�3%r�����],�/��%�
0�(ZG'=:�D	^�ݳ43����r/Y���`_i4u'&W@*�Q�&�)�I_�Bʘ���������z����(��ָp=�P����,f�����>N��pgF'F�3�ؔ��ݤ��{7�Q��^G�}H!P�ve\�Ռ�o�f4ך�8>k��{/%����)+E1���|y���Ɵ+r��w��r�9�ALv�f���7�zm�������<
\��j��>�{�Ņ&w��~�
��!t�&���R@�����(J��"��9�� m�E�wn\��P���6_�jǸs�6f���TP�8�����^����*)��XZ��G-bx�,mZmzH��P%�����~�<���&Ǧ��ǳ��K(�"��pv$�1G��6����प۱N�:��=k�z6�Q� �~�a##|��wp�jk���/~���WfB/��˯���u���oani a�C������<R������s;Q�Sw�[�s���|4n�2߳F�gz�w�&�!����/��ü��s��,K�P�}����f�B��~�+�[I�@���8x�R�H����Q�x��ܭ*�q�.n^��汪��OM��wfqr�%a�lD.Kqq�z?�H�fQ�R%�7�Ȋ�Rq��	vv�1;~�B� �"sQg�r��H�����^l��>��[i)m�7�6���R��Y��-OON��;��>d�O7���+y�ۚ}9��^������bii7�gln��n�
܎_Ǡ0�NT�Ric�CJѶ������Қ�U�K��}-��F�l`2�ʨ����M�b'���SO]5ؖ`��@Y*��ŉ1w��j!?�3�ꩭ�D%i�Y��"�0�:��w�VF%������N$���[ߘ��p��dH�b����m�%GR<fddD~}Nsm�SN�ƥ��b�${����=��K��G@��=2��*�ߗ�ã��X�'Emh�{lv�(�F' ���r�[�r_!���9g�d���U5���P����LN�D�h���-X�,��E�B"lן�˷��SQL�/�ӓBJj/�L�1���3�k�3����U��M:8a���G�1�陏�M-<]+	�1�Ŏ�Yュ��ެb��sy/��u}\)�_=�A)��F$��񢼮�����;9��A��y���mO�"�������!<�&�8���!����ZOUF��vdR>
R<��3��[�z��`�׈�gk|�bV��!���*�x��-�qgǒ����������'��h���9D��AZ�z:i�@Z��8
L�M5�JW�Ǭ��/�Q�� ��P̰��Z�9]���?.�ڴJ⪮Zh#������$W��^����BqK��<[U�`�Ia=,�#����:�-d��|�4�UC�R�T�Kk�+���M���8��/pq~!���5!yv�xo(�8��I�Щ��ށ��P[�R��~����l��(4E�z
7�.%�,̏�Y�#�Mi��P 9*9-�٫
>�j]��y��.2oĝ����Sg�bU����#��Y1:��Ψ�TM}S#5��W�z�q=נI�=uu���^4�^]~�z�pO!j_h��'ER��^��Pr).$�P/K��/队��˙��"+ɔ�@鬏�����.�R><C��
Mu���"V0:Z���8��qtR�Oq
� �JmP`n�a��� ��LJ��ڙ�uJE	���01�Q�}���!i`��)^�����6'� ,�l�C�<-Hu$�G�e� �ݥK�v�U������:������h8.w�c����M^��M^l
�`M%GU�dK���T���2��Py���S�[�X��~)�t�H�	(z�\O�����&G���E_
�jk;�ҔY�������ս0ys�߅b�K��.˗_Upxv�d����r����2�+���(9+_>{��ӆh�]烦�v���`u�,EN@��S9�\��7�����t_��#Ø���r_<\��# ��#Vr���9C]#֊4��b�u�B#	�Yr��81��O
�U�3ޱ4���SZ#F�Q�J.(˻�>��y��5\x�h; gU*�-=��]]�&�>�?K�kWƤ�*`�����\!���R�͌���֛C)�wT��kZ��&T�2�P��*D��,��MI�Q���p8U�6P��ׯt��[�^\��� ����X}�cj��}}6�)vBwF	ji�]f#�4Xď~p��	������lllɽNb��|�q|���⥀�/���bUv�h�6����V��>�[ľ$�Η3=�1P��o���]�;�^�u�Ү�f�)�*�˯�`��qZ����ݚĥw܎l��Y(��M��6J}Y��$P9o��?�{���J"�{������?�����������)���qxQV! Ҽ��jR\5U,*_�I�r.ɮl�,.��p�9<�?��R������#)���\�����[���A^i��o�;�bm�>ϩNWV�0;W��N?������>��=�Kj��{p���a������{��x9�GZ�B�{��&����#��B{,�A�e�)�E�{i;��M�<����qI˟��Dj�Au8O�I:a;�j'�����F�Q�U�N\�g�ծ�2%?�P���}ؑ������pp���+s���J��?�������W��V&��<*gk�q~~���.�U%_Ռn؃�4ÐM���Ǆ��m��?쫕�'��4,�L{*���(��!�]����x�@dWO%�Y���s�.�,���l�>�����J^��_���rG�<�#<�O_<�o>�'���|�e�<PEQ2_�����������#4)ѡ UV鲴��6�\�NK�j��e��<���}m� ��V~�V�U/_�ηIãBc&��U�r��Di�Lܮ���A�����"CQ��)�.+�m�ʐڅ���+<}�&q��O�,a �����N.j�y�],�N�S��Z�;�JcNp������MZ%�j�}$?%�b��+D�J}��(�{�i�R��L�/"�f��%��h��E[E;:��JvT�Ի{�)#�ٌK��j�6�{��O_8��wOp�s*E�>��\]E�����GJ+N��ZԴ��e�gS_߱a"m��5�zJ\r���ܺL�YW����E�wY+�����v��
_� .�a��yT�2��RJ���sH�n7nL0cC�����w���cvf�#9��x��=,.�������u��ڬ��|V����ls�D
f�:����J���tpu���b!��q�U�����4ھ	�)����禟|V��a�|l��Cx�ڤ2�z���6��wߕ;��p��ؑ;Uƍ[W13;��ZՃsm|�� +�4�ȱ��������8�")���-��~< r{g1h1j�N��& \t������w��x�ı��u }|�]"M�Ϸ������^�"�'��פ����!p ϸPJV��BkH�MǧMl���?���&1-�
}Ye�u%���?6ч��`�r�!vw���:88$95�1��Md�Q�c�/�����3��H9���b��P�k�j�lp��g-byy#�}��%��)�.����? �c@�I��ݽ3\P8.������^<�pl�X��j:�r`�v�%~�Fu��`,���é�:�O�(�N*.Ug=?ttԈ��*k^2Oy�m������01�ĭw���i�y�/�nW��h�����k[���$��L�ZF�:���qQ=�??��K3(I���٦�QY4M�۩��~>/�P~���,n_��Y�n��4 ��A�5��M$��8J�bj�w����� �.v^?Ӏ�E��M`�Y9Y|��9d��K�\��$]��Qu�J����%���Ѵ�D#�*N�M&Ն����q��	�=	����w�|z4/��2r �S�?N����t���MU��#����v]<��OHc!t+�����O�`V�����G.Y�������|���?[�C^Q�NS�����[��
��W��7�����8=?FI.���4��!��ЩV
+��K�K�g��O_��&@3�jXJc�m��۾3����{�:�B�:~��k��v���*^�z���u����^�<���i|�ۋ�����ĝ�>G�h�6�
�*⡂7��	����[\�&"��n������))�.W��3�v�
�(�����)��(���r�B
�c���v`� �$Y��Y�/6�A�s����67�[K��[=F!�ĝwo����%��I-`i���	�\�N��q��ML���l�k�BvW��䐇�||C�^_=^�	�+W�r���<�B�
Qv��RܽQB�ą��M�o�)�4��")��.�ji^X0Sň$�?�WI���P
�_��7Z��Cz+�q��3�|�&���p��I�3������וZ�S�����EP�ֵ�H�j8	�� }�NP;��Atʩ�C�@��(V�}_�+rE�	3��M�@ǎ,�U)���eKG��1%_;���
� J�R�d�.w?˺�ђظ��!I����e�FXq���S�c8��R�I����ΐ�7ggX�o?�w�V�����ɺ�+/�يP����2NNN��� "�X�p���Ke�+��J��``d��1�:~$)6U���䬼�N2I���% ^^�QSԟ���Z��;�����1f��I?>�G�s���;����/����o�!���Ϛr	Ȧ�i�vCw(g&J8����ƦJ�#Y@v`�^5���lVwø�sI/S���5A��0j�UJ��i�ZG'�t`�II�yQ�{fe)`�q���X�h2�R5Q
�h��(�miS��)|[@���Y�b	C�N����,.-������!���I^K�z^��T���Т!�����=��v��dO'I,T�9G�لĵ��Q����.��&�d���e�FE%_����f10��R�E.�r(M�ψEG�?�T&�� �$>z�� ����|����70?^ROÜ|���w%Wg�Ͽ������{�2�'�g���Ч�p�2*T���Jl��µ+�8���� ���Sy7r��Wڔܘ5����dw]#M�?U5#�p�j�`��M���eS�*�K(��J�/�����Ҵ�`�B����N��E��𲒓8a�Au^���vL�p`8��{�x��6�ǧg0'�`�͑X�8�8������5�����!�?L�]T+�F���ܣ�7�BZ>�RXz�ֶ���S�U�ǄR��ئ�Р2GZr�kR��1�?K��<7U�es)虩HA0=5�;�ͪB�����'�012�w$�sJ��[ƫϱ��ܗ6n�sS
�I)j�88:W+�(�z���ߪ.�Y�bbltHU�w�w���=Kz�1ƪ��S�W�'q�o|��{fM��UR8QF���3���V�)�R���H+RU-�����o��kz�7+xK�c
���"Ft�Op~v�����t�,w@����|An��hP̡�(c{c��oTl�Bj���^�'�KV�mi G'�r��NlB�.o�n����!��C�G�rJ��жrX��i7��d�+����Ԑ�H��	�v������0XQ������X���rE���sJ[��;V�I�#��Ӿr�����<fp��UV�$�e�RJK26u=��j�лg�[ ��!����;1!u�v�}��J*;�uy�[�i����[%���ٔjr|T0B?.���v*����+XX��*w�Z��g�+èp�GK
��C���k�����m/�T:��hV~_��Tm{r|L�]F1g0�\�X*X���;��7A`�#�5���U��B6g��R1��+#�K�;���k���V������f��(5��HV�`C�ҩ�ye��z�7U�2
M!>2|��V�M��	�(�,=�x!��6frB�n�V��ʔ�e{&&h����7��R!9���uY|�09�#(�T�r �%�/�䁦�Q��~y�w޹�)욭 �c�r����gԈ�?KA.���$=�Ҍ���7��r�>���,��crl����T�$����]����6�~s�%T�rU.^����wTB��JM�r	�|�nߞ���|�_��\�)�E��/�;�U|!+ �o���Υ J�/�4�HyÁ���.���
J��Q&z:r��8E��^�s��*
Gkr=�X���wL�r��(�":_�KJ�M��[��l��1��Jp�ǘ�'*S^��Ĝ����䉀��H��_E����|��7��;s�9;«���&%	�-�I��C����;�5.��sJ��$V�Kdƽ�\Z���s������mI$��vV�KfMB�NBmEK�0�ة�'��M�w�Ty�o�_=|�dbr��ߍ�-����o�����u|��[8;�����z�pb���Y��'�];NZ:]Sy$E�#�9����
u��D6��N�o��zѸ���n���9�3���~����
����OJG0N:�D�n����UI���ĵk�ĥ����y�
W������ ����)ƇK��}7V�ϟ�碴6�a>#ϼ�֮u&H�k�ճ�i��$���_�qz��)��<9S�FM�jO��(����g!G9N���!ȮUC-n΋��l_��G���p
��?�����wn��9&���۫��ŗ����7�%�T�z�	/SBO�OM q�eL]O�DO����,߫|���LF�����P:A�W�)ު�,w��Yc
���wٴ�s;��O����9�f�	���4q��Q�^�qDU�S܍"U;�m&A3�&�1=7����i}'�(ɝ����܄�`T(�%���S4��u�=,,�ꮊz}�y99;ǃ�^H�Iq������<޹����A�\��ȳI���ga[�����8��9�֘u����$/qnz�B5I��W/q~Q���8���?��Q��?��,������I,(��x������X^������M��Q�C�:��g���[K�]��̨��Gu\H,oHv����>?-�a���Nz�\�+s�8�未7�)B�\�1�����n�1���Q��{qm͋�n�ܗ�����3���7*���w$_MK�L�S���~|��ߑ<3��3����DR�{?&g�%��#g}R0�_�p\n�T
��wq,ϸ_
���q̌��27mB#��u5ko*x���7�r3���V*�INP�@��$�#\��#]�����J�|�-�{/�n���5�V����~+W����&�$oShq�F���'���J��o��$W8N��8����<j�6���vX��Ή���T��LyY�.��qs��Pl6A���;Cl���	Nq��G~^
�$�O%UZ�MP���ZZ��Q$�F(@��p�Ew�ϵL�T�v��d��.LO���˗������[J��7#�Wi3PP�V�"��>�
W0Z���ns}�#߫Zk��LJ��]��3(�_sBbw�k5����N��Ή��(Y/�@�?ڪ�M�.���L5�ի7x��+,���w?���� }roJ}9<`��ؓ�<��צ0#?���G���g�1�n/Ե��İ+��re��X���*ӣ���TC�(��qtG�����?�D|����y�ǘ�e�4":
�Q��|=�^/�7m$1�>I1U�MB'Ɯ���)��P�>Z�Ņ䇋&n^����E��Iɣǚ���ک+Gז�1%EV>���/�7�>QQ�Z��1}l|�#��U)�����ؖ���MmR����6N���!�f�cNaH
ҭ�������$>x������c)~J�+��w����c�	��O����}�՛v��&�>ä�&(&qlat c�	���?�@Y
�2�$nz��ȸF5c[��\e��b�-*������S��3ꚏ[3�\��+��}�Q�0l���8T���A]��������rG�u;��_������K��P��ť��s\��SS�=N�|�MdYtۡ�]]Tl�,%��\���AS��{�m����b�XD���FU��v	�m����5��9�����\}��O�j2;}E�Nptp��W��_\���D���C�]e��\>J�
��▌����NBS��_��SE��s�T���PԮ�VK��a��3e&:!=6�U�%a�z�1Јy8�U�	o%J��`��|���%�!Ʊ�j]�������ǻ�'�Z���XZY��k�^�	0�to�П�D7��RR����	T�-�����`�$H
�T$950*�;��An*��U�x�t_%z�0��*T 5�D�a.	���=B5@.�=���;X�:���7����5N�$q�K`,aw_��Wr�j^n���+x��k����jF�� i��J�`G�G���I�`��2�nh&�����R�z��%�]Z�u�<W���E�w�w��Vn}/����ތ+L��y7�Sp�@sjf\��?ï?���QI
˺���}��?��\�~m���=`��3/���CU��A%M�F���P��30Pұ����>2�����PﳖD�~I\�6�.�5�����٩�㵫! UZy\�c>��KܓdW�`�{���٩		�]�^?� ��$��H�||򝛸u�&���7�be�ݱ�g'E}��:pחT5�\;�V։8 ;B|�T�򵹑V�\5���
 7�7I�q�{�cŬ���5[|�/7}#D9�UF�n��P$0a�522�l>��'k���g�^�6'I)�/���K,�� �obxlL��+)�*3}��S<y(_�y�I��� p_7�g%��/�����U�xx. ��
^)'�M����)�7���EHD���I ������t�?WC@�9ff����89i�����|����Ĵ|�� ��S�ٯ�է/�/����>������k�-텵�XN �^�]�{I�*`|0��>�X�]�^UZiB���T�k*U:ŋ\�tj�f+�F1��%� ��3�	[�"��v�±�r�٭��R`S���JJ�n���}����&��_�O��.059�ݭ&�^�aey���-�����&��w��Ohs������s�W2*�c����i"����<��g����ܼv������yqr��&+@�2��W�H��O��.��Tm��O\���3�ۭ��I�:.I��˵U�@L���?���,`rn�++�&�d���\���+R؎���T��Ȯ�R�������O���R(�	��obu�T��C��dK��|F|B��t��?A�Ě�Jw1��G��(��fgpI��r�u�Rl��yO��j���T:�ࣿ�O�%�и+I���>����H�k�R�����=�5���7���/KlL��8@���
�����'��U��6$��}(q�@�ϓ��pqz���I|��J�*���z�S�����<�E����і��).ƺ|b�zk<��I�,beqL�f�g�V���]����cm��b�	�Q�4.sJ|tt������JK?���Q
7��	���)�{=S���c�S!
��x�x��)"y�J˦&A��m��8Eb�D�DYj�{�Q/���>��ɲ��(�������%�\����X]Wp�1Fpϻ�X��������{ߔ�����j����6����e��ծ�;yO�$��HG�'%��*��E�Q�pvʻ|!9�.gdÃE�O󘻒��J��Y�No����ͱ���KPHd�Ϧ�)�0�^����p?�&Kh���(d�x���ȥ���c���Ǖ�Y\�:���ql����2;?"x�[E�V�:e�X���8OQ�d9Iɨ�&)���8<�(n�r2��іS7:G�ʹ^u��,�Uɲ��QN#����:�G��q�ꗁ���tTd#u�N�w��K��{�r����w�!��o
lI!��Ƿ����Eg5��ܵ�$q��2�%FUT��쎸&3�_Rl������KC�X���s}|���j�_�2��n�(aU0�����</�DV�&��40�{ņo^�ӕ�1ŗ��������W/�u�}O�<��ԏ~�{R��h\�.�����S���D}cW�VG�e���cɹ�=65&GR��C�����I�U�pee4�T���U�����M��a����
б
���Ms����u�Sc�G7t�����=��E�$��oN{�c�.�>�_����xږ�sl~��0�j.S�R�p� �;U�$���'SH>3s$Yr��G6EH#}��*w��X���"_��W�(��k!������`~a�E��l6��D�����X	U)6���	���"�04@�b�x�W/���Ś2Ҧ%R��)�Ւɬ�:�y���D���=<\R�����jS}}�R�5�H�7�1�He�r+��نHĹ���K{'C�a�%��S�����-�E�.��x�rO����Čy(R���m|���(Hc d'mu�M����x*�����.�2�P�z_�����ݐ^E���כ��Y��SW�-��g�A6U�Qt�~�vK�ɵ���㠫p����	I��8���O��\�Ux�)๯����~���}�;r�nݘ�Λ2�vj����R�iH���8��/���u9<RDT�ʻOe��S$���ނ���.w-�Ǘ�������;�]��q�Ǥ�q�ul�������{.IZ��jg����E��>L���zZ�	��R����:A��ɒ�����Q9���+�'Q���u�Dߛ�j���n
}�J	hJ�B�C�FШ59$Ϫ!����
{IyV����;a�i[�0�%E-T/���a�\Cr6���o�X�������lD���hꗿ�9~��/0�0-	}�����ž���20+�HiV�z�|I������6�l���uI!i����6�3��7���Ąx���/=g��s�����_?tM�����_�kqƿՋ���YN5#�+��xD�bG����0���	;�$���|��ӖwT=��0?�_�ʴ�̸&�7�GT��z�U��3��˓�.$0&�3*L���'��\�5,l�-S\eG���Z�(m�Dw>���ܔr���{�#9k�������������7�~ޕ����5��+*�0eϥ��!b����zd��ΌO��wJʦT��������������³�)���$ޚג�D:ZlE�©5hb5�S�'�z�{�qQ���=�|��_���6+����(H����i�N���-��|�*Jr7�8W����m���N靻�pk�Ob�����ך�8�*���O�����E<~X���F�O��/��'���>����ǟ������
��앑���rƒhP�QiC�V����1=��Դ�ó�NW9-���$xq~Q���-..�0��U'���z-�t:��a)��Z�+X�'b����ŕ�Y9�"O�p����='���4�~���=�}k���y(ҩ�2�t����b�95�U���������g���/���A�IM����4]�SS�F���[r~s�~}PE%���x 9�輁!ٿ}R�c�k�U�{�LRkc�I<��	�����|]U���я���7���,�^c��F�	�������μTd<��_����k����ŞM]#��i.���o��c?��F�w#��^S�jjjJ��\_X��d
OWO��AOTN���^�K����A���e������
��d�VS{��ϣ�)�#x..��7t�玚���q�����,�h]ynZ%	���~��6a{axY9(e��8���:o�@�>#��X��dB�w�G��|�?��-|����c1�ƣ�k�k�@����|���E�2c�� ���#��{\��F(y6קތ�3�+�����}�]LObk}U�Ϲ��=�&�ϲ�t[bn^
ڲ4�~��12�m��b!��GI��Ǔ�ܩ��|𹾑ر���Q��y6r9���cg����3藸qxz�Q����Ig�g�T�9ƷBN��p�i�b����T�FAGi�<sl�b�o����|�9���7xdE�c��Vh����r��>X�H����KӸBE��O�ѻ��爞�W��Rd�����q��M������DpkGtNb���(�����o�D��R�ݦ��>x��[�huk;[�Z������Ջu���)]�(��{����#8:,+��?}&�4+�����ʏ�Ҁ�h�q'�M��g�GY`�XS�I)x!#糯�������F���r3s�@Z�wT����ל��S�4��P�YO��P��s��+�r~}�TW������u��)���.mJ��h�3�:,�JU[��N�Sq9)�"�Zih.����6E(<s|���|J�ό��+s��;����ݏ�{�#��N[�3�R�fT@JP��*%�]W[]�`�ģ�h$��T���"��ή�a�/�����=���p�\P��
��Ӏ��,Y6����4-�;/_oMpf�㣂wf$V�HΪJq����8&gf�����}�όcD���y哦2q�'M�J��q�=�r)�Lqzt*_+ą�MuK�*�Hx����n���.uc�]{�g���4_�+V1M�`���P�0���K�'v�C�+�(+�'_�
@y�A) J��js1�r��ht.e���]�P���(��c̮�i��S�d�_'C�S��!&FJ(�o*��;g�e� BXB�)��k�%&vr��rn\_�}��s9G������x�j�� >��v��֤�]�xGwb�N8��8�_�[��J[G�E�ߡ,�?��� @�o���fU*�5/�s��X��-���������M�E\X����W�\����k�-c�/�*��%���O&��s�͵-��p�ڲN5�殨o������?�V�/J��C�??�4X�%$	NI��������Y�h����������R^n�\��X�#�=�a���]<|y����\����R�F����ۡ�!tU���\�\6��?Y��Ե�+*����ϰ��:���_�k,_]£���"���[����J/]��'H�VW.ZZ�0}�#�+�{�v�~N����ؖ��/��Yu9��!x�X)mI
�:�1Fed	.4��K���	��|��
)���b�y�)W�"^��\tv�:�<��g�����@6�W��Q�`�ɝ;R�."l��:d�o��:�nڭ�X��`5�w�9�v�|/^�ၼ��׏�q���rF�Q�T��J��uIB���W'���
n��΁��C�"*�=L[i+c�G�p�bUbAY)\FqR����/�Ž��z�:n|��{u� �2��\5���+x�s���O��5>;NE����pM�uf��>��,�'��{�ͽ3->9u�gb���fQd;�6I0bv^�S̋ã�%|}X�5ʶ�@���t���K�0!�c���'XL
h,G��_>V��F�����+W�_���?~&��LE^��sqV�b�^�C�������,�<���(�P;k!�ȡ�)�����-�������I���}�����n$S�5�2-I��uj�o�c����͎Ď�p�>�6P�*d��r_}u"��d8$~�Y���#M�	��� �O/TjnfZb�:LA�s)�C�)��r�2� ��vH����	JEJ/��GY ���$��>��+�j��t�Fob<�����й�ۡi�3�VO;�s�&Ђ�"@d�MQ��S�T�3�h��S6���!��ힿ���?~�����92�=��������ھĒ��Px��&_����4��� Gq�ƻ,z����>�w{Z
4)<�}Ǣ+y���׿�1�~x�*�۞<�q)N�5�^ɹ�甘�G�-�&Q� s7�~�Y����R�����EU��"����l���Gx�lMbeR�^
g�� �v��{yDo.�2�<�]��������]m��% ��̼�׭c�T��Wqvv���]Tj���d���Q���foj���6������~2ih]Ǥ�,j �eB�F�FK�g�*��sG�:����u)�?�pejP��g�X�>�i;���S���
��d�$��P[�1�d&�2��?��՗����arz����D����HNVwv�z�v�����4��D$��I/� ��d�t�E��LL�5Z���g�'�Nn����N9��*^���<59���^��\?|ə�o1�ԧ;�����I?� �_���H�<ը���$tџ͠8n��S��+RX��s0��Hi�f�q6�|m�95J���*�Qt�h3v�Ѩ}���bPK���=�_��O��-��m�m��`W
ݼ���3�~޻�ج]��ĳA�ň���m�6�R8����+�ͰP�-�� ����@�߲�r��_����+��]�ƧJ:}�IB������T["4������urǻ��u2D?�9c��h�k���J��y�-�`^�=lU�54��D<T���d*t���Ǔr���Ȓl�Sδ���Z�,�.���������u�X��f�ngF-�"�������j���C='��3v�s���15���Ҍ������IA�\
�<n����i��+U=-��kEƍ咼�$��v�(I|��i��<��'hiyW�Ƥ8ŉ��i�X��^���ĀF�Hi��TƦ��"!��A�=��cR�v�~��h3�Ob��`/�����/��4;;�>�,����J>�b|rPEo�+���(���ђ��,������Ĺ^?��Q������מy���2�=�����	������ǧ�s^+�����nh�^<H�ZG��W&1=;+�+���E4�]|v�$����#IbZhO��S>и\����~}U		��=�t���:Re�J���"��0#I6e]XNsȩ�t����ڑ�c����%�p�ėE!�a)<gf�A�]�!ڔ$+�v嚎Y��ϰ'��?Ƈ�+ giy�o���p�ĕ����6����M��g��soz��Y�wW;�C$�9C��h�Zi#�P�����ibW�H�1@�����۬J���9����B�FT �κ�5�=�9U	�N+�Y�.�pp�WS�
������9;8����S����Y�u0WB���L�)�=1���l�ʤΕA.;���f��7�\ȴ��ä�8a��#L���z�}k�eۺ�a����$c͞�ڳ��[�����H�.�IfP�c��oY��@���p"GD��ʊ=��e�FǞ<߶���wwӆpO=�:��t2��ʫ�V�[kv�=�W�3N[��(��$�K-�|Үm��Հ�<:�1��{�m�͎5p�8���H,(�OJ��z�D���-��Y�0g�"�$E����ܯ��?@ Mg�KFl���u$g��}����H3-~<� ����T$ԦZ<~Yr�Ɓ����!\4��1���!iT���Tw�5�Y�#䊆U�D8�ãc{�$kn���~#�t^i���^
���vݲل=yzl�^���, �Nfvek�n^Y�?���@�;AEb��ټ}��_�}�v-��
�N����;�߅3k��J��?����]ݚ���K�e��@۟$t��sf4���{8K��E��c�G��m�yZXY���7���$[�Yu{@���Y�֬����,�))L�ф�����&1�:'��acцݎ%��.甀����*8���?m\��m0��v#x7��Ƭ�#m~��k
��#v���k�x�N�*�.艘c$l�<R]W//���a`5K8��f��G Tj��IY�X�o>��L���ܴl!�sUq��.'��O��]$�c?� �ܒ�?�n_��?��9�h���?|�A䅥2eW��8��H(���-&�ٌ+�����=G�i����w�чwq�o�n���/��T"�� %o9\쳳KA娱�>a̾�|3r[Ι�q��  M˖��c8Ŵ}���f�^� ;?Cb:����F��M�a�s�A���~�3����ԛs�b/����������/�w�:�Q`S�UU��)�Ӻ�#9b@�k���yf�ͅ�y[ZZ�>l
;5��� �"M,>��r�~��ϑ�G�����o���Ck�{hK����Z�tϮ�ܸ}OT�$���!�苷��7�:;�f�Y$��a��D��#��rٲ��F�Z]�k1gow^[|P����W����2�cv�`�������H�F�5�)��u��8gd����9-�D¢&I,��"�K�)���{7S��u;��"���@�rv�DY�N=ո�,��ꇾ��uv���;5ᄴ�w�\a5�,�����cgV�7Y�H�"�3���Ͼ��)/���Z�F,���_����"�UI�(�:H�NN�TL��?��ݿ���jH�AB�a��?-�g&+��[n�?���ڍ݇xFO�����wlk�L�ԕ"NƇ,�*l��~����L�ٳ�jkQD�7c��/����ն8?+��O^Yq\43�g/�,�ݞ �O�tO�D����D�Q��?���z�@L�$�+�e��幂b�F�%��F�7Qyb4g($���s)���V��c�tr��KE��=�TtX�z�2Hf㸃��a�JMs�i$pd��ög��K��crv���mϞ#Aޘ�Y��$�h6�?��ث��ӊ��.����	���`���N�rk �z�����+�Si�xv���֟��&�6؉z�'-$�u�CiR���͕3v��&➼��>���Cظ��z�G�.��Od�X���㑨C�p|""�c>'\>���B��Þ�pm��w�������n����R}/!Xv,p��w �A3��Y0mAx!D���X��a^��ֻ~QP�g���={����ϑ����=$Q�6;;o/^���f�#	pig�Hh�s�;ۈ���;O�ve���?��-��V��6���9�ݷ�NB	�_*�ٯ��C�a�	%��\Y(��PA���������B��u:}AQ)=EA[�<�lĜ�%3t���pև�g8cyq����gOI>ׇ0Y�~Dߐ�m�D7�����/�?Ow��=�1~fD�%�o��O���.Mލ�ig�?x�g��e.ng����J�kd(�x�W���83�;w�񵌋V�]$ow�l��k�ޤ=��%������6ח�G��tz����ā��
��|2o��GV�ul��M8�{����	F#o������>�����Y���u��ɌC��'�H�fkx���/#G���g�J*��j�R����v	D���ۆ��ص2�!$Ҡ��E0��ϻ�2geGq�Ͽ}%�A-r���#�~�Quh*�=m�N7Hhj�	�;	R7D���i�b!�-���5�0�sp&�hk��L�/���?��;[6�T�Z+�m\�ݓs�E�>����$SH$\�t���)���m�����?j��d>��O��Yi.k�'�0^:��~��{&_\��w���"{�4Ħ���h�C�%)ysأ�o/���l�N�O�P^���>��#-f-�}xR�~F<;�svj''u�z5k�0���g���dm��� jPz�[�¹���������- �[��f"b#��?w��+N8'5�1TB1e�
	,�t��+ �a^��<kd/u𥸃���x�z��ҶV�>CŸ�/�(x�>���'��*pn~6G�s��-�˫�~Y����)�WG��i�I��-�R�z^�=�$�l��7W$�J��8��T*b-���8�5~,l>�z�p(���1'XN�� {�PN,�O�BZ�֭P*��Ң�sp�}{��b�hI���FS�H�Jv�{�`�AV�)%"�o2�a)]?��U��3��R�Xg4�����HŚ
l�=�{��9��{�±���dډ7�L���L��7s���9
���3��څNϋ���{��m�޷\���H��#1�xl��(�9�������-�@�[vu�v�P\����b�tZI	������X
���i��~���雺��1�@������8%1�{��i&�2�i�6��\Ø��A�Hr�I���]�ܰ��Hp���譍 �P|$�]B���>��,�ٿ��g2�d��^�,&)|K���6�35�qOထP,.&l�x���5��a�Nk}r4(`B�O���� >^8�=l����_"7`��*���a��/�0:�^��)e?�������z��'��$�ޒ�n�JZ�l�fmb���/�S��e�?��|o���b{��5W����/����u�5&�M�U�
��e5��%�=pr=�a�t�S��N�,��4�	;���f�]��LX�XI#e+ö���e����[���Ev�M2���Y��~|�ڣa�~@�IF�aB�7���:i���+��R��n���Ή��;�����iMs���!�?���/x=��O�|��zG�|��L��:�%��=c])�0d0��Sg8@r�e�q��1���g��g��ｱ���,`	3�[&_�1�C��v�����O��"��rϾ|��b�����
ٴ�V"'�NH�Y�ث�C{��{��$7����٥J��uh&�ˉ���"� A>l }�<|f��9��u�������D�K�V���g�������I����]���/�Ч$Dr�c�P,���n�y���������:Ck�vt`�F���.�d�
Y"�ǉ��T�,q�*��H//t��4`%bh2��s`B��	�>A�0TD_=��=c�tD:��5�xya�';�&�i$t�N�NO�q?;��:m$qCe�7�b�H	r��8��=����}����8�ݗ����|W�'ė����c���h��(4��3�E��kWW��p���R�j��Ţ����GʖL�[:;zQ{i������ۏp�9�8�ǝ��b�'���Z�:%�K1�W�c]��<:}��(��ؔ�r:JὋKh[�M7����Wa�yw��>Qᇳ�Lʷ����M��ڇ`̜J�G���ŗ/�=#�sQ<
b4�ܹa�̲�ۼ�f��c���(k���Y�>ei��a��ga��� ��b�!�T_��\̉b��ݛXH|C��L&��晡�d�����!r�$T��QSH6eX8��"Ԏ���`,�3E�W\���W��X%FR)���Q)<���w�g8ߝZO�ӌg���q�~�1酾�]&F=S���4��2�&dO"�p*�=߁����X��������^~h����ߍ#�>��JmlX�_��_��}%*�Y��̸���>��ɪ��ʅ4�H�)�3v�x�9d���*�Ϥ��=>�ı=��.�V =[Y���D �w�
{�*u9�'�A�a��9$�}$�]%��� )���lee޾z�J3Pq/�AZ���]��.	]H���la&guV�|���<[�j��Ȏ)u��M��#U�"�Cf�U��j��Χ8�r�S8�*IQG�ZzX	���4M]������t��Ԥ����O��.W,�C�팥G�B��O��9~f
�`�2�Y9��:���E]������ؒ⛆~qmAY��kmK!1;����#i���&M.V�]jۑq�j�K�sŰ/��p�B�����3��8;ST�H�5uǁ�.ř�b���!�xq�d��Z��a�#���W.�KH&j��$����`;�H!Y��E1�V�U6������)��U�����8MA⢂	
XL�&����nN�L�^����caҽspC�A˞�&&?,h�">g�ꭊD���` �,�!����]�LY��d w�czQebUC�4�_�ٟ+�[
B"VY%|��d���={�v���\�{�/�kB`}1M���/w�����SVׁ6�j%2�2�rЛݜ\\Iq�ZѾ1`���#�s�Vp_�\]Ep�'�N��fK:�d�;9�؍�3�K3���y�!IS�^� ��=��ЎyOG1�`�Ҹ'��3���W�x��y�K|κ�a`��3r�@n>� �T�u��x���;2��L~0�J&PJ�]�iA{E'L(V�H-���/G,�ب���Ƭ�����&�c���Y���l�ç�v��k?�����������c;��T�Ͼ7�z]ŭZ�geؤ?��5+⮼|�mg�g6�숥��0����H��w����y�ډIrV��`�SZ�>�muG٩���HA�����V�<�_��_��ږ]��W�G�q>��=;��y� ܛ�!i$fI'����R{�vE��C�����!F��%	;�p6����`�j�KT6���&rv ���=��&���� ����iE��$ﺇ㉊j�a߂~�f9�Ci�i���ڊo�����.m���v�Nm��� �9���F�z�;������b�|�����_����c��g�������t�h�6�΅Y����X����*lrw�TRKA�º�P�G�&A�^\E��8B���X�ڔ����[=�k�ܿ�i����������������[vx��Y�W�s���}�6+�+��b�,]���!�Ap4L�X�	�,J�.�I�-6��(�K
�z�����Amܨ�ȸ�r7r�/���p�׳az$��.!g��p�s��῅^�&�c�IG[&������8���WmeƷb��y��x�I³|�,�n^����>��U`�Ұ��|F�o��ں����g�;��!�ʕ���/�-X���������ꗒ�htI��"�cqvQ	��,X0Qך�]E7�nR6��j9M^:M�'�m�-��6��U�˾bK�C.��4�i�?��dV4I⭤`�x�L(���O�8D��<;�}D�#H��.� �A >;vQ�#h�i�k�(y����	�$�B��I2t{!$�q ��Лr!LSR���RD��0,�C"�����uq�/.�������\�x��%��C���\Y*����2��ˉ�d�)F��ތ߆�?����Ǚ|Ԇ���q�+�78��s��F,�,�2F�L�f�,����9Ԃ9H2��7�������y��nW��T�Y^ۀ�L�ӗG6a�LB�"���6Y��$a�?A�N�G��ɟ�H:k�0�$T0�8�Pik}�$��� ����ٕ�&3(�A���aB��5�I�Fc������f��'zW+�{�z�k2�)ø���(��@rG��C,A�\���;Cu�cѬl�fi�/�u{�=D����7o�˱�q�s�{����&}<��!�	[6Üc&�b���W��${�F�zdNK��'ʐ�|��I�|RVG�I�	��~uhs8+��K��YŎ���,�Y��sD�L�����wCV���t�]uu>�KG�ISذ{����K��]�D�WMas��\�H���M���mޥ�����=/:v�+�#�.b�j������s���di���T�%'Ȋ�E���'���~�c7�
���h����:=�+ I���yd�ڞ�w���H�v��{��F�U��󕬼y�nBS�͏F\��aе�t�A��c��}^���c�/��κ7������5���ى]^�,����
��Qk�:&�	s�e.��4��jq�T�ܫ��:G -+8�bn�>�p�C΢f�'��[�#i$�Ĕ}S뾧�*�
���!+VS�BWYR'ι:�Wǚ���98��bc ���0���b1eKs?R��KR�p(�$(C<Uą��9�l&�5i��G�������W]��G�=����w�v��c�������O�g5[�GP�o&;��G�5���lB�\�aH�>	�0����h�,�t)o������J�NrQ�����D�.e�(.�g�a�]ȓ��	%���и�䓡�kι�!��0�NxiU�z�e�=���8�2ko�/m�F�;4'h�YY��7�F?	5��dD#!�P2���$0�?��p��⁗ɪ{�N`�'��@$�t�VVV�e�#�D
�[�΅� �
Z#���:nɉ$�y� h|�荵��67�A�A�G`M&�'v���>�o4��s�SQ |�dnO]cVf�p�p��~�DR��:�1���XE�waN�RvZIzhN�]C��|� {�����"Y4;�,׈��QCw���D2)�.�	�G��`����D�SA����K�PVb<��ظ����-xVH���ʼ�^tl{��xn�>E��)N�\h(64_]B&p1�� �s	Z���`U#G}�9����܃X4��N��|ͤE ���'���I�b��}{o���_��޾8���ǿ�lɃ�>���w�S�X)S0r9�y�ʖJI[B��?���q�?�F'�#�g&N�}�J���bд�m˖���[f��!��=E�uF����.���h"ICZ�h
2C(��xl&$d�}�k�{�+$�����?���c���_"��Y�(�	+��	����q��	�Y�'uF�����W�e`1���tt��W�Ɨ� W�8W��l"b�ʡ�O	��|����Th��nSo��9gG#�$�]/5\�+�=��i1��3�j4D�����V���<_Ϟ�ڇ��V4�z�g��o\]GBti�?mG՞e�Y؂k��k�1�	-����g�Vƻ��'�����k�h򷏚����U���������?؍�y�ˏ�B	�xkU���ֳ7G����}�
�E�Wk.r�CD��ъ�D�D�~����U_�a>E]Θ��(Qټ9+$D�a�d]Τ�4�J�ԕ�=�tÇ�uG�߱E�Y��l�<��b�78�^���=�$$��ӗ6q`WV7�����Hj�5ɦGb��C��N�uW��9�>A	�����.�::|��(��N�R��,���e�W`3�I����;[Z����E$�'v{tQi���I5�Y�?�#�o��7�G�֭e�߹MfA��6����q 0��lXA���%m8���i� ���Ն����fTq�0��cL���	�X6v�b��E�K����e�xv﫶t�s{��-�Ĳ�t�P0�����?�8��gw*�,��(�1���@�:�9�<�#�cR3�Q�5���RJ��P�U^[RIe ;�NYd��䈨�g}��_ETp�B������4)��r>�t@�&��]�d����{n/�>�P�����m5;g_�>�\��|nN	[��~$����y;�����X���4e)�|�h[�������+�]��{w��%��S�`~��N�	l|�3�.�8p�6��@=a�L�Cih�������"�d�\���
2��͎��q��lO_j�5K����o�M��J�}=q�I,�c�x2��$�!&��煒#�^��d��wHL|c�.��FLH�C��H��BFf�J�6i��`"y�L�,�<��M��8"�Ս�ΰ�s#[][�+ˈ;���{C��*⿉?��`�����.��h�"��j��5�,l�ڪwi��I�m&L^��#�;?��K!g����<�YK��*t�F���)f4{<�����Ě(� ib"�uM��/G�b5֥�k[�qm��gm�(D�,$q��q'זvm2��q_�xs�s𜖍)I*�(d"�E	��3;�Y��]���
Į�9v�lV�YF�T2)�	�`#G��z*��D^56r��z���-/&��h�s�H�ȼ0�eq��ĸ�h*��ɼ������6?c��<�`6m>��	~ړ�{���Q%S��Ë���g�I8��;h����JmN�Z��d:��ډR�j�Nd6J&pk7���F3)	7`,�q�w�:�� �C@�X�$$�����\Y����(츹�s�@I3�43�'A� B�x�iFdϻ�Z��J��Y]m�9<�x���B\1�㩓փ���܁V�!���##�ί��MA��WX�j�u������}�%u�(��wP���lY�I��R������p58��ĕS�,�}��K$)p^ØU��4��F�0�!r�R9o7n�ڤG:�ֻ6hR�����e� n��u��aHE3yQ����H2�v}a�5�(�ì]��J"ڳn�ewnmY"S�/�h����]<�����������K��f+�VOMDA#Y�$�fk��_Δ�(fl{���1��:�d\d�ʠ���ϋ��RT_�DN��i�)��¹��"۔林3s0/^V���~z	=��ר��d����E��4����W'v��K<�*��W���Y{��;{���J!�5,~�`��y�w��]��i�e���X�j'8'�fIC�F���c�p<XW��R��C�|q����An�F�x�F�v�Ϲu���[��!�����8�v���ƕy{�|��H��rĎ�:;����D�=o����l��W���$�	��ƺ���D�!������U�?��kvS�O
IGO�i	�u�c׽w_U�Y �ǲ<S2�v� �'�2�JL^)+���D2�Ni>#8`��w=�a��R9��7��k�"Ib�«�G�F��B6��ֵ�����\6b���W*�J���`w�.Y�m�_��W��v�y���m$�M�����r��}��bϾ��f���Ɉǳ*T�	�g��:c��x���l���r��ER�gO^C��i�nܼa~� ��3�*yT���OW�v�bSA7�4q����X%�N�!B��:�u:qU�i7b�:H������M��۳��;p���̟x
$i�9�;�J�H�9��P���b� ��P�#��))π��<s��]����ѾX$��3[�莊,���n$�)vFKsV���oNw�5<�+�E{os��?��GV�_�����{��?;@�w����������O�ܴ�����$e�n�?��m������;�GV��':R$�3|�(�����{�A;P� �F'���J��G���*|y������QWL����Q���L�xY�#ZD�R��n}���k��� A�=�_5�Q�:�i8��%$Uݤu��d�|�E�սv�>��A��� �!���aw��m<er�<)u��+x�����~as��A�f�����?��̌�!�{���`_���D"z�"xnO8K���Ͻ�����vec]�	�ђq����)���U��4�5��Ӻ�����;W���T�]��SW��|l/�*��ZDcd�v
�^8�̂&���0��HےH�*@eq'��H�N������ݺ{[:�=�4"G�>�Ǣ�(����%k��YO��8u��0�SG)���Y�c�{3v,�L��'�G��q�w�Ȏ����MIP'����خ�x���Ȟv�&aGIp�p���qd��|�MT<apL�� �eO�m�w���[�0c��>�m���@�8�3��G%/�7���ѩ�{Ķ)�
ּ�<wgq�6V��'M{�r_�����]�GŘN�DR�\�������քm�v��N��&_\&�nԄ6Mg�"bb�T�<L���%��h�s�큋;�Q�fs�~��8�u��b⊈2����.9��#���11S���W7���qW_s�E�a����b�]q�ki�9��ơ�M���3���]�?�<����n��ge{�K),-�X2@,}b�_"�C����i�O��#��(�5q���7%_�Nm��aѤ�UYUg�niaV�Ʊ��\!��6RX��Ec<��x@#?c���#�c��Ms�2�p�"�Laϱby����z�e�k+v�ʆ=z�m=l@�|��Xz��[9��[�H��ۭ~j0�� pgؼ��_y,v�%]�q�$~��|^��l�c�+���(Wb3��Ć	���#�!C��b{-$�r $p��Ě/�lڵ�k��!6�1����C���	��O�`#*��-.���r�.N�����&=k��Io�P;�z0�e\������ܪg�K5�0����d%J���j3S�CH+�ytJC�皛� e_�|��if���{v����Dp&�0��G���^(��|K�	"Q���2]4v!�\�.�rE�ڍ����h_	Ĥ�� 3��r�
�U�6
zv��XY��ꩤ����)$0�p�#�ʉ�,!�Z0����~y� ~����j0�04,l.aC,�8�s^�Ū��
�j�bѪ.����[���gN�a��d-�Ŀ4�`��;<Y���9��(�;��B��h P���pF
jbKe���﷐�pF0�x����/�bGNq^&"���%	��K��bK�v�ֆ��ľ��}�������e[��O��ͥ��	+S�ԫ�9q�P<
��lJ�=���?�Zr��b;x��@]J?�`8W�s$S�{x���)F0b)$�dt	�����gQ�b�4��;�a����//�� ��.���CT,:�c_�pH��������Q߹wUڞ����"1�jم��'$w�O��8&CeO�U�d�Q����:vu�l��Ś���M�#�ܾ��i���	�U!�!4�'�-��K�&?.��M�6�N�,��H3��!�8>=����k����_�1J�3�N��Rb�6��\(�:��)[�q2@J�j̎\F����Ng6���l�^����UK�fl�����Kg�&W�|��� �����i��;�\��p���)q�y����[��%��!BJ+��U���� �-�������?����uE�=n E�2"Bg�̕�=�Z�2qy�)���:�t DP�듌s@�`����Kp:�7��D���rr�c�Q����H/��b��=�H�(2���3�_R3�X!��_����7����w����u��-[�߅=��C��Т*��A���Y��������mv�h��r��)���A|�ؽ��`���2`��5�.h�!"A��t��#��pOB�釄P·�_&�
7Q$�����v�]���{.Aвb�]���*���5nÞv��>3g+�<|&V��S�+���V\�!B���M�[9 (���H�������g�w�	۸���	����m�̐\�����ÈX,����j�<���.��մ͔��wTA0��jY���󴲺f�+kbx��O?W`Z\XD�U��'�L,
2��2},���6r���z8�;�t8�7�N�V�=��!ҳ)��.�nS��˳�$�FmB���ڪY�0o]&��P�\7���qv8�|g3�*һ@X����(�qzZ��pH��mg�U��6��gq�f�_Q?���]�>%��tk8k1���Mp'��zc^o(Mx��z�ݹ���I�j5��a[��w��Zgsޮ�����*�]ۼf[�I����=��l���8�����KO�R:�C�����'�"���+���U����x�g%��(|�p�U��8S�~6�D�ٝ(0�c���6����ceМ�Q؅v2&�zO�Gw|H��mΗ͋O$��"zI��i��G�h�{)��}��w�f* ��ų� ���+��YA�u���&Y
��Ȩ���X�M[Yɪ����`��S�ɕ�A���2�aLD�����gӰ�\��c�!��}�>&��ټ`���hB$:,�w�c�6p=ƃЗ����VjB}�2�L�Wk
F�:qv����x>ӛ�S�9���iᮖq>��{#W�"�"m��ݐ��q�7����3��ŋ!wJ�+ɡ�� 9��I���;v�u�nVP�둊-�s���v5��A8�8q�=�]B*�0�w!� �O�I��4�%=�y$m�nߴ��W߼R<��~k�ᤉ��Ԫ�v�Y)�������#G�D"!��I���	lY�ck+E�"��=Y[�D��̹���?xe�B&���ޛ`5|Ϡ5t����|�ݞH���e��l�$�).pRW����p:�7f���������x�I�X�S��q���A\^��0���;�Bm��N�>ه�Ѥ$�x��D_NO�1��D�8�y�7d$�|��8�j���,*P�vb2���Z�V ���q �JF���z�6֋H.aܚ���_�p�kx�������
YltA�5l�P]>�%6�
)�΂O�4v�4v�I`�h<�-smNf�Q%�Ms�߻�i�sY;�ٵ���o����O��o�g�v���5H�g���Ea����Hk0�P3&�ڙ��	"qd�tYI��
�� �W��e�۟��X1e�R�.&278<t�=��`�d�
'(?-\��_������n~��Hr;}U�w�:���muu~��ODZ�O�B�]�٥%��Ҭ$&�Q<[��F���.*)�ُoj�n{�����Y����;�N�n_���1���]HEK�j��*�0������ �R�y��yɼ�ꖒ1^��P��%��*ba�&!䁖NSi�V�XϒyǄ��jPA�b?$����R�:~/����_�cLSwB���X�=�E�����e2��a�!8���R��f����k\<�(S%t�N0�M��jF�xm�?�+�֙
Yc�0���g�=��	R�_`-:��?���gJ��w��ѣo�\Z[)@��_3�^<��W�������k�I�Xmn%����9�ؗ߾�<��ζ<=����6������9�g_4ڷ>��÷C���7vp�ts,d,��'ġ;�!�aB0��}Rh�No�N/�$�I	������9����>G¤\��#f��q��w�LGa���u���5[�?�*#��IT�u�M�܊�$@�2��l77�g�U�ݢ1� >?��S^� o4��f�.//-us���&ZEC"'r�ڔq4��M�Z4���ڃ���b�>��=�quŚ���W�
^��{_��rg�đ΃]���G?���/����E�%$�d���7/��Z�F6W��/��׶�˸���|ƤѱGO�lg��A�Z�@ZJL2Ȝ�f����a'ۏ2�Kt��0s�E{����.��h��Ols}��K)��W�ا_|g�N�V7f�n��#�>?��ʮ2=�_PT̂a�0����2�fg#�k
�E��lg��W+[*�-��=�����
��5%��):�9A�b�\����S���T�f��W�(.4@���t�6�<ݾ�n[WI~�v߳�ܬ}��O���jw�l!h����|��B1	_wϮ!X��`)����o���c;G�TaG߻���ٯ~l�6c�P����{f/�T�=�����b��Ȝ,��PyR[�P @��%���L�8KM�<��cɄf־��K��<�>o�T���N���g��H_"�]�3Eu����쎥Օc�T�i8�!qJ�#ѰC�n��'�������zs.�5S˩�+��lc��k��G��1����Jz!��$	�������>:ɐXXw�'7߉�a�>�6`��$-7�o�ݛ���CRŹ���N[g�XH#��/�8S=�I�<̊�5���d��D3�G'#�G���x���+v�ƺ�/�,��.$B{��ǔ#q�e�.��C�(w�3��e�(�R��O
Ŝ�O�fG���@�l������}�y�ƊK+b�&����+V.��ŘI��	D=�@$��!�^0r�RbGvp6uR�Ɇ���� ��J�p��ݰ#$�q���pԍM�Ɔ������rS�� �I��`sRm���:MuX�Vn��F	�.g]&հA��Ć�-͖ŬIHa�h��P��,���̖&`�q��#����F�R��>����|q�ѳ�gGJ�����up���`8VQx�f6�qQ���.�{�����/1�E��� �Ǐ^ً�6�sE��차��q�h�	p�8��L%U�1���t�Mk�nΐ�}Y`1�ri�g��$��;��X��l|چ�ڀ�#Q+,���"�����)��M�оkV��خf�LzĎ �FB��T�?'MI��
�B>��2q����%��6nd��֬�����ǟ|(��&��J��\��ٓg����J�_���I�f��w�=�	�]X��t����uCZ���e�u�����������V�wEx6D���eb�}!�5�K�y{ �8��		v�!�2���w��)����Ō*�QYF�^G����gA!��1��Q�a���g�W]\BU���_��(�
d�T��K�mb��c�4���8�2g�ȖU�<�f�aKpw�A߼xi������f��CUji�3�k#���g_��R�|p�6�����:�/V8�.�p8GV�pޢb���S[��޷r.�ڱ�۷�����[ĜWƪv��c��Ga5�sø�D���	�'��%T1��R���y�"F�)L]qU�b̸I��l�^��8@&b����e��=V��A[��b�ù��e�{$Ǚ_�b���v~qi�:��x��c��VH��ȓ��M?dh��N�0H�����(���[�K̈́�؋\��k+����խrQ�daN̬�Å�ǖ�g��ڳW�m�Uϖ�2V�&����f� �]��e�ֿ��$�A�ě#k$�vgcӒÈ��U+�a� 1,����˦!�P�'���
B1��=�WE1�<������aێ�Z�_��/a�e�=o���:w$�!�,�U�&�m4Q�i�D�z��/�d�'
 ��"UG�2rA�C@�,!p���;�'m�ն54��%�I�0RU'&2 B'�KN�����ʉ�XG��w��1%���	�.�܆������p���h��E�1��p�؆��a�����墌���\\����ve�?�۝��WkH�0Fi숶	Ep���a��$K�恵�Kf�����{�#C%�%��#�ut�u�_ԣ>��ƭ��.����{
V���u/�לk�Z1���%�!+d�0��&�c/�+񕁃��spX������:M��ΐ�Bͤ桢����.�q?WmЪ��6}tL:V
�7�Ic���Y��B�9r��\ �vC��
G��tF�@?�����Z��n���������������
���O��ք�I$�6G���[���y�`O���+u;?����1Rǒ�����W]�3�t��9��L���~6 �-�KF&�,`l��:��Q.��������VkL�T���4��3�kVlq�1������,!9�#p�&����*�;��y�kv�Q�]9�3lF8�7q,��;�����#!>��	d���{�F	�v���>�&�	�D��хB�L�v�
Lؽ��KH�2zO��]Clk���%����Ϻ����7����'�|l��wWq��"�؟��(6)�|��'�(�`��#;�~k��ó�H[&b�!Cu1�C�S������K;;a�N�D�P��l_	?!D~�\�<=-��zJ�.%)0?WVg����v����]k�SZ�����>:�����U̦|y� a6Q5#�/��D��)p�~��X�c�`�~$��5��ND� .P��{m�̤�<�9���V���Z,�S+�?�H9��DA��f�̦��I"���f��!�%��ceW�p���_Yزo��g�v��k�N�VWK��_|d�uv&�8�IP����]_����S�
��X�k��F{*t����J//����f4~щJj����g/a�ag�9ؾɖPf��
�;d�e�A2ޅ.�=�+2Lz��������6�l1٢�N�O.��çV���I axO�D�0�i6$�ǀd��u\��.5��=rI�l(3 ��\A�n���kM�ա��vc}�z�d�+�SrOp��Z����Mu?���G:���\v��P
$�
����!�[c�B��;�lk#k�>�Sʮ��Zy�lW6��6�#�6�(ǜb�-,���e݉㳦��Q�Ge2D2��n�״b�(��:�'�-�Lp����K�e�YK�RjVh�Ā2�G���x�\�'3JI�¤���>�G2Q`h&�`v��%���-�&�	;�C5H�Kǖ;����H�(i��w�wŏ��qg��?����l�DSq��tť�Mbfo�Lr>�Lk�3ȟgrKR(�o޴+������`���8���g�~���Igmmy���gE�Vm�q^}�0ƛ�{�������ɸ��:�,�P����l�I&�r�g�Depb*b5�Zh�p�I<c�������QJl2�3_�#GG]ة>��(��T,��+�o�:B�L�����DryX�ˎ�T�ׄOW��d��!1�Cj�.�Ѵ)K2��&��`AM�Ns9��w����N�0p�*t�F*����,:G��\��zd�s�[�ę5^\�Y�kY1=k��9�`1:�s;;��{��Y�䰂l����'O�L,���7��+pֻ���l�n�(c��2�����ݷ�pVd���$J%��Z@p���7v6�j�����I�<�R�ð!��uits�r5vU�f��˔��R����~n��l|_�8��Ic��f���𰊥t���IG�������sxb:ґ���Jp�T�Չt�&��%8o�i���G���I����	β���0T�
�h���O2�(u��9v#a��u�8���r�`���dC�4Ҡ�@s-�\���Ɋ�%��=��4��e����-�.�����t�\�Ե���\\\��Ō�͗���>��{#������{�-��r6u�9F)?�b;�4B�J��;�:��av�-���,,��ƲT����v��,O�3�I�t�|���_�e�<��u�9��ge.���<�{=;�����/h�-��x�(��HX7g-B=���eeF�
��	8��.	��
��Ś���7���	L� G0����ݰ��%lԫu�Y��2����b`��6Z2���e�%[Z[��\ڮ���\�\�z�j�>;�}�+�(�Rv����ꂥrq$W�օ1�;m��G'�wA��H�4A�#QQ3���NBV[Q5�<3IUȪ�5	������ϧpVe��鳧���6�6�IF2��`��II���2��߸wE���EIc�9M�{��
q/9���~œ8Ϥ�������N��b�j+�?њY}`}B�|�I�BQ$�$��IT�xU�E��N��Q���$!�|<r���
-/-��Ƃ�`?�yxhϞ>���8�����}��-���wP��/ފ�3{zZoث�8�loUL��fW��d,BS��:�������H�N�p�%>gd�ܢ���I�/�b׈�^m�<r]P��q�ig�i׷fmn.o��i(}x�Gp�E{��"f���_�����O_���x�f��."��X��SJ�N�iu��뚈
�QbFI>�/�{�$~��Ax���fΟ�e�Z�8++�E�vR�C`G�)(`b��3�~$���,��Q�?���Θ�C��T���g1*U���B��'����G���=�����5o᳑��!�k'Hh(}�����s9�˳k��أ�:�q~���YT�=�%��O����6�l|/�u*���)In�zw$�i�[��D�Y�H�s�|_!D�����Yk�����L?<{"
���	�����44�֝[��y��߱�%�I���<�Nr��	ΐ����w1��2ϑ19>� ���R��`ޗ�b��=��}0��DZ~`���9��S���>�P$��o
"�=O���<>���r8.�ؙ��΋X�O(H����U$V��=��=��!|J�~�˟ه?�"��ٙg�^�Y�	[�)�9���b*�������e�V�
�Q2��=$ʃ�BI|�6lg�P6�Z�D��y1�8��Kt��
�~0�q̇D��l�m}e�J3%ܯ�>�Bڥ쬓�"'b������ޑ�"�e��� �����"�2����V-�_�9Uх���2�&rJ�Us3�P[��I��>�A�k�N�"�E��^Q������(��&�O����<����t�~�H�x�x�I��/Qf�9	�T���q��D��MrF�I��(-��Iw��ϸYT�#J��D��@<�?��b�h�3�#�=Z�/�BJ:���4m���ܐʲ�o�3F���,jaJڙ��\"F����Y)���fՖ��lu�,��'�^�۶������ή�U/e��Y�̒�w(��H��Ӟ;K�F9�������༲!2%�F�D�B�S����@�B��i��R�	��v(�!����^r0��i�v⊤$���w�@N_�ל��$��Kke�ZI��܌
[�vShÛ7֬��h�+����D${I[�O����,b�$c��@�M��vz����1�.�v�o��g4?������Y��R�=C_���P�ǚX8���8����(�A��$�'�?���G�4S�ߍ���'v|zj�;�	Őy�6b���Nh#E�'�G�&��Y!�A�n}����xA<W�
��4+�r>���}gr���m�c�ԓ 3	u=���+?`�!:�	M���2y%,R*�C��ly!m�9��b�/'m����1jKHKH�����d����[ë�k�� UN���j!NOj���ٚ(����[7o���W$���8���?���{Mll(-�1�8������R�aia!+(@	J�u~~��E`���Ɗ��0��_�Ѷp�����9��n/<[�Z��$Ŕ�`���&�ꨅ(6%2�S��P��� ��IAX��}��x��V�ឳ��uP�a��iԽ+̙.��)��dzݗ0��@sLc�4�{�`�mX���bi��O�����?z�j�u�yg��#�:4.�vum��*Z�~�4g�Qۆ~֞�>�7{��3��Śg�~��U�y�d1l��Y�N��v|شݣS�[F1�x�� ��AVb�=QZ�=���¡�s9����+��+\�[�8�9����E�ۛQ�j@�����c�������֚C�^؏{�����j�8�験�\��L� g�Hc���	̤��V�X��`��w���E��Q~��M�G�u�w_S{>M(�K���������,ms�d�o-���Uu��"Ь�۶��l�]Y��t����5+M� ���ظb7�>�Z"�&�Z��ӗ�vpZ}:����^ݰ_��&��={vi'kT{��͞u9�,�Y؇��|r�d�B���ٴ]�Gvz�`�v	D��_�6F�M����������}8r�i$q$�t��2����A�s1	'�,�;?����������GTCIv��P�@s�.X�S��4�pokE��?�@"=���*�#7��}IG]Ň��#��`<~w��C��&��NΪ�j�?����w%6������o�|D��cTB���������rֶ�#���4�1���c�'I�в\	��$sڏ�/�4��c[_[���u�$������`4J����l&�U?�!xϤg�}qb�����؃�����_T4�re�j���������H�"��s����2�ub�g�n֋l��(�-�:��]p��"�w�7g�I	� j�@�=��+h�<K��������  -��X�ߑqy�7���7,b�p�����NJ����xA�+J��!qm/w�"!���ԶO�zm_}���u���HW7q�;;�Z��7T�%�u��`��D�o�I�j8��%�E�w/mo�D4�s�6��_�ɚj��6̓��$��fn���t쳂mZ;�dm�^e��ݸQ�������SuF�儽}�c�_����K�Ŭ]oMs��ɛwn�����AϪ�-AD��*%�]���@�9�`ԘBbz'��F]�Ix�n%
v�Z�$N�,X�=��������K$�:�!�V� ����աg���p&͂�<�^]A��%_V|��ra�ۯ�Z�C�}����olv�����e��{�N�8�Ȥ�n��d#o	����!:kN6B]���۽$+oU|�?�����])�{��9����;�7�2S$�����
�k�w�m������o�ҙ=z�D��߻�y��`G��TrV���QU��xߗS���\rL����L�C�nV*꺁�H�:x7I+l:7jRb����l�N�F$���B�DB9��%��<�sU�P�@�T?L
5�kF�e+�n�[��Hv��O֪Y�z&tO<����/D �$�|L&a��Q�N�~�]�dy�D�+/�=66�{��P���B�xt.ĳO��dZ�z���n.X�{�3�G:8$㇄%2Y����o˳����d�o�-����b��W��������~c}�����v𽫖�E�_;�R/�H8��$�������]."�dF� $n8sǛ��;v@����9����5��lφ$���Б�ŋ+�s��S;9���MqW�9D����2	����#�f�v��5[��Z	�ӧ۲q��޲�[W-JĎN�V�u�d��J�6����gVl�L�fR����"�Z#>Lg
jZUqO���H2��s�I�,ӄUfvU�0)dl�&��^/�}��K �>��O>YS*]G?+_$��N�̧�:lV0ɟ��ܭq��}�\a-�GB4��q�Rw��9�m,~ �g�嗼.q<{1����Տ�B�y	ύ���L��v�|QV�|���b4&�*.��ڒ�.�lk1m��K$r/mii�~�p԰E2��" ��;�����-���D5� �a7kȄ����L4��5a@;v��-��_o�g�:5�d<��;��F�"����������� �:�:��!��K������/.�-:��Λ]+��~� �6}���͎X����g�V�y
�ƽ� �\t��{�&V�9��#c!E,K�N�(숐Z^�n�8��ʲ���XN;� �PRf�o-[�ޡ��S���#��ZX��x��91���;�pn��(U�%&?��Xz캓<D��,����ۀ�������ݳv�gY��\�\�����=�g�f[mr�ߦ�e+Ζ�,���վ:՚��f�`�3����c'a�rw�bgg=�]��D��2�f�ʟL��$б$b�Jź$�o���@z���Yi1�rMVI�2���Up��X��k�-�/ڟ�}�5h¾5\�T�yVi��"����:S1s�ϸD�@H�7%�p�
)/�(���r��s�x칪O�j�D�HG0�^�6tc}ގIo]�s$c�\�gX���\��ʅ3���0���t�{�Te��0f�|�ݺV��gO�᳷�>���l�o���|�=�ڗ�!�k�-��N!،�8e1{�S�����i��m)�̫3L8%	ڭ�=}vn�0�o_�P��i�(HARG2�w��x�98.�"Q$¬�� Ѥ#�[����y6[�$�d��ˇ��{��;�[��O���.ZF3V*$���R1��A$�����M��Z<<�;�������"F�i�v������H$�ȋ��\N��$��DH�����~��8<Y��s�@���fu�v���}#�P�뫒O�`"g
�j9�*lLh�TRw7�N�¼�X�f�*�jy.�;�h�eo�H���H"�9�J1�����@Z] i���p��2���H	7�Cȼ?
��s��S�Ιl�+1��~7/vRi¶����-����vB���@�:���eATҖV���	�6Sް�y�=��E���YR���b'�"hXT�J�w���Q�3�y��%lTi�yzvo�OA���}Y�E{ڮ����)H��q�@(�����텉>�`�*�"�MY\��q��y6��L��GU���5�@C�k�H�hE)���C�|�`�}�K�c@�,V��	6f��W�6����\2��A��~K�˔�!�e���Eӻ�ϒ,���qi'����1��{�������m���]�{{Ξ?^A ��h�i�+k��;f
����"@ ���Ҭ͗����}Mm�Y���s������+ ��:! ���ϱ�X��c��	-��|0�g���77�S�r����J��C�@+s3����W/$Vsz���B�sp�)�F̢^(��w���}
?ԵN�B���L^Z�'H�^a��H���-���z�&ɲ�:�ZG�֙�Y*K����#1C`i��K���q?�w�ɵ]rͰp9�� ��鞮�.-�RT�V�"���֏���z؃D��������s�d�Ɣ��	�V7�c�����r��o�^�"�g���2�Q����d�Bޜ����P���{C�42�aO)q�g9�\�n�)��@��ELM�11����:&ǯ�����bms�xK�`bf�>��^�摑=��{���a�5�<����p���1�����=��<[}�6[h*]�x	g�e?��,H�մ=��籫�P�����?K��p�F�ۊ�Ue������wX���Ue�0��$��"����ru��o�y��J���I���(C9~^O�1��-P��4�ڰH�{��d"�LR=9��}��Z�N���2�<۶Ѩ̛�$qt��d���I��N`d���ɑ�EUN��v�~��;ɸ*H2�]��(�#��p6.�PO�D��C�N(�hB������m�f^�%S;�i��ER>Y,%�Q��b�॔$:�tT�ݨd�<6�S%Q��ŷM3���Lj|P�s��Œ�ͫ�x|P���9�$�q}#�;(O�O�U�����b����w�d�*:r~~&{��	a�(�8�H��^�r�!�G-�;,��E3j���o,�a��ȉ!dsU��ύ�z�ZC�	��8����ajRο<�����g����=Y�bP.����*���w,���+�����Q����j�w�5�`����==3������3��Ϸ�O!��GU93��ѣ��4�[ԖΜ���GM�41�1����PA���l;;El�\���>�8���yY�1�clmհ�w��	M�s�����2V6^�@���Ӓv}��$M�3	�rI�%��Z!ll�c��X��TF�u�G䠦i$� AyϪ�q�4�
�Vg׏�X�K����h�oޠ]�"34�La�L2��0=3�w߽�G�W����[v87�L����I]��0��) �mik޷C���ak���lE�f�}~�l>3;�@ɋ2J�&�<���Oprt��$��<0��i~gD�֠�t�L�?H����Fu���PL��u:���ߐ�f�H@���z꭭oʿ��9X�9��v,	mVAQ9�4���݆����ճ��}�hN���f�Ri,�v�{ؓd�Xia�ذ��<��"����k��1�,v<�*��/NId_�׳�
@����"�� ���������;J�����X��ƫ�5������!�k]�M�
q)$���*���TviAҭCɟT��|�R��4i�����ֺ�I�H�I�
�Q�N`�L�&9+�i�ɥ�_:Й~�$"�����/���1��g� ���̺��|�8�Gz��=Og��>����$�Y��0МG�I��/�e�L^� �~b5	`%q\�ⰸ�t��$jQ	J�xD�%��/@[���7��x�����p��+c���C��j��:uĔZ�v�ۆ�C�p/��Dr\.�s��ڸ0;��ז��?����X~g_���>~!��9���_���Q<�l�O1�0���q���p��T���܄v�T���@��!�h<���7�(�D6La���-�:��Q���*��n��o��q�=I��8�b�͖Ğ�����Yd
�(AJ�J����Z*������8��i�jPe�V���(n^���lHŐ��H�"�pT�AҙحGi�� ����b	C��e/Ix8�b�\�����5�C��!�1����G�h��$����xA%KW��|}/_�Ȟ�FadZ���Ŏ�R��+��θ��I��pV9��G�����������o<y���>���$����˷.a� x��	������[�<D$Y�='�>�B��&��:�����QM>�Jo$0hKR���!�:�r�Fu�"k��bUY�R��*�,�p�9�'4.����ɑ^n��%�7g�40V�r(�]~=9��au=��E*S�f���)��1c�ԕ$;��U�b���*�6L}�i]'����3Tk]������N%��^N$�Z��n&�N��H��W3��Q�8���׵���gx���sp��\�����������^�4'f'�Un�@�E�4O��Ȱ&�w�>�����?�;/�����O?��9���F������*nݼ��>Y�Q����>��ڜ�r`�JL"EJ���^ӓXh�[�͞R��R�!o`��^q-ߨv�r��]��������&; 0��|FLrg�GPl��6,a��iR�E��*���xS�X4�s�E�U�TD�|qI���ܼ$��|� ƹ�T*6>4$�Z� �2f�c(���*�-&֒�y�H����#��	0N&С�
��������^*��$��%�&�"���`[p��c��ĪӐg��"պ���j4OsC����hy�[{x��n�\���#IN��157���C��M!Q��*��U)bi�"�Ʋ8���OM�;H=�������q���.%�ԑ`B����O@-��]��j�e,��?���wř5_�~��J�7�ˣ� -�6w�$���
wt���+!��k*�&��Ѐ��J��o��]�CI�}�Z���H*����zB�n�A6��BE�$��F�C�$i����"��I�#Q��b5f��}�]�Q��$-� S�rzz�Shu����e�K�3��y��Z��*X�o�|%����WW�q��nܸ��O���&{$'	_Z�L#9y���ΰx������-��(U4���G
�������}�5"#\;��;V�_��8��\�$����Q�pXoy-L��cwP0!u#�i5�]Nڰ�T��~Z8���\`��&/^�ǄU�t}c4(1 �y�6�u�$%	1#ˎ���3�%Z�q�����&YNuYz�Ai��İyLzÁz���S��YV*��}K�}�{Qꆰ�̄��S�]�Bء�W�TYI(��19��tǻ�Q�at4������|�Dzt�¨ܭ:��䧆t&�XW<a���z>i�ϩoF�0E��t�C����X��w��1aU�
����}C-��X�ɧ�<ڙȾ�)�[�Bb Ꝅ�aO[�F1M���͹���"v��p" ����*���Z��r�#U����z`��J�|۔�ZD�TQ^���rqi��lX���+�{����3y MIKp��Piվ�QV(��v�)s��T�T����ǩ�Fc�f���=�����ݫ���?��o�j�%n���}��,�v�w��8/�?�^4mv�dg�U�\��k6zı�K���¡T�����j��(-���]��z���n��#������8Y1Q5������.��Aہ���X�a��x%�F)��9C٦��}��H0<�M��r��m`�ʉ<M4��
k���Y��rK��_�'�9�L��pԴ�];�O�yǬ�4�rA'Hg�	�D�ESO��N��*y��p���7P��p4#{�L���{oX����F�P	٬�ͭ�$�js15���Scr�$����?�L�YO��
  ���O˿���#Ϲ��0V#���N@W	�&��ɯ������vjm�:�T��A<�8G�B%�̶��:��_��A���U��\����V��w^����<�ѣ�����u�]�vl�R�?v��jՖ�iI�#�Q5Z��VVx��D^�c`�>:=��4j�>)��Y+��X#�*���|N�=�^]�C�x�Ǉx��._^ƕ�p���Zug���s�`�v�h�ݥ	���k�#���T��'M;��]�����X	y=+�U�Ү�[��*N�m9t�`	*j�3�!5�5ɘv��U�^ja�Qd�,�YD�lx�"c�O�FJ������7?ס8���S���ČR��l����Q����EQ)Q�1��|�HǄ��
-�%�w�^#O�ƙE� 0vPk�s�ت� ��{����x�����bc�X��P���o���.��N�g�l4%�DRgz�l����f�̮����_��ze?���:���o����W/,`��v�vT���������wZ��BI-v)K�7�C%��YQ���n�g?�ɱ�gQ#Ǩ��Nر�r�V��/K�d��F�h��[uU�a�F!T�*X����\0ΆrVF���F(C��@JPR�.\�DmT��E��#�rT����c�<��c�4&f�����t�?�����i���Q�"g>:��f���]4�l���O�`v.���O?�%��͍�h%�\��/>�W��+GHd��E����a�����Z��'`���
���/~v���O��G����{�T����;I��w��翼��$����T$� P�J�-Ț���N���x�4�Ӈ�35�0�c��<� ��B�g�0���� �*[�z�#;��S����fج����8�55lG�BTY'�*!�1�
}ÿPP���I5�n�����&�ɔ���쪇G�P����=_~�F@��i��Ιs���W��f�P�UU�(&f%�%�{�]z{x��Ί�HI����{Hg�8<�b�́$�5�"s�� �%���m�ϊƒ*G_��c����,.����En��V��ˇ��i�'Ϟ`���G�#�-��Ow%і5I�U�X��=K�g�޵J�p,y����v^U����$׬��!eS�������I���)�M�#�&%���9�&�2����g|��l�IO&��(�׮�/g���T�yr,#�wH})�E�F/;��OMIҪMLϣ��}O{*���e�O�,T�1��,�~4	`l�k�aX(�~��>�3}lt�p~��q\^�������e�h�
G-����H��Np<���������y\�4&��E�=����S
�<�����-Fp��-?���*�ͩ�{�!
4�	m��z�=�N��s��6�4x�uQ���Ֆ�^��0���)�$�C�8vI6�� Ga���!�
S53�,_���2�Ȫ�`Lk1y�8z�:��p�C^J
v�ͪ�����R7SCC:�������(7Ԡ[�Qh7�o�N�Jބ��$"���d�(��r������1M���h;�f#*�m�C�z���j�m,U�yI���B�x��/)�%�է=�(�}�V^����Ǒ��Z��L�@�b4j�O���b�#ۉle8���_ձyY�c1��v��Pug��[���XTK�ؕ�8�k�b$?��S[.�5�4C@vi~Պ ?xON�$X�+8/��K�G2(�wpx�F[K	Qًi���N�me37$	 h"5�EJ)��`�J�l�v�s~��I�B�%���#���6��,8y�v��7�#F�BC���=����@c(�� �I��^���1vv� ����$�Uـy,]�&I��<������B:�*���ch N �뙄�(z���X�:����o�m��U�\.-I�(��k���Y�v�α��[�	�A�H@;A�ta��x�,d2j�pn:�ѡ�\��}��Q�n���D�Z�88�j�=Ijw�@1&���IRLp��3QK�b�6� ������΢�.i�W�Rq0%�[UU/��"ߛA����3<hZ��v�B�vwN����̔\b�_�û��TR:���$��O��D�x,�)���$�8ؗK��SN^~�\�	�ϵV[�wG+;�̜C�&wƾ#0I~����pa��3N�ң�V]�_�&�'����A,f�ֺ��[�� ��~:� �0����������O���O*���lY�T_���F�'����ȺEH�T�\R[��a�`�F���oat�����z�mn������$��r�!��)�N��:CNB^^TI�N/���}��Z�3���٪���|��4>��:^=}���"���(�,��loV�pv����W�,��w��S��?"�V�&�������2+[,F���d���'Z�	�D��L^�1������W��j����CER5��4�b��*�"�\7_����C;��dB&��x�g���;G@�y����>������=E�0�j��Xg�Qԫ{X�v�	��ʚ�ݶI4��������D�&Ō�=v�%nIޠ��KrV�f���=� g�`w�ۿ�K\]Z��Y[U )�Ҕ8LO+UWzJO���yQln�˯����p���(��|��%"���%�����>��/qa:���aW;bL&H���y����[�����h�b�W	�����~5&�W�=dq۪���¸��� ����YoV��Ҳ�Ѕ���VV.?�}P= �ew%�Q%�~�T�4�g�Z��kr7ʾ�G�L=������ͫX��(�ۈ�k�0���"�"�r��n�"hs 1�)�J���^�`nn������W1���J��.����Or�P�L���:$����氰�uN�Dwo�9
)���H�>��;�����Ȝ���i���`x,�?~���k��Gu�EI�T�a�����k:�n0�k�m��I��$3����R�F�L>{z	j��3d���I#(㫨���B���[�	Ba��	�"	��	��T�H}պrG�H����2!�QB��3���� �Q�J��$�;7x����c�Y�ع&9�Gg�X�b��dR �<�>z��$'G�����4v���Z�bh���:�v��kf��|ʹ�ʢY�������<n߾�/^��GU�Z���MI[�����Q�m�T�(��h��F&B,2���=;p��x`��q����}f�ʳ2�Z ��Mԃ�|&��2#�NJ����m��"	ӱjw����\�A�JqC(�tM��ºw��\�g-ܻ���Q99����X6Z���nm��Q)����Fc	����S�ca~��U9���F )ԉ�e�����瘝��!�����؝QurG����<o4R�n�t���u�`��,$���l!����`G��$C��YF~hX�pY�(�F�.���x	
�z�����/�W�P�	S�1Z��>s�,�)��p�-F1קb_�70�sz�~�c�Ƅ2�|s�^��ՠ��b�g��(�5*�����ǌ# �_��	Iz�����a������z�&������+h�
(:�+�,���6yN�%4$��]Z�\���3�ZCYga3k�&y"�a�T�V�V������-_��R'�e��IY�	D���a��J��]�B!�C����E��r���n�a6/0ʺo��=�����_��*�F}��� ��u�O�]���h�*��vL�1s�������v` ��W/:&�S�V��LS<����9}Q�TZ}8�P�Ng$lk2qx\A�SC�MKpɁ��17n�V�R*"�YJV.I�%UA���X6]�	r�._�Vo��ԛ5���l建� Po2�x�NJx�dW��������&ܻ��7&��4��o�q���n��9st��a<}~�r��yy?�p��1^��^] {*�L��~�-���tv��N�  ��IDAT��5>,�a �H��<<<$��>�J�~O�	��F`�t������=�KhիH'�,UF����qy˲^!p�]m8x,�o�#ɻP_�G���7����]�Bp @�N����Ðo�;\�viM��S���w�R����6�7vQ/�1?Ǐ~x��'x���I�n+��7`���X�g'�0$�k�q�G�v$(^�O~��_�����X�_P�Bz�<}��"A?��mI.���:đ�]�z	p�A�)������vz��)�L���sp9�`b��BTq!���ny2ɋ..߰eĄ("���F>ٱ���h~�k?�ܲQ�1���Q�����[�K녬ZA��2)�Y��VǤ�spO�*8�����RS10��Wf�R�x�V��v����9�Jm<y��W�̕O7%�%�G�|��SYV��zaRX�>o��t�B�K�O�|aGeܽ������~r�{�>Ĉ�M����~��*�߽#I�8>�𦪻=x���#��
,��q�����\�o/-k�}	���:�����<�QS�6��q����_�A�H��u픪w���Rl{Ɯճg\E+�4Ɋ�g7i~!I�]��� �����jᎀ>>㱙�DJI�3iٷU�X�����-�/�Z�oɴ�����+�%uf0.rN9_��s�p<x�TU~(��_��U���΄�R5���� ��,��>CG����Oi��O��Q>�Ͼ� ������\���yE�ɋWG�:��S���cY���?o�������$�L��q=A�s��T�[�o}����P?�Վ�Q��w�'bjmѱ��zw�m��E.�q1���0[����d1-�"!ߏs���t&���*�J��'��{//I�]��ɾ�a _��(Q9����=���;�Ujʦ�Z��s}_qR;�m����J�_��/���ُ?R���P-G�X���6�#	Gm���0�
�[�t�xB��>x!��ǭ+K�����0¦�+�(���&��h�nJ����}ׂG_���脙[���,}HՀU�o�\BvԂ&�!O)�Z�<)�]�g�-�5��DvY�d> ���@P����[���\HgW��`8Z�% ��z�{� ���ch�=әH	�N��64�S�E�����͹�T6�,#Θ)��R�`X�^[��ϋ�$pǘ/�_��'�w��$�����I�9�`T5pvw���l#�$Β�g�7�F�\ëW��6}�
>���=~��|nXU���?���-L`c��o�	Ȗ;����ņ����3�Dц���1��1�����Q"�]�)#֞k��j�T�L���6S�>��-����R-�q�1j�,9X��ƚJ�����[��eF��0b�&B�
r�2��u����(q�gY��<���}�59g`�7�v�k�6�,��p�~��$E���9c���:���J�����>sޝ��^?���:?��㘞��xB�ێ�;���nC����rgl�R��H4&��EJ/&?��v���z�a
��DC��k�o��~�J�e�x���10~�M[4��J�1w���� ����I'M�D�Teֱ��Q��\V���'�J���V�)�pרz����G>��hT���;-�O��
ia�k+e=q<-��Y}}��$��G���e��0+ɠ���\hI���1m�ɚ1g�:Fx�s��.`~*�KW�H�Y��ީ�0�Ob}uOG�FF$����V`;{G��H�,_�{܁���ѪE�1��	K�M�)5�:"Fk��>3�b���
�BZK��
|9:�3>�<u�49��DaI�&��:�]����d3�CX��*e�@���!j���O�8��q_.���ِ�t$u8n�P�t��j.��)�
+n-Is�a|��<:�a<��g�WdQ۸�<���QI �q����7�m�̷	�k�S"H'ɍ�`��6��\���	�~�<z��r�tR�-	������ז�O�����ڦR�\����
����Sz�TS|��	����VH�P���>93�z�8ni(4	g������*�:�h�j�*h�Y�^Ĵ �t�xa�:{R���lD&*=��䲓u����ї�EjK[�q�! }/$1��"����̔�B����u�C�8&�)K��&ųS9L���`r(+��.����0�wo^���De���	p����~O�)2(���om���JZ��~��`mu�<��QQE'���@�޲|�>����
����B&��HVQ��t��a���������+�ւ��]T��Πg�bz�y�0)k�I%�pWX
V�:���j���9�V�$-�cE�
e�eL�g�Cfo�Pg7I�J%e[.z��N�K��P���!ӤGQ?�l5�5@�R̍�i��u>��|^.�ç,�:ַw������B�縲<�ա8*�3�f�ب���+-����}�L����_�b����������o� � U����{�l��g?�r�)�}X�KI�;NB�	Z�H��ju/��Ԁ�����4���ǆ�M��j�g�6Թ_���P=��Rq����YcX�!6�]�x6�z���R/�tJ�����^��@�VU��wn^�����
S�6Ԩu�O�`47
OֵS�r�N��.=��D���Mةz��5��oz�u���$M���?��q	��_�?��=����f�>Wp���Э��)�M�s�^S^C�:�v*U<{q�kqt�&��N�0��V�̓>������:��`�,����'(�
�|C-�M%ӱI�Aߪ:�?�gd���$-�3�(�*�����Yٕ�c�jJ��1ӷ�6�ox F��	�Vυ�������FG�)��F��C�^�U�V�?i�L1�z^��L>a�R�-�R�&�]���,k�K��~��41& '�gE�j��K�����o�����g?�!>z�
����:A�|�Tf����k��3 �{�尣�/���j��.WQ;[�Ѿ�+�ȦH�6�����˕���Q�����[_HX���d>W{��U�c�d���F���F��i�7�#���fU�����Ym��u5ĐR�T��u���-�x�Z"�(�"��	8���}B�`�N��\K�I�xH�Au�7���1}���(E:��"����{�I���֪���k�X��i�M��$������+Ƚ������_����15��~cQ��֥�I�Xvh�U�2� ����f8gGlk�b]o�ta\�Z?����)6BfϺ|Ϋ�]+-�#h4�z��Z�j�?V��*L*PwMRȻ��װk���ۥ��Nَ��H���M8NY�"^��K�x���j��>��}³���{��hl	��]�����H㜝A{{�VQ��1ۭ*��O�	�d4d�\����H�����j��&���s�!yQql�kXy�R�S(��>Y5j_���};�E�F��Y
D��)D��������z������,`|xB�eI��=ݕ{��R[�-�^�R`����¾��tn��X��k����Ԙ$�T0M��v������'��pMN=Y��4�"2��ZUXgиpl�a�.��P������ ���5<��`�b���Ɉ�¾܍���Y���8CP�g���-'���'�M��A[�(z��Z�d3aܺ���O�X_����&O���"(�cp��f��I�?蟬f���J	�<���G��$�fKbr�j|z��OMdq�Ƃ>�7��ԃ4��)���{Ċwzs̪kk���BxEU%�!a�']C�tbaM)�V��T֟c��i��Ӧ�-���5-?D����3F+�ty�l��[Җ�����^<�D.M.l���8�����q��dՌ��ٌ���*Z!�<8�|��r�7" #��ax6�d$�F�+���飯 �ׯ����YW 	 ̓�u ڳm��JE����
?��X.�[�^����{�]$S)<�\v..]Ļ�TP{��
NNJ|��$x��@Z��S�98�J��p�ʤ���}��}{y~�8Ƈ�&���6ի�F�;E��ȳ�.Ag�������f"�$��Ҍ|�l�&�4pm&��!�|�!lM�=%k��u�z`�����,���3mɳm�ZE�2U1� (�x��Zؿ���v��Z�ߺ���?��K<���ݾ�~:�����M��^M�#���+e����[�:^�\ז7�����ju�dJ�z��$�#�p�
N%�<}���
N�B�����J�;�΄k��,h0����J�[*�*�_	��iLU]�c�è��.���?�c�������l��������c⳧�A}���8���o�yS=7cj�ڪ��K���Q[
JDBc�kx�6�P.X������8ǐM�������G��ɇ��D���
�FY��HQ���T�$P��<�[2�d� ��:ӳ�;���� ~��%|�����t	-{h#wUN�%����G���T�����kCm��$�%1��G���Z�cO��Q�Ɔ�}�.�A ��Q�3�}ֺ
Tfd0��tJ&)D!{/r����5*�o�J������E�D"��5�����.Z7G���W�:c}�*�DSed.}�1nH�͹���S�cI.(7�(WJ�;��9�ת|�Jj�Q�����(%�����3�3�~�:ݻ�{��tq5�о�w����'�K2( �,Bfs>�-�4�079���$&rVV6���+��"'�6��"���ڬ�Tm���3�P�3�a�%e1�]�l�� ϵ ��F��`���c�$!S}ˎPz�$��a�F��<�eL&�H��T��/aPL�ނN���zi�8��䚄��$uI�7c��Y�8;-c�����#L�N��U�J�B~(���wp�ʼ��6�ӎ����ͥ	�w�P�ٷE�� �3�d�*\����_��������{�`uuM��yv)P�}�3V����ŭLH簜��<c�k\�~�ӏ05�Cy����KR�ë���=˪�K�Ȇ��zC�g	�s*�A��W�o��0�������qE�;�~��λ���g��s���!1�va-�߻�]��p������ {p��ۮ���,�x]��b���`Θ��q�&�e&��5�k'U��#�kᯧ�dB�k�jg;����Z��S�@�\̞2D8�'�&��K�(?��ӄ��ƺ�����M\�:��r����DU/�<׸�j�W<�R���j�C��N�g�}���s�K�����1,�L�nnbw�T�Vn��	)ݓ�����6A�.AG^BFi����&s���s��h��
f�FԲ���gXK���j��6Y T:�+�aǸ�&&�4>u��f���~HU�#NLT��$����p�� n�������6��Eڌƌ��o�u���[�#ch�2/�Z4S����=�HDP.������	�pT�Xp��]:��o'�xw{���n�]#^⪆C_�KɊ0wQ_�.��
ˇ����y�\}"��k�M
�l���&���U���I<�A&Ƕc��>�3�?�z�?�>c�/���f�m�]|s�n�e��ڷ�S����Zl�Z�?6c筶�3oǝ`c�o��a��vH��<~D��8Z�ixh�jH�C��ٕ�t�7���� �|:��)�Xz:��j^�mo�(m�j��#ۛ�:�Km����K�bq�iD�T�������ʶo���sz�:��>B�T���KX���z.��قZ8%S	��嫍�'�I0���<�BEnH��-��x~��j���&����5ڵ$+����xk������u���&�PelL�rY�AS���Q�3d,= 7_��ƫmY�8����N��$Q��_������'�:��*�zD�u���wM���;}�M��5��B$��}q�����?�|z���'$���x^Scg帪�c'�@hw$hRl�WǗx�jt��/")�d�6�2��Z#��/\� �)�;߭ae���e		�-�ǔʪ��T��P ��LU22&�&�3C��a�m'�B.e�OV���9&�	��ũ|����1(�Z��6a�����vu�����z��ojgot8.?'�@�v$ar�:��aŖ�a2���x��Ȫ0E��6�Y=�z��7�Y���>�����G_|��7���eR�V�~] ��Y���.��x�{T��T���:��(]	GGs���Y\�~�W��~�2���^����5�V$I��<ZWgH��s�#m�����>��®��K��2ʩwʯ�
t|[���+���g'�*3MJ�k��ۉĀ�a�$|vՀeQ2�6�xA��e�n4�{��s	�t�]�:�v)Wm�p8�l�V�4����F_�#"�˝�"_pP:=�ӧ�4@^pQH�L���tTC���@ȹp��d�4��?3�ү��
Ƈ��+�5�x)I}�nݺ���&F�"L�Z �;���j�_l�!�[�>�pL守F~�w�m
<��V���9����s�AE�X4`%�7����|5��6��\zJ���@�4�����H�܀2mב�	�m�������s�U�}�r�۷F�g?{�����d2��)��=�@�H�r�Պƴ��(��Y�韜�:����R�a{���Y��&Z�"��`lx��)/�j�q|v���/"sV�q��朕aͳ�ﰘK��B)ys�y�5���i����8�=W;�3&�d�{\6,#�/G��Dܔ �5��]U�V#�D�i��v�9�i��ynT�$]�w�
T�2ߪ��ƕ!�Me�̽��D/5vJ���?MlPu,���K�
C����tp&`����@7���-���qm�^�Ƹ�=Ŕ��(r�4��%^�h�؀�I<QZ!�4��raw`�"��D�lR�V�VY���;h�j*��|uQ�_W/_�Dp�S� {�Ԓ�� �s�����p7�w�JGp}&���\�ƃ��8���tV�x��Y�J��A�B_�*��ZdIÐq=��{��^�8g/�GSt��S�j�:L#����5	����~C�\��T������$�}c�X0�0(څ�3m�%������)���uZ�o3N	����9:/b���ƭꏼ���z] iZ@dW�12�ě�׶R�	�ݞQ2L�\��J�ݑ��߇�T�#ё����cscU�n��r/Q�kogG�Q���Lv��Df8i�Q_�n�8�Ec��21:�[�䬷]<~�5���k:6��{*k��Ħ�j����}th��I-������ER��:p\;;����֕�:C�/j��5i���>��l2�)}�`(z ��۳	��:�e��`�ӱs�A�M�s�8	�d���*e7�����糳9\�� �uL�`b	�&Qoİ{�$V];�C�-��\Z�D&W���1�����͍)����� k��L�bp�F�QC�v.���yWg��:U��]�t�]��s��*ᝪ�*rYG�Ӹ�cÒ��Z�p*���T��qNC��E��6�J^
�pFbaD�T�%à�n�q�K����YƤ�&�{ߵݤ q>�6=7~�;��P�D9��τڱ�-!����t��!k�	C'������8l�Z�6�rp���OciaI��z�q_0���19>���ʉ�5t�a��Y!�����OozxCǄ����4�-����#��.&�'qiq�zEp��]�[IW!��uT�q�*�zO�ie�F&�p��������INr�8�ǲ��c��OV�{,�ȫ�g[�zzXޞ�{����F�"��Z�Rl��8Rٖ�2	8���BVW�_Į�'I���taO������yYRF?$I��2���G�A�J��R�RKm�YI^�Q˹�!�+%�� M.%o�UU!��8�+�1��ĮU�b6�e�3YI�\�fmG �⸎w�]�܄���J�mT��l٨���x�PM����$6NO6�\��zw�]GK.�\�W���Q̶����x��5���SW2w<S�ql׋K*��h1;n�>kAr��9\�\DT�4߾G_��ZO0��zM��F*;�N*x�qU��.�ou}���pj�ն(=���MǷmd��T`*���-�Z�S���F�T�Q�(�q��4�M�
Z�Ѕ9��L�I7�ڤ��{����6��$R�����o�$Pȏ#'����-���h�,76!�U�eP��=��M"4*��t��n��"��*�|u	3I��>*�N*>^����QE�0�U�V�W��ΩԸ\���r��qEik�u�ʂ����	���o����������IJ]�<��q,���M�:����'���9u0:oQ��HX��r��Q,^Z��΁�>i� ��`brL�$��>���(���{��	�����"
9�t����߷r�I����ܤ\R33r)��������q���~��o��_��6���~خ(/zJ	���,��TbA�|t��#��<C��`kwG�I�S�'�����)߫.A��6��;撣�T2�����b�-'�����c�v\�n1�v�� 3�ط>v���Jڠ��X�!��ř��	Ө�����I��s=Yu��cΫQ1ل�d�g�V'������z�n]���R�T:*�J���K9'�_l	��������;�p�bO���pK7���$>�&	�P�������=���'WЫ�����+�'��?��G��ĵ�����
��w@�O@���+f�X��<Gy�J1O�q�[Ũ$����0:6�o���E���un<�=�s�\�h"����m�.������`/ M0���[�X� �u�P��ʀ�m)ܶ_0��5����y�R
�B'�Z�6	�������ء��$�/B��4��y�X�E6?���!�����E�M�~�c|*��ܑ���wO���rU��x�$���&g��O'��ywߠU+IR��'ޖ���_��+����E��G7T������3v��%��Aj*'g��k��������ky�)�Q}�����y�G&�=�Q:<��"U-����,f'����c|��v|%�1cX��kr�%��j�ʒq�����m��1�_���Z?Q���9h�S�A �!�@3H$����;������e�H����Ya'Π�����FlC!�^����X*W����'�Q��˵udSaܼ:'� 7�%��#��C�m<}���tnX���Ɔ���ppx���m�3���.��\�i�(`S��T\�aI ��y�B�o��f�H�'I���4>{����1C��C:������OC��H2��|Rճ��5e�|��tC]���ưxX�-�h^O����%�-a��<+:Q�3�g=OV$M�8w�1Q�pJ�{��{@Vn�oU=S,`w���ħʺ���B�|Xʡcpg.��x�c�*僤^֘���˞�7c�X<L�b$A�6Ѹ���$Ym��pVm��J��ѧ��Qܸ:!Ϯ�d���B��x��ɱaD$Fn��F>�ŵ�i�%��������͛�L��J��C<3��ʎ$#}��`��~���Ģ�+�R�d�z���sR��7�����D�/Vq&��bA���"a4�01�3ōN�4AX�Wʻk=����g�j�����L����������ޯ���PD�5޾��Ӑ��#z~ϳɉ�! �+��B�:�)fqm�!���j55qa"��Wf�,s.8�I4�s�3�N?+U�f5l
��c2��yW,`0/�b�a1(�R~��{�3���٤ܫ�e�e����'g����V��gj�V:�b��^#�����4�	����|�s��{Bȥ�gH/��EH�=IH�nԽM��kX��Щ���?�cY��tN�휧c1cώ�9�P�)��t?؁P9�a��E��1u����l��T�	�����>L^):r������3[G�MK_���ffg��)�.�C���-)���J�m�澪71�Ԍ�� ��j��h��wQ$�q�{xrMD��sx�s���^�p�nfR_��EO/{v!]�ױ05���Ώ�p�K5�u��瘘���QF�"q��[��?G���p<#���6����.���h3�m�!y^v=�t%X�Ue���T��`�b����F"��l[��!��Q�������՛�@[:�];���pj�o;TЃ9���gǱ���	�`Nlo�1{a��-���5	�4j������q\�4)���R+��4��X�Od�& ��&{$��Wn�j��j����xv���x�O���c��<��K���I�rCi���v{}���#����'I)J1�|p	iI(�_a��N��8�.������m���%г O˳�����LN��5��T?�j����G<���]c�ӽ�꩏7�J��.���6�ꭎ�`s-��3Ɔ~g
 L�y�u�Ɵ)����V��P阺g:����:�;����S<�G�I�2ȧS���θ��*�3<Gnd-�x��E��+tg��V������silxae-��L>��Z��t�-+�s^>E鴬տ� �.�t];r�"�X����ԫb��\�qy뒼OF����W+���m?:�/NH""A��)����$+\�@�����qC���|�:�#]U�i%]I&��}[ݳi3�H!���jDԟ���/&����X��Ο����
����$h���F�W��VY���Tj�k��Az�tsy��)��|u��k7���u��ɉ��U%v6��#h�ɦ��g�_û�SXy���ۿ�G�~��ז�����׮���?���$^��Ff~J�(��{*Iɑ�x	���O��'d'��2>��

�q�b��m���;���zCl|�]\��vV71�4��ޙ�;�g�l��bS�=z�dnD�g
	ݻ,��u`+�V���"Z�`�^�X"ﵐJ�!����T>��|R	0�f�����V��NI&M���O�#�^�JRC`���5�Zg*!�#���[����.�ܝ��&ۇ���%����£9�!]O�Β|��I�yAF����~��eI�#!�|bn���WuЗdyl|�~g';r_�g?��F�����_���>����o�_������-���?����P2��HX�z�ߒ5�al$�bow����z�poд)�9f|��m�e�7����	�����{r�N�¥y�NO`yy_~�O�6Pn�YL���KgQw�%V��c"�Z���l��r�r�l�b~|^��L�TOF�D&����ud�ԏ�:f��)V�筚͎���;�zfT�2-1��j��qC6a�i'��j�-��W+F����V��jf29P��w$����*���I�ZZ�</711-wb9�]t{;�:�[�����;�u6��Yy����J��O��kbX���p����>8��븰�Vu����ø$�?��c���e�}��E�m&�<B(����3��;Rա������tQl0*���\�����	�9,I�����#�{��h��KZ�M�[��"Q#�"q������g%c���S�.�
tI,��J����>��� ���C�a�W'kL�^E�<U�w�f�	Y�9��ll��EM���2R��G;Qr	�0� ���hJ=���������F�>ˠ&�����R�d�%�����P�F����t����%�>mbw�5�$q��8�ݵ5-���6�@~�����~z��5F$����JҊ�(��Ě�.U��"8[%�bS^G	��pi1���
[����(�&�W*�V�Tŏ� ��B�i|���b	�ھ��"�_`T�$��>*KKa���9v��
ג1�>z39Ż�5&�L4#C�e�i�o��Ο[�x�~mX��jhn+��FC0���B�榇�pa���	h�u3:G�{XD����P`ՖL�xA�p�O8"A5؜`���a�'�r&� ��������M
�q����u����=�K���6��XB%3��U"���'�~<��uVW���Sl7�Kɽ"�/����A��)N1^�}�+�s�y���@8���D#l�Bu����pȮE�:z+���y� �S���6%ϫ�ŮQ��j�-tۆa�����5�0eU�Zm����d���a̚~c�ё��׼٩j����x���Q���*�	�n5��
G���T�=!�agk#n^���\o<��bK hM騬P� �|b��6U�s�
B�~S�� ��Wp��1�J�xx?�/WpV�G�Mk�r�H���]�6�*K�5����g�դv�h9*)ېC_�L� ���J�c�����#L�-�8A����&��_����>��Lu%�k4q|�k�>J��/癘�ҧ�����p��o^��?��K��Oib���#(�����&]�ظJhwpeq��QTd}�D++���/�����8O���,�ǲH�eMW�\&��&ǳ*`���yd���Ū�U�6�w8����s�)V��P\.�&�.Np��u��Q����h�C�K:'+���6
��:��x�7jt]/���T���T�פֿo�ޠ�l|�LbF�_�Q4��R�4A�����R�6A4�5f�<Ke*�z����D�l ��¨e��:P0�Ε!ܾ�����s��w@K�W�x�|C�Iy���p!��s����gkrV��d|if	�r���z�Zg�n-/�����8�211���ql�~#�e�����;k�/��\��q*�ܓ^�4.��7��C&���IL͌���ƫ�jY�H҃'�f?!`"����>�IŬ��Y^���EM�#�I�8+u�2���d���Z���~��S�ؔ��T��,��H���@ ��0�ڕ�͔�f|D�x�YS^ �����  �ؙ	`���$�vv��c�4���e��O�crdT��%v�8��n�k�q���].c����7���M������2T�M���\F�����$����Ϻ�f
�J�N���TO�%���	�I�L�4f���3
��!�����ć�����xY~����+y5��<;����7�\O���r^���_���hi�B�-�x��W��Rf�g��d�4<̎pzr�F�<׍ڹ�ͱ7O&gڨ��
 �:pև��N���PV�)��D�o;�4�%��V��sa#��p���HT�}&VZ|cN~F.��$�>X�3��)kG]�)��]}o��xo�����q���[B�V�]���mYI���	@h��D$$�N��|�n���Iy.����76wp�Q�/L���_����O�ރ�:Α����Ҫo�g:�Q�W|��}3�l�A�,b!9�8��Ƌ��u������t��_}��&�teo��P/�����yጘ��cbO�9��d�8_c��X"�oS���~�"&1St��$�MiN�[Z`$b�z.��zP�1jz�t1���W?���VOZ������TmhO��DH��SMo�8糚�p�����q����k�w��WLpDL�&���<��!��o�ƙ�?����(g��oΡ8>,8gK��Z�̺.]\ܽ�D���8����.��/��19�a����q�*D�& �s=Z(�vQ��%V1*�pqn\�|��nac�X���)H�꼸aT�1�6;]-pSlKiҡ��Sv�e��/�ի6�4
�L�Hy$�󵉘=�=3�F�#�;R�X�1��>ʖ!��>�L�I���{V�����I��B݋J���8��P����	�eo6OO�޻����:�VK�^����175�>�ӣCH�ꂡ�IGԯ7�J
�hb}}_���\��i����c8<>����*�9��)����q!+�O#uƽDb�l����{�|��I,&�q�b��-l����'w�������g��d1FF\��Ex0��BV���y���`jb_�:j>פ�I����3H�D C4t阊�kqI_}�|#��"��v°�<z�I���-,ٵg{0v�6@T��䬄v�,1_��H\��C�����.�O�8?��%���&}�79,.�H���G��]e�s�,R ��r��q�[�|e�sy��Vq������9G�s&Ì���9�B��.��8+h̒016,N��_H�~j��&$1��9>��Q�;�rN$(�K�R�E]�z�S�V�J�d�hSt�j�9Sƶ��1�M9�<L�ۜ�������L�M��X��d�[���(��ä��m	��:��AT���J���k.�HB��'Ū��7(�����|��F2茣�J���<}���Sx�\��V���A����{<���/���.M���>ַw$�cnzƐ�z�D��\�S�˒��Cx��QԿ{�c}̴#���6�p�C�(qO��5sd��%}{Yj��7�r;B��0(�J�?���{�Ph:�T�8sYi���,z{����	�QoU5��ᶌd+��G�S4N@cP�5�i�
���ej�$��z��JHd�-��Og�0�bd!�������&���1�_�bx4�A�E*V�	���]���)V_I�	)��Vn)`|������d�:f�'���%Y=�g�.�=�?~}��(,_ƙ쇕Ǐ�
_H'%8���x�n�c�9�'++Z��y�1٘F*בgsI���u%Uֽ�_G&����	�O�ً����IY�2������Wf��ְ����l@ި$(T�e'�`��nMr��dh��1��D\��v�B�����)H�DM(����<����N6yKm�S�PT)*0@Wt��gh�3H�����|^��G�8���eE�B�N7�~M��e�HBQ,Ue�S�<�Pr��E�{m��#4_���|]���a~4�/>��_��+��$Ǜ���x�!�'ٸ���ww���B����t���z�-�HI�%��5*I	;�[�H�Ø^�����Q��l襺������܄�Y��J�h���ٱd@�\F���A�R8�]���\\��Qev�≸����W�J�J���O���~�b�	{��)V&�w�i�2���"�aV�(^�zI��9Ȏĥ���<iMܗg2�?��������h\^W�Po��i�=5��I�z��%��w�>��]鞜�5�3\�<�;O�XY�B,����	�ܽ��?��<w�Pl�)�E�+ $�/�pR�mFD	����İQ�*����"�#�3lK""����X�0��,Mc,�9�{��W[���82F�"J��ƛ��?�ʣi�,ɚ x�y���Q��rQ	�����K�L5?5+��c
��9��I��*�&>�&Z��?�X�{4�5��>\=C���i�K�)Ԫ״�O���Hn�T����C
SE�=���/�ǃ��x�|�p��$�-���?[��%iv]����gf�w��LW{t�	�á��%.iIҋ����$���<̐��̀�� �MUu���>3"�{����"�	X	TugFF|��s�>g������b��f?̤���u|�`��?�����l�A�����s�&j��_}���9��{��4����2����[�T���":/�A�ULd��lQ����1tx �y����7cƣ�>���<>����<��/^�L����==�w��p���NH�l�<:5۩9�r���;�+�B!�g��T5u.T�_F���@= >�Ng�=&��{����h���ͦٞ�
���=������k!d���8l�>cT���4��g��9����ś����\�uag�ѐ�]�V^U�J=z�z��E�S��x��-,/��Mr�vZF�7�8��X�S��3���J��|�\���
	�@���܏ߍ�ĕ��=����e��Ǐ�
l�*��y�b�k��:;3�s���T����#$!�Æ�0J��o�gC�� �D	�m\\6���a�Q���M��	��B�f�݂��Uщ���<�_�{Ev�g������4���y��Y�,07�}����khf� L��V6V��Y}�K ۱�������N�/�<w�����IsE��DARI4��n����ϯ�ա�So����XG��9G@X�s���RQq���DgE#Wb����O��`b��!��T��%�aއ��i
	~�1v�OP��cv���R����eeE3�:}A7'+݇'U�"�3!c��k������n�6pMT
z��f&�J�;��?�k�贈_�㬜�t�^�#Ӆ�x{As�]jw���˕�i����8ס^�X�F��|�ug�_`�Q�����
VWfq�}�k7� �.�8�9C�%fT�ޣ\��k1?޼ٷyY��$�#�j�@=W��`����z�ʿ�w$?L��D��0�F:��L>���+�TP��U�-�c��]�J�@��Q{�v�
�A�˫�(�V��4��-�)W��{g.�JT @�֬s|A�K�f<��<����A�_KLO�73(J�����(~/��_��������AU�tؒ�F�g&����vY��$j�s�|��2R�LPV�S�sq����8>�|WM&�*���������5���P9,��`��`�vJ8-��ed�iT���8?�/fsC����sY<z��<�Y��/v	Rn��A?K�>�)Uy�ZF����=5O=,>�6�E�;4yv�,0I6�AU�n.h�	8��]�r}�/<p9=lp��'�㪜����J~�T���{'�w�j3pZ�P��2d"��!����1sq]��Ӈ9a��"� fI|S6�
�dr~�.K�}�5����������D��m0������~5	��g��Ŵ<�������?����NuU���\��/�6c�4��B.�D��&U�V��?�Dq>�^�����U�u#d�����NG�L�͜V�y�F�@ła�u������21�%i(�	Y7QjzC�[�,�:�6+��h4�NZ���:޷'�.�[g�!��W՜�#};EsluI��Kf�r��4��W/v����$�N�U2��V��Et���o��s\Ϲ����'�����ON��W�7���X��A���:F�s	�)���S�z����pRo�{L0������*ˣi�D4H���0��r�������\,��-V�ե}|���& (��2OOـu ����f�gx�v=Ϡ�t��B��|H{s擩�DU�1�ݞ]C��$Ьv}St3)˪S?�x�x���wyMgU�p��$�z(�z�Π���:�����S���������nu��ͦ=C�?��L��1�n�A �B��$�MJQ�߼����2>�侉˔Ύ1�$�|��vQ�\�U��<O]&��sW-L�����z�������E�H�t��^2��cbFvk�L(�G��1/�>���\j���I�:ܻG ���F�	��XZ?�S���ӺQ�t�JioJ񲂊��{3`�� �c�����	��r&���TmnY��Jɩ[���W+q+���x �*j"[b���e�������W����U���psϚ���Б���U�؉��8�Hy�{-�w����[�����=ę���Qu�͚C�`�gܯs�T�{������u<��ų��5�ݝ�m<}}�3q�������CQ�ΚH�I��O>� [wo�𲆯_����r]�13r�ߔ���e<"`�j6l�>tDu��x��|^occy��K�a|��
�
�x���{����K��ј�e�� �(IH�W��0��@^[��.��;g�V{bs�S�i����U�	��w����o����Fxsa��)�)�+��2���_�W`*�����lc��
���C?�&A'�d>0�H�b:�ؗ���	�$��=����[R�J'��z�1y�\��j{�Wx���TG�]���%��GN/.����y���*h��!hSP�ã3��bFY�4�u7�-�W&�1:�}Ya�s�_�qq~�f����,s�4�	$��r��=S��g�ٸB�F;ԥ�ؠ�߳��=bk����ا�T�Rk��Xȳ��tzv>,9�xL%�����pZd�����3Ӆ�	��Л�{9�;5�w	+�.��}��n��~W��k�y »<I�8ufh���h�����Z��_���b�k{kc	)�L��<s�=]����	���+Al!+6ɋ��.����C��K���\��a�]od��a~���8��k�3R�A��k�\={�U�Ս�܇	�X�c�y��'�\��7׬=�"[��ϵYy�9u=ʬ�1�4�vV��	lӮ�l��+����$����8�7�>�.훮�����)W�ま����Y��.������MLF
��'�,�t�o�wy���:e�<kp�S`/-�Q)7�{��"6֋��;�$�z�g�y�4.K��Q����S��w�&D �k�ah���]]��9r�2&�L�����FO�h"�iuy�fy��&c�&ʨ���;%�|�:�!�N���,�V���V��*`��[k�q�P(�ΒnJ;��`8��C;���_>go2-dۼ��E�*�8�p��ւ�a�(O��)/=�0]��@�6uo���W�H��Lf��Z�������\�x*���)��K�X�O���'�/������7�������}����e�柎Mf��[��|�}�+KK�A��{��0�3kjq��R0Tp��s��ac��gi���1 �`qc��"���ban�`��;��W�<噒�D�)J�G>���/�'D��;�$~ȍX�2Y릑��x�F!Ь�QQ���^y�1�D�]��9R&�l�-�)�xT�)��}� ���/ڕ����pb@ydC������M���Ƌ����S��F`C�,?�a{TG]�z\V}��?�7olp�X_�1��^+#�IM��߽�~v��?�+���C�g	�^��+ͤX�e���2�����P� ��'�$=�~�WϺ�q�6�V�����-`ie�,D��.1�R+��(���́'wTeż��N�JωϦ�}�w|�Օ�H���%�A��5	�*����D�X�*X�9�C�T#�ә\N��&^b��95Oӌ��*:�N��o�I	{��k;�U� ��psc���^�uYJ�0*%�0f݊ ר��%���?��#��!R|���~��XXN�`� 0g"��?�O��S����*��C�ɢ|��<�����9��K�SY��I���TӔ�v��P�2Ǚ+d��� u����<��������'?���	��E��������M�,��x��
LLRZ�QM��R;�M�!�U�L�'%j�u��u-�1��:
��K��±���<�ޝ[��;��Vd
دsG�V�1,Z�ԊB�|��&p��3d4��e����Bب�~�q��j����&�1A���͵"�K����_|ŋbb3ۢ�?}q�da�%��=���lǧ�J-T���I̯�cJ�g�\�����S|T�0���_z��@H�
X�Ǳ<?�XJ���-���Ɠ��E������8�C����z��Ha�\ߒ����p�GR�U�Ҩ�y��o���OאId���������v�)���3Y�(sG�E�p4f���:��:gF�	:!]��iL;�yQv��&PS*�Q�T��;���U���8@��׭0�H�9��Ƴ���1~�M3��"ܗ#>����SJM%y�t�b�bqnw�����,����%~y�ff���F��!7������@�h�G��Ǧ*�dB��U�O�_�7߾F�
@��8���hc#g�n����a���u|�Տ���+�}�����Ox�͙����ϯ N�����JE_��3e�lá�r��ƣ�i�ƒY���o���[�F����nR����^�n/(.���3h!��S#f��R�ԗ�{���?���Ta�ͣ�F�hdI��(�Q����*�0{	B:��|s �6�F��F��8�u�J�DknX�� b�����7ħ�@6�1[�7o��g��������"��	�h�h\����E��܏�)R��od^���)��0UqE���n)�����S1^�9�q~a��"b� �Y�X���&��K]^`�9ڌ@�	��O��Ty�R����w"8��c{�w|v�
pRvn���̦�lA�^>�J�� ʦ~Mۣ]{��)�i�l1v<MNߕ�]��{o텁�&YW��𼏕��#��s��fW�5\�1�/MQ�u����J'Ӹ�����R��l2��n��ʂ	l}�b��ڗW����A媌ӓ:V4������#��z��>���Ϭvc��s�G����gN#������F��L3��y�~��q߼�O�u�2����1Q|��u�D��#�S��6�L��aĉ;�M'.3	�L��R�z�� k��:��?���|����Pp�<e�y9�5�#}O�:¼)��A�)*kݜ���b��0���?C��3����E��wT9�'�o�޹�i����	��Y`��p|t�T:�u������E�Vs�kx�jU���[a�丌�s�?GS�H?��N��D"��J����spx��f�g;���5������g'5��Z�&�d�x���yZ'f�N��E�R�5[7�f����IWs�M{�b�F.��,��Ku�b��-�X���F��MG�p��D�)�b������D���T�P�ʃq||�SB�?�j��b���Y�*�$�F��Nm���V1��W�Bh������˄ݾ͡h��	/чw17�)��`=G���q��C�irǾ��S�5q�K���/�	R�&�����9ic㾟�!�O�/cm&��T?�>��U=��G�F7�$P�ұ3Ŵ�mq�g3K��^`� �;k96'�<�C8=6���u��T��}��|ь��-��ĔN�n\�����V[~�;�u�bfLS%?���y�:+�a��8��>^En7΍z&�n������2��f���_]0�����>��3��t���'L�bX�XǓg�����YgN���{Lgy�-Y ��G�de�����=1��J4��ؙ���}}G���v�g%)^��j�|]%����$򳹨Q�f
I�|s���y6�2������ �EL`d�TE�vG<��v#X[��V����;�yW��]�tt�����j��5���x�Li�����Q]�M���T�-����u���y]A7K(P���,�݇�1	������gQ{ٷL\E)�`*���}R9�|��x�s��v/Κ*�+�D2�l6o�w��>>�����@���&���8>���!�Y�r�6A��Sִ�5�x�{Aj�-&�~���B��}<ke&��^=C����{�X[K�tK�s����Q��R��8i A�&�#��J`ls/}T�a�,U<��܏�M��?h�gFf"����F+j"S��g�<v�g&�0q8�w}�������	�VP%oj;0��O;M�A��y�]�;�ӀJʡ�W� ���A����)���j8���@k���bKs�����'|��K�����(�
&%WX\\�󯿰�����1F�8ffR�\��oͳQF�d�ay}����?��19B�/���%e�W���YVņ:�m��bO����/���������.:#tx��:i��Ql�g	x�(>9�ώQk��|�/>�'��^�IW�5S�3��o�o�l���G�H烨0�T��v�}�<�{�<tĒ��8����, �߰�Z�Nɝ(?�0���ǥ���������(鯍��Y+*�BaH��Kgg��^E�J��	�P��n����X �ը���U����hW�����[��N���b}s_��#S�7��� ��ac������o�-&}��a���c�����ܽS��?B��wsYX�P�4༸���YEmUR�L2#��#��w�ȧK��2�G�P��/ױ�9�_����r����Hr�X��$���g����,��)���"Ļ��f��v�bg����������^�/��,�9��kd��g�75N�h&�|G%�
2���H��ëF"o�mh$f��3��H&�u���  ��W�����c��I�c4K�i�u�(�����b|��U��3s��U��W!cO^����)�?=��Z�Y�_�@�t�x61Z����6n0�Z����ĭv6T����Rv�\1�mw���ݾ��u��W8<9A��n~y�	)�s2�[[ܷ�|��%�Ԫ�d'�Ub13�v�W*�Ea$8=:� �=ƃ�;>�*���b�U�=���'��dX��ĸ��3��|N�����^,�J���]���@�	IL��n�l���QPU(mp�oI*� �*�	l׌:�n���m�0,��τ��2��x��������-����G���OO���"�f�^�����.s��}�no�ť�2�.M��oc	>g��?�Es��������QgG۷f��F�(��^�a��E��U����]!���yVmٜ��,S���	 �R[�BW	��̿N��:��L̄�\��s�!�&�h������=�U���gz�M�^1�:7_��H�S�7P/����U�X��C+��y��xWƳ�K)y��l�Q"Vױ�;da���C�դ� ��рd8�.�HW i#?W�Nn&�2��n�)]��T�ϘP�X/��C1V�nR�?�|�������F��g��kf���u���,�xC��xE
����̩4�#։���V��J������L�U3��A�ｆB.�$�F"4q=�h�ͺ14�^:���Y��,�=[��6p�~�qLC���iZ��3�L������k:r(S�n�h��WW����9&�L�D�	����US'6g&�����?��%>�`oݳjڷO�8�G4���%N/ZX(.��x�	�,�D1�����6�G�%~������rfV���o�k	d�j /��4t�b��x ��4.P���]�/��"��G��]�����&e��.z�丯	�׿���ka�K���v�si&��t
���d:ox��{����	X[У�xݤ����>x�5L<����B�;�n�E�5F�R���{3y�hx���ɸ�����c��z
QLڇ�2�'^��D$C�AN�Q��ah�f�@�Y������)7x͸�1��9n�`2�fO�ah�sqe���3�9|yh������l-�Љd��%A��0`sNJZb|��%&�~<�a��n��8_��l}�n3��;�^vqY���Pk_3J�r�YDU��3�S��1��erv�ow�z�J��u���j��E�y��wH&4�eRK���7U=G�p�5v�;>���3W�ֻ(]��E�z&�7��G��
	>ov�<��L�v�^K��HD	+o
I��ay�%D=�{u���V�W��Ɛ�fq��-&m�j&��D�e{y	��o�{����:�u�g�e
�M�_t-�O���ӕ<;/\u��\�r|fR�t~<aDqsy��7�s_7�,��/b��<6W�3��x�W��oJ8�l�5�b̠i]BU~}.�WWV��>w$��3i0Ж��啙�'c1;;K���F�щL�^�d�G�0ys���9M3��;J�{��5��{7�dzV�`���:O>�\DX��6�u�enx����ͳF�1+,uzut���K&��BΙ��TxɟU��K6�sxd�'�_4�����eU�4m~�������?j�J��9T��,z�(�71U�L�A��~חQu]�Q�����>���ظ5���>�è>���am��>���$�q?��`��8�]�)�L��wNQ{��if�#�|Nͮ�=��oxAǙ�/��XKgl��Y�en�a�W)ߩ�9MFv�$�j�L�Co�>JL�ػ}䇳<�G�s�N�M�����EG!�ppb��D��4^�ŭ� �W��Y�?p��YI`$��뷘�,u����%�'��q������}�>b��{���U>d���;k'�w���O�?S�@L��C&������h�Y��,����!}ߚ�=���������"	�w�/xDPe��d�g9rK�_��/���e|��>�jW ve��#��3��联eO�������M��X��Vl�V���S
��������{���+Tx#�o0��NA�=c�H@���'���P~uP5Cu�ń�̦��0.�|��g��T��DpX(��*H��*��9aWG�i��$^<=��o�E��9��X��>>��J�e�����[���{����˗r�1Y��M�e�8K����s�z)���>'�ǰ�ƻf�s�l�FP-v�螙d7��8����o���U	W�5󢔢w��dm)�t~ك�����C��i�Uqj� ��h�G��T5�~]��l
E��B�p�X7z`109q�����+n8EI׹����ŋ��":�q�w]�w��9_�c>�˯��.���
��>�\\�GД��y��8�d̍F�>�:<�>`���[�9q4#h�1 460�"��L�V���ZX	ȧz	E>�Lښ���^]u�19�zv~Ax�LT&8���!pmwF���r�V�gX�bq��'U�GƦzohsǑ^��8�x���e�sQ�,v,ޙ"�7�(q@��M�X����HǒF�WgE#:*��Cq;w�+v�9G��OsX������w����]�:=�ӎ�Ёz��N�ry���G004�!F��#�d�x��lЌ��[ڭ4����)i�饹Y����֩�$b^�������
3��x�F���.���	��s��Y>�\����G�.�T��Q�`jokF\Ϧ+q�f�ry����2��[��TA���h�T�wa�wb�
{��~c
4x�M>7Υ���u'^�`b_jf�dO/���\]H��M�BϭZ�{d�pb�?�S�G �ٻ�����Cl,�a�\�K�`��2��������M'�j�3Q� �hM6n�!V"���>��X���%"�n.���;#Sm��%����Z@"�����Х������O/pz^5��įM����5�KU��_���#f��X�,�8�����E<��ͭ9�o��I�����W�88>����aS{�x^s�=CT�<U�z=&�ţ2nߚE�	ɰ�a�H]Z��DtH/�y���O��Q�|����0z�>�H�gp���@����vO��%�S;	���eB?�XGP�u)�jfO��ZsD��$�� /~_�.��4�{��i���]��|���D�K΀vo��W_�cr4��O_bf����������l�k0�����O?���V=6n�?"�P��̮�Hz�XF��W}�e�F5ں}ŵy|�tO_�a��c�?�E=���<\g`����2^�>�i�ʀ?���Z����=v��2m�A�,o�d�62K�L�.�Aedԛ ��B*�V����]&@Y��TӒ����.`8���n��>�@3ZK��Ѡ�^��x���ܪM\�q��b'Mm~��72?p��Y��@W\z���(����
|�I�p���9|�p~&���L�cV�k$�0[��&��;���<n�[������sm+�������������ʀ�ҬW��K�,(����&m�>�Zm>�	�6^2����y�~�$�_����k�1i�I��ʢ�X0�D�g��>�B]��`ں�P����o|A�������w߽��� ��3���"�l�*�&�gJmE+���&#��m�@l'���-|�!P�%�z���j#o��w}�	�Ԍ�(�{<�{��a�-��0C@��h/�|�؎W�*.��r���X$	l��_m#�����=5�P*׭��gq^��(��y��������p��u��h�@�N׏�UO��1C�pz�	��S�)4����ִN� ����x����!���*�K�kP��.�gϷq���[�s�E,�����<66���k�	�Y�{d�~� Y��J�hť5���_}��>�<k�����(��OD*i��D����أ�t�܆SI�	��fs��:���`��m���\j>��Mz��>�Zt�T���e�	��5����PȃۘM��g.�L �Q)���{o�P>9�nd<Y���;<���2��x�n�����*����g��s|f�x���ͷ�3��1���������"�ϾivHA�M#?�j���R񔀅��l��_Z�Dy&��h_Uq�z�-b)��L:˽B��D������[("ʊ7����9t�1<yy�*�j�5���tm�;I�}�,�ss�TJ�FE.�ٴ�}+4(n����|��ٳ�=�uc�5�;j�3���W���F�5h���Ί�U�}F��6�$߾�j�
x!�;�W�F�5b��c�`Yj{[�KVL�r���:׼^)�2B�4�{W�V�M��dy��R1���&f��9��2�,/�3�����o��nJ��] Gǧ�O�)�;���P�^ >ǐZaC9��,�4W|v����d�)D�\��3O)sS�3�n��+��%p��1SH��C��6 �h��q��O�ݳ��4AP�^���������[pf�.ɔ5����=ewU��X���󅞎F�>���Z��}����1�z�H4~[g)������)+򆱲���b:�g���J�14��g�Wo�pĄ�@#���nbw��w�&旖�yk�犷y[j�c�J]�\��G��wpt¸-;�4������ba�� W*�\aj�7;	Ju����`^jV(�x~$���D2C�V���)n�b.�{�����L�m涵.�M��bƬk��Q��1�O��˼k{nFPtKQD5��̪�v���p|z���#�L�R����b��În:�@�o
�_�����B�>p���=���?8�Vލa����/]�nhvL˙k�x�	�L�W6"c0���f���� ��W/_�{z�=�yZ[[Ǎ۫�;�x��-�Ƙ�#�j�����Ӳ�T����N.<1����N�n����6�;B�dmƖ�0��׶1�|!����	O�/��;�f���6��?��$�.��{T�8ok�s�M�q�Y@93s��Vk��v�y}��%��a��8R8���LX����ќ�8ܽg��5)��x�������7h�][�Ia��qK�ԽI&��81&�M�::�(��[ԣH�&FQS�DsC=^|�sy< 芌[����1��d�d����gr���O_~�� bϞ����!��>_�oՓ[w���[f���	��G&3�6�	X0!�Ag��ŀH�g� n=���A��_b��J,uf������B>����9��͸W��ԯ�� �]���YnW�ͫ#�9��I$�~o`z`Ju�z�l��)A���sc�^�s��sծ������$���� b�12���ޅ7�
͸�j �80����4�ڱj���&M}zv���/��옉���F�2a"��r�ä�7	��0x����m�@�y�/�B���5\]���7����~�=�4O��_����A�{>���Ѕ}���'��kX]\~%�*=ԙ<�k~.n��A������˝�<�;�~J"]i�P1e����E�>^�=�z�L�L$�Ɲ�����J��; ˒0�u)��&ݱ�&�� ��4�Ъ�y�l.������ߋ�����^�G�N��m�@�Ur�L�L��`K�g�?r�S�ȇ�oT	Y�Ho����Nͨ�5��pk�^1��<O�Zb�ń0�ש6�Lj�*�Kj2�r��X]� �.����1޼��L�3L,�/��/�受���gw�u��j]>�L�M�Dɿ�7* ˤ�z�J���_L�obE�'t	ɚc �'>�ӫ3\�n��&�Sl�K�[|��n>X�7�_��A���{��E������"�簘I���)�{~�=��T"&�E7?��+���8gT���=��{�T�./�0.�7dc�=����TJs^Ҏ��&�+��45��=2r�Gu$u�te-���Lͫ��V��5l��T�W�7t �����Yu��n�{�H��)�M�2~�._s�$i&ģ�e�r�w��7�\6,)�T����kL����]�勊U�����W:�(sE۟G�3���Ư��x��D]�g~�s�X^��Ϯ�5{KXBd�.?K��1f��=&C-&�!+�+F������Ed$�����E�[�n���)$�1�Ĥ�
�M�0qnb%�����֌>4v�K1Tj��[�q����p���p��g����h�݅V�E���P�3(��x���n9&���9���3�̅F�����J�UѮd#�������n��}-O;�%dI�Q������ѧ��~R� �b29�xm��,�qk�&��:��_�'\\���=��ܧ�G!��0�GdS��JK�d�"�d�&Q�Z����_E�E��2[��/�ۇ=����E���fʴ�T��y�^�e�c,������6�.��(���T��|��X����n,�۫�S�}���N���^���|�(���"f���3�NϊD��1�����P^�9Ĳ9>�G*����J0N��A�(�0�q�5Y�t"l���ϒiѹXڍ6bkAƇ��Y0�)�F����1d#\	1n0��h�g����x��M�r=cX�(-Λ�F�gj�fo��?\��G?Z#�YƷ�m3���?隶���%^$��n�L���e�;��%����G'��"7�c�TG��ua&+3E�EM�r�UĻ�ʅ,���	��Ĭ$.�����1���	��AS`?�y˼f��6n*��T����1��_�9�.�`~�{k�gw����Q�F	�+͐a�~�Qɸwҹ:�^�_�12�N���J����`�Ԛ�����^�����QKpGF��Jr��y���ռ��DaL���A�R��z������֊r��n�:�4�����5�_4¼�^�Y��K��êY�e�<z��ٳ<��i*�����zλ߇����*����~#�4�׊R%���o_!����C�E6���ű���g�<�T�;��0W�E�i��
��Y�(5yf�(��-��T+��5��i�O>4�.��ll7�:+f�s��%8�Q*���Rq 3q)ny?*o��n2�]QWzܘ�'�ʫ������"�&G؞�X���W���hdL���Ol>Y�����;pg_���sj�z˻�XV"7� ����m�3℅B
�����܌��u�c��Ku�uO�30/��nXB>��m�Z&�*�8����MA����踆l����1Ê��vd��2���\5��)k�hnT:>?����H-�oL-Y���EHq6���,.�*�T�`��?K�cI�%s��}&.��{i4����B	��0����R�KwW�.��9�i�'~�!��ǩ���5"����'�MY�f�\	q�,,�Y�f��;���
H!��[U{`ʡ�e�:4j&�g�O�%úT5���J�&�|�ԑ3��>�3lޞë�~����!�q�q|x�Gxp�6���Q�\i�Y�TI�U��Qwl�_���7N�)j���ڛN~�t�7��x��hL2V-h��v޽����|��.��\��;����f��R@�7y.s���UTC�Z��؉�+��4��	OG ��G��e�X�%#$�Z@�A�w`M��	_ͨ~J�'�k���'�{=;3��P�p]
�O����2�$	7�&�x�S04�90��:Q�,�EN�TE[PH�bxtw��Tf�=�~cq;V���y�T��OL�#X]���4�T#g��;m������S<c��wc	��_�t�T.땡��[��Q�T�|>����g��{��uas��������Q��9���~u�j��ȋ�{����,�"��5��<�>ǯ��CW�������5B�Hϥg�(�ǒ�g��lv\�y�y
����_X��������uy$H�q�w8�(�V�@�T���L7�Q�ǖ8�s(����5vJ�>�����C,%+��XT��fS�},�Ǚԧy��qr5B��ar�Lj�:�m&�r�v�kHg��UL^��'y��pu�M���5NK8>i�۷���m�͒�Y$�=(��ê���A����憬#��x�A�����w�dS��8=m#�x�k�߻��W��)�TQ>|C �!�n���J��L�����>��0/ِ���j7�)�(yPe-7;�Ӌ3�������]�.u�� /�a@��g4:�d��ǠcD1����&��g���I�k�>���o���=̋Ѭn���3�����'�/.��|ss��
Ͼ�5~�c���Ţh�L�J��?��?ƭ{+�IP�x�j���2������d[��X,���"ɋ���Į:D���{zh��J��m��W๸m�y��D"��C���h�%��<c��-�z,�B��½����R�������+��e?�03;���7qsu���LX.�~����˝2��$|qG]W�h�Z�'�� $�FqƯf�b�T�7����y~�g/�yA�\��)���yM����Θ��<���L^^�o��N��=�a���l`��s^tcS���E�k3���A�>����.]�3?W��0����X�{y������Z��Vρ{��/��_|����%�^��?����s�8Cݾ�5����2r\���~�G�{^�:?D�IAs�{��T&���c~9a]��{�k�i�ז��mVV�Ţ��SO�&�m�1�l�g��������|��*���p��-�,嘔�nF�����7o/���[<[n����N�mF�C3-roTpu�T��ݒ��?��=���1��� `�$�B*y�*VN$P��A�e�ȟV�q˲�~%r���y����F�{5b��Y3�tM��o @�H���
�>�A���Y��n��C��`]�z����@c�lrO���UǣÏ�����̠��aB��ոPX$ �5�P�5˛Ãc�yn3�Q�w�o����HGMhgrX6�����#Q+F6KiS�ވI�Ϥ^gY���^�nb_�k�̩<F��E�t��#_{f6M@5��Y�����f�s�T�k�L�06��|n<�$2K��輄��Q�a*���6�f�=)�+GS7E�Q���ϸ��<�{cɈ�D��8%f�b�u����=��v��S:�S�T�P������uӍ�|���q~z��Ɔ����حb}}?��ޛ3x�sa�*��vg`��D�u�b�SS�N���8ԉ �����zf.��ՔY��S!T�#k�Xl��v[]{�Ac&�О�5��� P2#u�.ߧ{b�Xg�@��ڌ)|�UPf/W�>�1���U�N�M�!��S��g{<3��ݞ�\ş�ԑ�����\����x(��%F��QO�&R�g���A��d�n���[�'��ko80�:k��8�]��h�6�	鍭3�n�0O�s�9�rQ����s<7q?�E��q|Z�s����s��{�[�Eܹ{��f�i`�5��32�׻�s�k���6V�0��۳�yq�����f�c��u����	K	��q�n�T������^�`��{&��/��DBd~\u�'>�cc+�E�h*��1�9��4��h�^��Ｖ�2�/_����Ā,ױ��`*�.������HPs�j0L��\MdxN`Q,2���ufC����=�Aw�����` O��W�r����,\>3c�9��2,����U��M��U�a����31EL�g~i�{�C�����d��& �B�8��y���n�����]^R��Jl$�A���r�dč��@#S�rj`���0���(�Ǉ���
�c�h8��Un��*g�-����٬�ig9<�ᒠ��M5�e�� ��Ǔnv��L��@��g��{�YTe<�d��~�
�Gi���pJi�lni��y]�\���=�F�7����ל����x^�Lof����|U�Ϳ�I�um!���׊ Y�f�����9}/ޞ�b�:h�R/����<~�'_�B�.U�$]�l�qY*Y5H�6�򎌎��-p*���a\�	D�yT���+�N {��U��z��S��ګ�T��lN�8��5�o_��a���lG�3����Q�%ntQ��
^�A��X/���2jWm��h�F3v���ϭ'���;��
/��϶�l�T�Hz+�Ț�J�yIym�k��IT�)���j�EeNS��'k�s�	��h�����G6�;��J��qY#+( ��5���lm�ban�39��3�����;/y�f��W���.�W�Ll�<���\��{�x�$}q#��؜�Y�\�u����3�}��kTO󘉫������Z���f�8���U��)�9��S��k	��_���1����K��|ޞKci&��W%&U=��)!\�g����P�=��� ^�
Z�@"t���U*{�-&��`��*?��9uq���vc��h\�"� ��,�,��[Q���h��\{��j��?�Q2��w�oʁ�錰
W)%�
Ƽ�5Ͷw~�'�3�J�31R���׻sU������B�ϳW-��RˏnEI�~�W�������#�s�{LD:|��7fqcy+Y,/�p3�j�����߽��ŀߛB~vU^l�u�f���3�w� �g���3/
���<��wV�����ᰂ73���RO� @���m��i�I�	*-�VL�<7gT��.���o�JtZ�s[�&�s���]	l�}���g�6�~���>��y,�ĭ�(��l
Y�ddϸ0�%,�C%#��z-�p����Q�C!���dU�FER��C׊�#�l6��������"�a ��ٷ���������$WN��{Pʚ�7� ̡�9�gk!ƻ����-,d�3�X�e��C �Dw�p$�����R�;�I<%5���~���21o�Ȉ:�f�d'4�`*0�.�*őd�f����J3Vv޾����G
76L�gqu��̘괺8���������IM/���e��ps���0q��V"r��*��˻��߯T�K���W��[77l6hV`������o���}W(3�i��� aGkZ��W�۽�������ȓr�(
D����)|o1Ɛ8�KL���]��e�b���/La�J����f�X��3<��c���S<��׀��E�^[����O�1���>����9��jsl�=�d�\�3�{dq6��b޼�Ԛ��)n�jZ	.R�, z&���\w�D��q��Dj8�!S�����kX
-�ܙ��6V��q��t�F8��!�x׿>(�{g���T0��*��fߌĳ$[�
��R���Y���'`��V�"ν��Em����-R#�V��q���y��A+p;Cz'��g���T7?��p�7c���'o��$�#A�B*oU�g^q<Sc�`,g�z1�4�	�W5���$���ML�H��f]l�z��W��f�9��4������ͦ����e̚��s�3�y7�Q������ol�^�P���d���}?c�%s$5�3�_�������T�><�Yq�𼊚D�C)[?��I'���[]�f�b��R����\f�^���.PA�J����.c)���Dǲ9�[b|~��X�XRL�*_
�N�W��K+���7S1E'���2ՉQ��#��qO	�L���|�{����Û�1�C�QB���=6��<6i���8�iΚ(����k�qq�<�U��i�F��U<��[3E3��tּN������0'Ts$�J�ڤ��e���X��낪(»˨��'F�m���Qb��쌌�H��!xS�'��S��;q~���\b"�x��{��n��������R�3��SQ�i���� �l��	jP���ĩJ�8m^��5V���x�0#c]�l�5��}�Z-L%=�*��(����Z��)X�K�X<b�z�厉4zCl�b�	:���������Iܸqϒ�A��Snvq���m.FA�ѩ�7����G�IN�9j�̪�<^;�]�c�~�)�ݬ�	rx��wh5&V)K%(s��c,��"�� V�б��X�Xjc��QN�sL���2�Y�C�~��GƟ{�9Q�$�����ŹU�ꭞ)��DK�h�bd�EjU&��{�7O���'C���TǓw��km��Z�i�����u�ȆS#_��Gk���ŏ?������]kM_�r���:��,�؝�������q%���k��gX]��6�>���<r����0���R򪓷�D�<��3s�QX�\5a_@"0�Bu.&v�֪r�$S��U����
�/��+���E��xȊssL@v���ڏ'5�	zH���<�FK0J�S˕B��K晉i:����j�mJp����m^*r��:SO�%��H�V4������z�!��̘uw=o#gA�h��f}Lz&�w�X���M�WT��n�.�BLjTi=;�����-me���-&)���>6�q�@CE�g�����7�/f-���S*�7���e�^�-�Q����;/���Hp�R����0��\N��ʼ�D��a��Ⱥ����j+����f�pGLj=posU��wC�Z����^zK(0��^8-��r��_��� >��ŀ�+ʰ��y�R`S��o׍^�TB���T��$��.~��hĄ�&a7��f"���v��)�I�����y�B�K>"��'�g9�7S6���&�[]*`�������i�f�fJn��?�#ln.uEf�����!��sg�|�zF��@�%n.������ je`o���7g8��+��y����"�W���>����Ƽ�����W1=��l��$r�Ap?g���z�dҺ/�DE�u2�c�7ۼt{�\��f�d�=N��������V	8<��Tޏ���=/�7߽�^�2є�����cwa,Y��F����Sܻ������ϊY����w���������e�������5FF�UR�����@���%\7df6�r���f�&�wE5�Y��
L�Z�&p�s�f���j7;v�
p�wm>�3��	��Y�\^^�w�Q\Rw;�"�[j�;�5A��g|~R"���~�a 1~�����o~�����{r�����*�%gw�����c}�p���?��_
�p�Ē�fJ��:��|coNK�C�SJ�%Z��X�T%����0��K~m�3����L����z��?���#<�>F����C�M�OTbӢ�O#�IGbd>��_bk5���
�]T�U�����ױ��x���k�k&��t�w1A��1����3�+;kW�'��P�E!�����Y2�1�Ѡ}�x�h���T-��0SW�t}��Id,�2�#�J"������/Cq&��f�g��KH1���{�����>����Օ��P�<��A�g�LP4���qR��Z�C �k����� ���3|�x�ݗ
r���f���Q4�!��nM%�R���D�k���sQ2�M!���c}���w��#  ��/v�{x�jW�=���	�]A�/a���J�E�w{Ѵ?4��g�oTk8;9�ݲ�䝠ey��d�a��JE���`lBp!����H4K��-���g��uF��z-R2�=BǺ�\k�黫���L��ޞ�ǟ�F�������w:��3��2�^U[��TQiT�K'Q��g0W�����U������X�{1�]��*�\Jl������ۻx�j�1�o4�X<�d�`�?�z?���/#�q4̉_]׮ٚh�4�|I��R�.��v�X[��^��������>�eM�Ȳ̊���`�r�8A�<?�-��H�����do1����+���rIƫ2�*Z��bܪ�`a1�nkdg\Q��9k�c�IdL��1<�J��Nѻo�>���u�5^4vL���?k�ŁA��(�f��_?6�$y��z���A�Q��x掎K�˯O#�?���(�3Kp���=�dŠQ�nV�g�(`�si	ue�~��'���1���5bd*��ȥ��H�����ˢ=$n���Tp�����cie�1%n�I���io��p|QCK;ᔣ+����[��ҖX �TRS�7:n��h���'�
���	�	F/�͜D-�@ �>�v��^q{:���dNU*�B|b�3�iW�������==85�2m�FW�E��Nae�&��tݼvZ-7C������)�>X[&H
`f�`�A=��� 2G3��ոq'���+�m?�E��5�U�͛Y�gy�ĭ�������xڪA�N��m<�S�l�ڨV:ȯ&�0[��٩�\l���Qު�4���byi�@#g	���7�.�r�� X�������ޡ��I�@��:��Qi��^��R<�@�{=��E���SQ��T�+�z�_�$�Ǝ��� '�أN!����g&��_:��
jpX�VI`['�l&L�s�q��o����!�sb�Z�}ט �&=���}�}u���7�)�+���r�@�܇�D\� I<���	ψ����x|���1���Ly4˵�����R4]����������8u�&P%]R*M�:{V50�0S@� [�;[Kx��	�F�h/�|K��s����y��a2��H��<���`��E��l4�m�;�T�AӟC�t΄�?�&V��y<5�E��Q�y	�1H����;�y�u���M����/ЅJ�߉[��@���`��(�C�0߻1nnmX�����.�>�@��\��|i�����pgs���Ե`�
oLsu�5���3���Y0з�upE1���Eg�:��9�G0����`��Ǐ�x���,Y��60�h���㌃M��gG�]]7�V��{|xL ���q{�h����޸������o�?�w/^����B�I�L�{�U7��3)'�
��G��zK28���y���_�T�c�g��Ox���;K��%������Χ�I6`r�T��^��Y���l�@���H�ى����ݿ�����@۝ұ<���!�U����)l��G|~~;����^�Ta�͋_��S��ي��Y���<@=ƙ��s�kD� �U��s�䫣#���W��3(&��_Σ�h��یY�&�n1i���M��hW�5A#����6pu~�o0������&h�caa3sy����y߾<��I�&B�����Fj�<�`��F���V7oc)?��~�5����T�����Gܟ��ó��3�=�t�_��٣��*XLb�<�} �g�{�ժ�f��o'N�]��Y������%�v��r��,h�T3��|eR9��2Y��L_�-�ɏ���U,�'FoG]���1n�?y���w���%I���kv'�ٴ�b�͛��.�1f��J���N��w|�hp3�3�z� ��s���U�-����5�0�,��������l)�iu[|�M&��?}�ܴD��XL�dBfF�j���~�����#8�io���Y�\G�0[��������]�ZK���)~��_��;^b.�kk�IP���nr겞�|7tg7Gv>�H,�X��Sޡ���X���4�mđ)��j��z������(���(�f�'6C��oc&��l� ��VQ��o�����!�Vt��������O��ɵX�[ޛ���~fz<f0�X�5�riV�d�"$�_R�I?)�Q|��⾷X���񦧽�.��9��`_���tW��}�'3O�#�-�l�TC#�;Ĉ�_������מ�4��z%�x�ҽ�F��t�R��9��_4\)d��*�A��^Kjպ�WU�]�Q�'��o��\�A�Y��{N\�To�TOlPz#^�Υq�k8su���ܸ�.�4��,i薜��ًr���B�ɉ��_C|&z����iVX7j f��/-��ZD}�Z�wf?��Ţ�5p����]�I�$hs��x�����ڇ�z��猔m*�x�'ƌ�rt���0��a��k���}d����GG'x�#�W7rIzaŞ��(^�l��LzE������!ߠ������̋��ln�H
q�VG���K�CС�y�%/.�q�X���,��H*���k�p҉BB���=��Dgwy�B�;�ܑ�a��nGm���$
�Y�rMy����6�y�?�k��w�5��mrze��g_�����eI�Wc���3�{�p�K����OV	��R�)�VWN/H�����]�rBm=]F�n��41�ڊk���Z�1�^OMqhkQ2����@�i�[#c�f;�,Ԇ�]�h!���$�x�7���{KV
_�ە�+�u)cV���y��%�����H�������֊��	#�S%�Z.���Q�Ԃ�G6���X��\�X�mc�N5g6���
=�N;�=ɗ���q!��q��3?�Т����������j��p�5�C5�4"f ������S�7.�"6Sq5��S�َ�����^��GZ�Q'����`D�Ѻ�n�86^���M�S7������ک(�h�)�+%��Fɿ��3y��9�_@=\&xI�fK<H��PLn��.�QDb��m�?E�(�0�dD��E)��ȣ����dAI�����M��L�OzNf�1T�i���K��_82��f�;~�� oN�zݦ�X��^xRvvv�le��g����_�kW/��q�n�rRy���(�P!<ܴ�1ѹ�i4���z��6T]�;; 
J�^dsR��䏟?���Y�`�c1II%� �OG�,b]Z���儚��sUe1r���x<t�㟪4}4MP������������
UuK��W��2���
���ˍr�Z/�H�``O�ܐ�y�̦" (v�Y�t
�.@�Omܨ6��ޒ��"��>�׫�G��}u�EZ�B��",�8�I�j�Þz�����LFI�2{( m�a��~O�uU^KF�riuI;Q�nm�{��B���o^H�5�&��P��,����Fp>F~/��[����p(({;{���Y���xf饭Է��8,�73R��ty�ٍ�� ������99����jP�ւ���7���S[	���j�Qy�S)g�K��_�D\���j�Շ��蝍'"�,q�E\Ju�Ą^M�HL�k4x_�[�Q��#ew��xq�$P��;���~&J$�{��\w�	){~!/�� p`9���P=8����$�y�H�sy��U�����(iQs�g��{�=������M|�8��9-:
Ş<xZ�g;�\Ֆ���!��`�:��q�LtWЃ�Ѫ��X޼uE.��I&=Т1�L���"yPX����_Jw|v��˜�3)i�2UO7
&1����w���� �5�H�D�$=NHs�paCw�Gj�t���8�tJlT�h�\��ܿ�N���#k�6�b2�IK��e,v�0�}���%��7S�����'�ǲ����k��ٺ�0�&��O��峇;�Z��,�M�|!���#��y��' �R
0�-���lK�1���h�"N4oU�'��p�d{5ƶq�ǝ����I��I2�Qp���c����]4d�O�?����ߕf��b*�C�^v?�b  N�#��,H�d�`mQ��h�n�a��\��yCz�Eyx���QOKR+{��ĲTc�Ӊ̆-�gf���k�_�\��&��5=t<v��e�y�Z����?����#n�Q��*FA�n�E���iyP��ĒQ����(�뺓5F����8�iU� �=}�Tv�Td�����2�� o�ېG6�<;����|�t_���'�r��?Ȼ7/�*r���%�C[j݉Ҟ�p?�橔k-g$�Bj�{����'P�Wr-U~tq_�����tXE*j-K>�ʓ�Gx�i�H�_�I�L)��Sȅ�~�s�>rO�V.�@�7��J2���ۿ�>����RM���Q�}Q�E�֧�Gw`k�E�GOj��I�L�X� z�^�ҷ�#�=ѝO�-�sEa'K5��ʌ1�n�T��?(�nQ���]k�t�'�����g� �_�O�*����ɇ,>���t�
������3VG���'Od.�67#�./���Yi������$_m��YINOeخJ}.&�� ���C�|kKv�{;���\6��еˀ������#�\��d!�H�$������\�����E������;g8W}|n�o!Wٱ��ԎF��P��V-�����R�._��E��^C��FF�6��>�<�׷��^�qC�>���[lKy��+���h���O7��NZ���
���ޭ�G�V��u��|�Ky�.ǎ��k�eݱ�% �P����/���]垶����
|������	�z�4+Nw�e}��ɸ̢ȟ_�����,�:��ˬ4�x7����YT;�����ޗeqރ{5��BW���D1��#1J�S�d��6��>�Y?b�X	�`��ϓ�Y�y����C��)<S��{�͚˨$��JG2(�O���ͦ�*��R����_�h�Nox���ͦ-'I%N��0�E�|��s��u��E�K����k�'c;�ɟ��F����B�x��>;�Ӵ����rp��\^��;��������h��7T�Zl� w�����B�¯D+5���@��<X�]j�gAL�g��.��Fp����QYL#6.�**6��IH
9��h��).-�IA������R����� ��6����W���NU�Jm5�wXUC;=�!h9��&WO-����6^ѐ
]u�5�rG��优�� <<�+�����h��9�"^���tʨ�s�핽<�d!nV\��_�)�S*9�˄�]��c�DR�0��A� ����xJ�a
`�M�%��(w�,�����Ɩ,�]� �����N�#\�2�7�)�O�.�0.��/e��O�R,��˃pvZ:#�.�SX�\Z.,�tjvtX<�-����IeH&f�2Q�(Ȱw`xS�)���9��ĥ0xxҒG/��x_���#HDU�30���Ϙ�it�M�� Y�����SΞ�ɣ�;rxt��wa�K ����z��g�h�=6��*�J{]�t��������&`[�)�֟�4g3�=/�D|g�~���@g�("Rr��Mٺ:/\�.O�A]�Wd+"�JS��>O����^ wz�����T ȡ"��yImN��TU�I�\|o`� ��R����5��u�G����by����8��Dwj ���(�����T|iS�!�O�3�u�
�|(��m�!U��wU��U!�@�\^�gC����9m[�u��|.�g�Q�h=�����a�Ewp����T�%�U?�oJr�6 �W�T8�����H�J����S)=��ZS�i$~���Nc��dbǙŎ�8sG�B�N�� �� P�T:��������{���fw�(�zU���ϖ�4=��}�U��r9����{)J$9p3����4[�yܳ�H������)���ߕ�?�yv�*�d����[*�244n�ל��Z8��x �jM�g:�)s�s,Ov
�}P���"��m�&����-&?�"]z�iq��/�xHn\Z�7����ޱ|��>@ש�\�}O�^�B"˃GOq�(&JrtQ���Z�#6 ���Yh��FE�I�J�N��;n�C���P�G��F�5UArl�I�hZlP�9��ӳ2
Ԓ�]� >OA�ê}$�`rw�)2+c�|RA��;�C�y��p �H@�Q�d�>��=I�"�l�����-��=�B���+$��̭�ʍ�o��Eި��4�?"�u��5�}������k��dY^�&��[.*#y�S�O�ڕjo�;�$����bbj(�JH�a,�
%[�  {�Q��v�B";���ْ4��^$9����?����ւjh7�9���QP淍(���s�c[Ea�Ƶ%�yD���"hE��z��ܓPugvy�"��H}n&*
ũ�4QN���F@y6��i#��>��q!�G���z	�u��j�~<�^��xl�$��_ �Zy����I��~��7ߐ��3'��em����ܖX莜={ ��3�����z߸uW��ѻ��
���V�(�F�K�ֶ1h&e2������|�q2����b��[��w�q��,�����*���zu�F!O$��ӣgc���F��p �)pt]r��T�3�d#���i{u��%����-�C*h�������C,��+�_� �!�%�kF2K>�U-�(ۂ��)�b@��%�I�ۖ#PF۱�@����C��ϢE���X��R���+r�s�AN���L4�W�F![��0�� p�?�L�ʀ�e��jKțqI�\\��`ȯb]�.]
K�̉RI�W<�����K�b�B^a���ٴ\M���b$_<ؑb��7V�M�.�\!���������nuu�k(��YB)��W������� �fJ���� ������18'��7�2{��n �{M�@<�o�V0MH�s��{�*Z�:J#����y�mK��ŸO�K��%��Ww����<g&jK01��\��N��L��f��Ks*q�a�Y��Ǧ)�q�]/����!
��ψ��߻�i$���6�=��3��F*c�^�3@����>��@py���N#���e�DA�j�{�����/���Բ�*�|�l��PQ8��M�FXL���zIo�M��ʭ����<������L}I|�8��W�ٹP��u����R�Q���<��n��;ߛ��N�tz�E��a��D"�B: ��2
��u�H��o L�:,J���q0��#��(ߘ{���*Z���3�w����u����H(څ���� ����Q`E[C��a����c��K�;�D��.�Z��^���C��+J���L"��<#Ķ*�V����%Wi�ϓ����A�vK�{mmM��QW�(�'�	"Ŧ�-�}FD��Scs�t��cTZ[8�v@��<K�lI`��G��QP����嶭�m�2���cC�U
�
Ռu��g�)��s�*{��U�z'<�WT)��n�W# g�:���đr�޺
9�5]����F.������������@Cl�Q��D#
*��`@�+?��q�wI�{%��X���4;\�M��^Uj�^�Ǩ����c5Qp�q��^o��YUZCF�$����>��f��K��'R�6$Ǘ@ ͬ������;�����,�}p'���c:�.�p�#5M#���8�աl�t_� �b��? �;����I/�@~/ʴ��m����K*�^C�x����Ϣ�˗��woˋ��<AQX��P\��u5Y�	\����F߿�ȧ�~b�t���(<H������x���:3U��%��T�e@:�w���8Y⡬�����G��t�B�qs�Q_���m��8�5��x}!�!yo?;�Vޥ�ՉdLn�L��ڪ\ xP+_�ȫ}#I����T²�b��7�\Ͻ�R��,��rr1�kH�r��@3`ҋTqqb�K.�O��D�*=ܔV���)����)��Ge��hGv駄��U��6nd��\���ْ�ɣ9 o5*r�ʼ,�&Zr���{���s�l������V���Z�� `P+� Ep��ߴʬs���qt�E�N(�>2]K˩l�Оt��E�td81�Хr��SRj�%_~�X��u }�唄�~y� �+�k(�+rxX�_�<	-���.䏟��9y*`Iʻ�!�޸+����=�;�ݵϣG���X�f6�.��,�~�ǔ�u�9h���˗���h֔�<�l�Mo��;�W�V�\��Y.�	? 1��^^�z�
��.�0�M:���*ΤN�=��e!��|$���\���\��*��E�`3��ݧ;oU|�*���Ҽ4��v��5y�{|�,��$��V���l1 i=�,��K��5͊��.�r:�S�
������T�1�]���*&��nn]�Tث~���	#�-����!����>b�L*ZP'�^�v��'ø��d�81��z��}�О\&q.���enyQ�^[�|�( ֳ|������ i�D�}$5����yt���.��q��>�7�pbV�������vG�}�EHB��~OX'V�VW�	'61���3UKI�!3�c�1����G�����?���ȫg3�%���{�O��=r%�g���o�g���̤��w��wA�z4��_�������@[Z����+����)�[
�m�9�rr�D:�8�D'�UgTT�ΐ���F_V�V�,:�Kͼ��N=b���K �|s�sYX�(>��=�g%���X�FE�x7X�_ڒ+��I$hi������q����
����*eټ�&7V~ ��]�A<;;�W�v��_����ă@n�2��,<��kĨ�ڴ��
�׋[}C�ܾ�
�<Օ���K�4�����{'�*��u����� �R�o0
P�.����崴�|��W���EY]�������>�Ã�\�zW��:�?�	>w�WE�R9�'Kj�l���^V���dT֯��Ԍ;W�K�wL�g��@=V�z7{�� 
ݨNxkio@l2�P�eL�-����o�7Tsr�^2��{Xŀ_���4IYO̡�驘R�o&q���n{.�\b�{g��|��w��bZD�X{�/�ݸ�5�_��h�� �>���5�����h#��;M�ȫ�xZ��3�2��NLf���_��E�_����g��y��n�?��n7$�`\mLh���ClZ᳤:6sd�_P ����٣��F!�JD����F=���b�(nEL\r���4z�RH�ȹX�{��əߒ�zF��i����$��?�iK1Y�5�?�k�ݴI�ɉ��b|����ØI&duiK��� ��p��nl��q��IU�2m��B�R��$~�՛�d�;�������xkis�n��D�i&*��]�=%(G�A�/�e��BJͮT{T_Mh#m������]�D����<#,�ia�&p�GREN<ɕP��s�{Zd�����b�ʹ�e,5�Z�S}�\���q��,���'�rzt(�dFs�p��݈��j�[��+���ó�K��>�?�S���dQh�΄$�����r�DOƎ �w���=PE~����MUE��u&N٘���e�-_9QoR���Ά_w箭b��Ϡ���}�!ڄQt�9�U��w,ɘ�?.1<�h ��jYڸ��ۊS�	I�/��k����3��Ɍ7"�"0m��?cE�8}�b9W�&��c��H|����w�B���KX�;�����y}�9Uf���p�J�� �4l\pՈ�?�Cq�����i�Ϥ�j�U.����H�7{8�QEX��uPϕ�F�P�և{�VƧRB=]#�o��lg��6�	fO�E��2R&�S$̥���1�)����(E����x)��B����$[�4���/�ݔ+H4�v�*���g�U[vN8���ʧ��d;"���H����3�@E�Y�F^�y��QK��0���:���c�c�49�hd�~\
�P��R� J�of�(�,	���b��f�Z��5��r���ү-'ekc� �U&ei�<ꋓc�|��ܹ�%�<
޶������A!�ǅ�=�X���bʖ�n����wINن���u��u tڠFf�o�H��/��&w�fjR��ѳS���l.�iG�@h���ׄ�f��Eg08�`�RߦZ����|���cYZA�"������E9�u%[��� ���u+E���P��Smj�/�5�vtǺ�e�b�2�uz�_���V� �τB5D�K;c�������Ԥ�tI0�,C;`��I�E_ Ϡ�1Y�"�ܹuMi�xsu	��f�����	�W�7��s�p�+��h�����������a��{y!URc�>P�qU-����2���k&�N�TSl��F ��O#�Q�vI�jԛ��!aT �y��DJ-�h�B��V�4��A
�mF%�x�{��򪝗0n(H��UYx��Ff^z �g_>Щ8)��ڹd:����s�Bq?����9��^|�����.CqUJ�	���C�ٓ� 1r��B���2��$��G�����]��s܇��0�4vec�E<Y	�L,�PYa�G�������0c$y���8hʇޕ�ٷ{h�A%��|��3�m�,�� Q�h'�M�(t���N��V�d�t}mb�>7��f�X -�@X�3�yeQ�Lt��5��:���C�d&�!|���B4,���,�E?��z�L޼�#��x�w�H� ވ'�����H���
H��m�<"q��#��]��/X����'~�d���O��O{rgkC����%��_�f6$�
���P�H����c[Ey�ʩkC��܅�6���2T�q��	�=�ʿ���%��3�tY=���{�<BZ6;�|F�SK*VO�uuߪ^>F̙��}��<��>|g��Y}�s�&�5@��>����w�(������A��N��\��C��{u�^��n�ո�*�)��弖��V[���`�XL����7�N���T�Z�H0�h!���ї_��C�z u����w���goJ*�X���/�|��-�PRZ���]��Q
"�4�(�#B�wf&	��� �������_�G~��rv:��?�#|��|}��[�~��ɇ-�89�	��;���}�˫�dv�P���y��/�ޖF��k�$�*�l��u5�Vj�N��ggȥ�U#p&
��E�."�Y�Wjȓ��?�3��)����_���ɓmNQ�Q�崐S��k]\w��ʸk��S�n��x}�t��%�k�����Y�(M���(��ӆp8$�،��Z� ��G��&1��d�Bg#��
����\�ۗcr�Ӕ������ܾ��b�*�����ԓW�%�RWs�?�7�ޔx��ЈFiX���½�Z�!-�l����qQ*�}�Ԍܼ~��z���<��W'�,��s�0���l*Q��T2�V�D��9�4jrmkEV�(�Pt�S��y�"�w�q��a��
`?�e�P�B6[I�w;,�A߀Q�� �G�o��5�T�9�~��Ru���?�x<��~&�oߓ�+�hS���"M��4�ĳ�ÿ/�F�3������*�h�p����@FUj
�8�c�QΉ�8��@���gR�� �(��� ���9��U6�6S�D���Ŝ��ټ<��[|+Y^�;TQl54�r�bavAV��� U`�1�j��-e��DE0��W�b�x�Y�,k��j�3hM$�Ij�]#9@^�"��D��3��*d42BV�u��=�$�
y��HZ݁N��jy�����Io�˰W<�|3Q�t{�!���ͣó��;Y�\W/]R��V������_O-Z<^mr0^�`��[U�;��XP*z�D�� ��I��:}�Gu!�q֬O��y�Suc�4���zCTXF�?��_cA� �K ��!e����'i�{�b��(K畔� �k�V��,�����vą|�!�t�*(���%���-�BQ���)V���G �݃f��^�a)�4r9C1"�\����"^F�1|���ړ&����dK��}z�Ҧ�D}��:q���m�Zb�aǤ�k�`�Se"�x@f�W�
�>� �ɐP���sj�=���1�w��D݃��C�DHז�k�,����V�6�z&ʫm��� q/>x?
�qKv����db�>	ǂ
|�,]TÜ�پ�.#���Td{o/�XΎ�(>|�L�(�4��j,��U�X��JG�?ߓ�TDf3q� ^�~M�� r��� ��s�P���ȾO�t�>��tvc8��g$1� �[U���*��ّ��;i�j�QInq(�b�4�M�|�c�0���Y��>=�ɍ+2}[�J����f%м��$�_���#��\�îk�~�&
���&���P\<��#�{N���wRpȳv������^F�m� ���e(��rґ�]B�h˓'/Um*����l��p  r�1A��m�D��S|��Z� RCP��"�cI�/� �Pi:�ܸqU>iT�J����+u�*ciDҴ��*i���2���F��J'����C,�@��0ţ���ž\Z���MJ{�Q��F�ę���+�u�����I�$�}rvr"�V]fba�E�ȗ$���<6p�� s��S�: ,Rޘ8�]��#�D�#� ?�LX���7���W8�eR�
V�L���n��i�th;�2�CI�z�m�}l�k����u3���?�gc��R�W�VU,���9����1�׳�����H�rEZҟ:�v�\_~Wʧ%y��
9�Ga�~":���� I�mf?����v���2@q�R�3Q�B"����ɫ�|���;Ź�I ����s�����0�d��vL�}Y��8(N�I{��aVv^<�ツJ�߾}G��7�ȟ��/UU��İyu�SƩ����M���L�`�D2 �[��K&t�ƍ��!.�5�>g�z� ��E���,�8�uU��&�(Q=9�����Þ�??���ݍ�*_�6��i��O%˝���jfFJ���Q��[<{| ���#M�1ep�u
����(�O�r��QʞV;4f?8��7��dW�/��~|Gr5[~��39���ER�a5���C:�fK�.)�FH�xw�Y�L p6; R#R�qIհZ��SA-Gܪv�|B���G��LwM8����Y���.���/p�� ���[���O����D� ~���ЧMGJu7PLUP���H��.#��蕦.e\����t�$�)�S����0���h��� �E��K��( O.���ƊGj%K����G
�y� �#����Т��͛2�{K~]|�S�@8�xc��^U>�ݯ��Nf�G1�BE~�ӟ��ʼ��P�.H)�CL-�˧���g������F��[(���(��`D�����;
���L(t�b�çy�B �R���{�Fj�%˯���3�e��5��ۦ{��kbv����`��ʐ��l,F��7ȏ��+uy�{$��^A���}��X~b�!��E�������WL��g�8�w��|*��2�פT����չ� ��0�s�8Q @��0HA5���|�y3_�2�#�O�C׮m��ͨ�x�[�UK�]�s���AT��H�bڐ*� O�J�V�qxx�/]C��b�w� ���q��� ��s��Ҕd$�3��ӣ}m�.��Т�A�L�ORY4w�f��2��(�v� >�3��F��ųJ�Ԗ��,pb2-#� �<����z�]hƩ�).�lX�w��[�G�E��O~|O���YJ�����w�k>�m���kl�&�wQ̎_��/��H��Z9�3֦�e��N��[�O�AGY[A��!�k�X0����񋓰�LL}9	�W����k�H�H���LY.]ޒY`��|﹭�%B���'ON�j�"8T��Xz��weUi�2�Z�X�(�W��z9�L���y<k6AErU)�}ڜ��Tz�Z�-�NO�[,���EG�5|� 6�I��2��.��5T�0�Ua(1@^Q�z�:�u`D���8�E��t'�!6���<_�{����4�Ԟ�R���j3d��έ=!=����z��xJ7\��F�F��m|[�:\��>ߛ��ӷ��������u�����%�̸����W�(~"����xz}yS�W��R����􃓢4���k벜���|(���k���P��@��kc��9��n/�쵍�� &Ӧ��<������d��U�GFk%@�e����x��?��nd{�,�ٲ�e^��Ѹ=l�r��q��eD���\N*b,i���J��N�R�"~�����R�,�\�3�(�}�9��ѺAT���h]`��|9�*�xM.�		�������URE^�L#��랎��]�̾��k�o>�@���� ���XR�>U�ߎ��{x0�����
��#��-�.�o�*�T٪��O�Ha��$�>��s19`���$��q9F��A�����}�>�JbqQou�L<F�]�/�l-�py� ���UF�GV����q��-M�Kr������� �t&��KA�ǉc��a��+��`������g2h��T��o�������ߗZ��8Ë�痭�R���Kpx��R,�e��4� @`��5P���PF'�twx��׿^맒��3���;R���C5�]ǅ�u-�є��kH>1�qs]%�]�ޡ��ϗ;yɣRz-���ަ$.	�JyAH�k�W��n������}�X���߻��X�Z�%�XK��7[�&~$B�v����n��c5��3tH(�Ԭ_w�� t���S��H~�6��l$��u�`l�-�1S�>��.N��*vEQ$� 8�(��=���Y�r�
.#}>�E�� �HH�f��5=��q{�����R���d����8�ִ��1C���p�d�����9l�z`�SՔ��~�R�i"���.�鵫K���9�x睷L����]��2
����]|�����L�TO"q��q߰'9<�Z� #B!y�pW�>���Wd���*]$�{ϥ��H��TCUA&�#�mUC��@���D�n ��2s�����=�Th�J<��~-M*��=Ş|Z�6F�8;N@mcQ���J�(^�/k���p���]�VfI������H�hls���Ő�=J���zRz�����z�ޱ��$]�?��ޙBo�4^&ӗ��8�����}-��"�Ҵ�c5�x�.�J�9D�]�����}��\�vU���&�z�"�TJ�݊x#cYZOI�	@�f�fi��~v�����]5+�,��ja�n���3�D��Z�p�X��TM�m�U]�yf]##"é�{����|����>g�PT�و{;�Ǣ��*N�ܖ�wq���N�\j?���괏V�;"�%��oJ(���#��o>�9.˻�#��gR�y�������-湎��&� ?#�}�i�р�!�7��a�9Bfl(h#qzǜ_��NU	���mm�p���ϟI�	�)��3���@w�V�����/r�҆β��������ᾄ�_�.\A|�o����7��~���
��44�I9;�Q6$ d�s1R��h�����?hN����b�!_?z��reDX>��N!����v8�]�&���mc�M|@�9��,��/�X#�XA:	�}�zTI�~�P�� ��:�ST@�$�rtt.���y����.����W ���˺F0�^�?�ђ�Z�} v��J���3d��|EVE1�L����,�u��.U��G&Nr��6]����\9�{jD�^�hP��i���������Դ����u�g�~	�b��Oz0
��_���+r��uYA1Q*UԷ�e�?�<�͗���qU���\��]�7�ji{M���9hRYAm����Ȍ�dy5���'/_[F��[�8��!E��x�C-Hwg���b>��K�V�<�AW0-]�����<�Ě�9{#UC�8��ƪ�2�YB��a�bv�P�Jѥ��I���Y�?ؓk[����>���̤�_2J�$��C��m3y��zw�a�{��N������@��T�Z���h�߅��*�P�:㓛Y7WJ�:��������= �f��FmcM�R1c����� ��dqeI�i�?9=���?����*� 8��#�D�7���;oƆͣ����<so��{��,#ą�6�l�ǰ�F�ߍt�S��f���/�{��x�M5
�Q1_�x(>�,��ӛ��y��R4�e�x����L�i"85ZY\Z�hpQN���G�K������{V�����_��ڊ��	��IG�i�Ј���]ln�r��~&�o9;��t_P��_:-j����.e���m���BXj՚��s���r����&�Jk��Gҥ�հ.�����X���g������;�3&|�b�$����|���_++�|�A��PO
깬�q+������6�[\x�6
����E��Q���F}��Y����Mc�E9��9��y�����p׹��4?#�s����`�BA�~��Z��Wݍ)����A-�R[��L�x.q��@�\"]^م#G���bЙ�������	*X�]�qY޼3#/��ȋr�ƪ\���@�i�Y���5�%(�>d8ꕻonI��^̢��V}��CC�}����0�;r�ʬ���m���zqe�9T�9�CqX���o�tS��S�s�Ă�v���%�p`|�����3�)���{PʀNCp�CIp9����V`)>��e�h����U����T�T�w�6we2�>U��9if�P�l�@i���w^�n�H8��81+-T3C�H�Չiq��NƎJ�ؙJ8 tb������S�,Hs������y	���.��Ç$�� O%Гü�p��Q ��Xr�=�l�v�He �<{��Bۯ
�6�s��*�8">����}i�����m5�������./��ZB��C]x��=�i4O`�g��b2t8�c�\
 ����U
�_���#�*'��<��_e�|��^)`a���]O3U��q��ҝ��;PN#�߻{]��|:�"�aDG조K�4�̍	�U!TL���ʃ��KǀH��(�%���{���9=cGI;LZ�:Ş�46�4�֩���N�6�x������,��������uk]=.�cGnz��U)w��	 �����|7+��m��ʆ��B�EZG�jsE�W��w|���Ӫ�nQ޼>�d��������/����g���|����ŷ��]~� wt���!�oD��'�M�^�r��Fo�&�!�lxF�b,��&�5���Q4���O��`��N�[�^��ȌdueMF����� �����g�K���ظrU�ݱRVE��
�9���/�z 8�.-I��V�J��?
K������*Ȟ8���<ع�ή����Πzw�QEJ1�֛Wdc%"{�^�M$�����K�O&Zd/-�K:��Na���g�Ҡ$G����H���ݯ���L�6c8�Q
�����PW$�H�O~�C��@B���5Ψ'��Ey��#������c�*U?Bq�q����0qk�ͧ4�f�xP���y{��pJ�գI�'S�)S���rΰ��w���f����*?x/)�\�I6��⋯J(���_��P��+ݏ�����!8ۜjq�u��Ǐ ���~2�[��2���)�4��2�J�C��=��S-�?Z�"@<�u��ev��K'�ً���~y�;��c�I��o�)�1���CD&c���a-p8I:��ʓ�	���?��W���S9ƻLd�[o�����ZRi��R���/~�S��2����3pxr.O�w%W'E6$�(w����G�D
����1^t������) �M��H�Z�����e�����,�TMv$f�72`C,3=t;������T��R���1p��u�,����<~�7�ZԽ��7�V��8;/�^G=��y��L*��3H���Y]�H�$Z'��gP�z'F��Cm�XM�0��z�&�.�r�P�c�ц�@��ὒR){� ��{�DL�!���D��;����ũ1� �5�:��\��)�S6)kj����~�6�[��L%���E�O���C�W���y�M)T�(ֳ�M���sWq��1���-??���&_-��|�0����s�Ѝ���G�-"(�5���� ?�(�B��I(������⢄�3�������񣗲0��=�;wו��TE�S���8��elq��<�c��c�U�K�
Ɲ�|�/�5Tv
�`޶ci�=�A�f��IE��ܹw]��5=��(�Q���x��/��qi���6'��b`;$����jɵ�U�J.גr��M�KW%��b��K����"_�Zw}Ɲ��V��՜�)%�R6�-���H�QQ_�wÊ��`��Uy�g�*��u�ύG�A�S�2��ȃ`�8ϩUg3�/K$� \�Uۈ<r[�P@��-��T*#G'Ei�Z��L��O�i�v�2wi�{������@0�m4�~���_J7�(�-&W���a�T�P4���Ǐv����)(3����8;>�ݝgr��qF��̕��!��|ϫ�#�̺6�)�B�Ć���#�\s>�׉6�m�)�٤��(��G�"�k�q9b�������|\D�c����ӝNj"P�� ��['նͽ��we�t��<29Y��A%�*�sw6&�++� (<}\o��y��<���^�CC9�2�v��H�U$��_�)�?��Y���>���cA��n�vU��vk��y�>RK������Wp�����⇲��Ԣ
g�:i�2#�&�Sx'�;=�T2�Ӎ�lI�j��� ��u�N��'��������I�ݐ�SZ[��B@^��ώ�  I�����YZ;a�K�k���z�;���*.�@�ͺ�WQ��{I[�Ԑ��#��2���q@�*t9��evVÑ�v�~�㛒���B��� �U�7�8/m&&a5S�=ZpҔ7H#{OX�ؖ��U{Rjt�No�kR�kK�'����ȰO�/C���L���'�����n����0N&#��bɧ���GҨ��r��5�����oŏg����D"Q҄��-�<ۡuk$_�H�,����d23���8A!��n�����D�pRvy�R)[��Ԣi�H���[��/qY�C�H\@��jm(_}�X���,��Ni�n^K����N�6P�Aib�����C�p��%E�67�d!CZrH�_h𸲕�'/P��" �=�K�E��Gr��>'��^ۭ�!�0�b�($�J�`. Ei`�̞ )b谓��$-iS�E��s��,���✞���恜��J�Z���Wr���YQ���gr��=����6(�(jzx~^|�P�'�\�S���~�YV�i�n��qo���~�;����d�	% �Q
��:(�j�I�B2]�|k��ـ�;�[��r +u|�b)/C���
@�}�h���e���y��j��TU�h��.=k��*>M{�DV�w�X��LLZ�E��S��y�=�=��`,&[�������A�q��S1R��@}*5^�����$�d��������d�����ͮ��Y�N�8���F��  �-|_G��Y�[w�PTqOv"�'#y�b��av�O�;*!O����|��WR�lɭKkr�VR��3x��W��ˋì�&fT `ЮJ��ӣ#5��r[��E�"v8&��Z�X��T�B�PG��F1��.ڃ�l��X��R>?ρC	e��L��ӹ�H��v,u4n^oh�9�s���%����D�/�ƛsr��^�n��n��EW~���h���=
p�����+� ��^�i��]��� �(_.���zm22]o�t�GHe�U�ݸߤSɏ��6ŏ�%�wr��ޛ�4#+s�;"OU�k�ƒD���u�f������ʌG������?yK.�Cd����C� ��//��F�}�/���U<��;�E��#���3�*Q������{�'��Qac���I��gGAQ�p6��78j� �!3#�;���9C�V���ש(>����4p�.m���w�	]�����ѳ�|���?�+������>� �í��h�쎍,ŭvW'�T��bfb�AT�tjA0}�,�8�g6v(��Ϻ���7�H�����JӍ�&�˟�E�w���r ����K䮱��꒰ue�zNX������%���ؖL�Ҷ�x:�r���3���w/I&�Fi$;�9�� �r��4��F��*�i�0Dit6�h_�;�2g��u��Q�⽆b�g�MPƩ�<#������6+����W1�6O��@��RR���ū�X[��%�}����Z��dVd���(��?�S*~j.����ݜ���$
�y��I�W�󑙶��2�Φ������ rso��gM�Ü��T��㞗��YYXUF%�i��T�#/��>�"'�U(Z��X(�_�ee5�,�D<F�$�N[��r���*�~]O��(�ΐ��jVeg�g�#͞K�q<3�P���u����WyuU�أþ#"���C\r�8F����qԀ�hg,SWFC饨1%Y~�U��VT2�K��<ʮ��#9<�����_�OMk�����N���t8tv�]ڌ�
_���?1;įYj�?M�F��ɪ{�66�ec�(T�mrEѹz�F�2�
�����3�T� r�k�x����*��ښ�y����;%uK�>�&0���W$3�h�G ��\_� X�Łꎸ����x7�F���r��kuj��YE�\y����"N�׭ހ�Y�R� g�g<1�G�M!�ƚ��PuI��G��0����/�`cm��y�3�<8��O�FÈ]rR�u$���s�i�B�'G�涁ͯ}��� nq�)e���0��ԋd:�����s)���TkY�!(�\�o?���Y�rI"�8�څ�,ݴQ��ϣ8��ˇ`�L/������q�NH�a�c�D��z�ȥ*A�xT���A>��������Wz������g�)/�f8 $��R4I����ս<�������pc�m9]��9,v�ը�ՏdccN�[A[~���u�8�b��v4���>{�˭�F�8t*��j ��V��8�#��51����)�s�X���ח6thN1�ٯQF��ץ��6~h$4)�)�����P�$�˖ �����r����zH"\��w�X�qh�xGm�XA�s�ܞT�UY̤P�$��������WWeIq�=���vm���Q��'C�c�!驆;�Tn�z^�!���L��Ŋ�9��K捄qV�Z�P�c20�i��Ϲ)��<[w�&z�,孻���׫���z^�g?xgAܳqyp�K���߉ge��: rX�����! ��x*Ӂ\}�H;I|�*�3ᮅ��T����,��kd|#�/�Px�,�2Y�k�1��C������R_��`���Ϥ\:���nS" 0n �g�����\����q��:�!wx�r���mI�������.w�\G�sI��E��K!�ûE|冬,�I:҅�2 �o~�Ro�H�6�PxN���0�j��d��ϡ�(��b�Bp�o�2
���F}Sk����L{����lZ�K��4�t��ɫ�#�Z���BH>��y�����F �s��[�J�ؗ���	sw�6��$A��&����{5���F�Ӭ)�}=�������J���{����^9+���ׯ�q�q�`�C�v����Ύ�f�j�K��X4.�����J�s.��~NvYق���Q^�o7���=��������$�G�����7�pK��3y��Ca�8�;fhFF:�3�wb [@ހ�Y�7]T�Ŵ��w
�h��k��]�6׌��dZ[�沈�J����`6 ����K9��,��i�u%]���9�D�Ր ]1�<BA�@�b=��&��?�1;�Tr� fl���a��$3Y��@)v)>B%��?���H��K�h��~c/v�q�,�s�#>�-y��X^��/�Q����� �JMc��*������x%o�ؐ�~�@�w�)/��嫧���1v�*��Wvv��W��K �?��_�Zڐ��zv��� �Z~�aG�X����4������0��HPs�3w���D�c]J3���3�aɸG��5�z'�;���M�����R�I��q�*��Q~
��-u9�"K%I���x�.���34˨Cz&�%}���zc�/����v���ph|=�?+�ٝ���ͮ�Ƹ��d�^�0���x��\N?��kK����d��PB�p�-�Y>�l���g{#�po�1�CnU��q�Q8�[��%�Jꔊ��;�^�\�+A6���^�N[�Z��)	�0%Ã3X�קS
6�9壧-9�f��Ѐ=N������P]����D���q�TAw�l�c&�}u�r�U�-�� ]N��5HI$�B5�f(rI��We}}^��(k�?/���Cݭ��u"(*�8�g����z�X��z�b��j�����t� �S6�L��|o���Lk��8��r&^���������%5V�6���y�����|�EnR*(�È�4�n5�j�@+��9�ӣ9;�{�E!��(H0
����	w<']YZ�I�j��LB�e[�͡�pJE<̀5�&�K�6*�b���I���A���N�&i�\Ka��T`��rk�;4�8�ɋ��
���o<��j�C��b�(�g�����ŏd��!
C���6Z]�,��G�C�b&�!b�i�I�E�c���w�-�%&fJ�xc�LУ;��n�C���F��LB޹wE�^I�:Zȏ���7���� ��y���+��PΎ�.�Z_���}>e�c�&�#�t��3i��ܔL�%���EQ~��O.��0�����;���3�B|d?G�+�<�<��zK_�*��Bݪnk�+A�af���kz��)��i�[�zgHW�u�r�+i�nq>��\+(�۪�����3�.�j���644^�_3^Qop�l��d�O�N��']�(ۻ��>��q�g��:*
��E��Gd�\B��u\RI�3 G�}�H,��!
	��H9ߐ~s,k��R[+K6{����Wo�x�e.�א0fq�y�\�Xċ�>�����9��l	u$��P_�8����)�-��� �5i�X���h�K�� q�x�qab��b�*��є=����9��Ҡ�K��w(��o��ZH��fO<����issM._� H(�T�W��K�#�`�?4:����c����G�}��=Կ��q�ɦ�����|��f�ڋ�ˈ�^��R�b����*o�}I.��W;����=U��(�Xl�`�;V�X�d$/�t�FF�@U�g��,;�Y>��y��yD�� �!�N��;(�q���c�.T��1��2����r� �Y`p��q�!M�ݡ���'=VQ��>�>�Q���,��I͠�����Gv��q��re3%s�i��Go�A5����]|��s�C�s�vzqFV}�;�|�C��6���ӹ��.��M1h�l��7�x)Mmx�]���ɠI�f:=�s����K��xOJ�+�����UC��Ew2��<�"�B2sk''PJ��|�ٹ�7"�w�P��:��l*�B�BUj����^� ���]�Z�;�u���^��'/T�r��ęI)��3[ߏ[A;�����Nӎ�!~T�Mc�����.#G�\S}`i�X'�C'�L����w�R�+['8�cM�z�/
Y���m�n-���ɕ�Wu�q����-���W�y�D��K����ޑ�B KO�F�+�hTm6x�zc`���V��&e�f_����L��T@Sҕ�]�ׂ���z^+){�����P��0��P����8��)&�]�3D!}Q;�k+W�[w���kMT�̳����yI,�d��3e<�ݤ3���rYB(B� 
�&������.}kF�lgls��1,!��<���H���p9*~�R��[̥��e����M����Y�Ou���n��v�1R�N�ٹU9B���ǏZ�G�"�����с2>��{�W���}�l��XZ��P|qu2F�w���p�-�R�8����2-GTO��ӆ�����c`e�ݏA<��� `>y,r%�������	�r��>����\2��8�ͩ������[2��F�������x��X�.� G�Ցzr�uoM�(6s�*@QT����ݻx��rzQ�Z�纯`@}Դt��m����}-�[�!�ل��7Y+ 4*q��g���`��骡�)|e�8,ݡ���#�����	J8�8SE�N�՞NA��I�/����_��ܾ���m��_����6�ߌLP�5)׶�1�8lT�(����j�29t��mt�Uw���޴�'���l"����W3�(���/�e�@(�шT�.Z%�����r��K98(�5��s��p���1;�\���_cN(2�0w�)�hR}>;�5�G����h���$�p(��%�9����-�ų��D"6c4;B�U�C�t+�p��)A�T)U�q<3���-C/T�i9T��P*��锡V)"��5��y��XU�=�w������^'��Gc>����t�S�v+��+�_��F،wv�f��<v;L�v�N#�&���B��Sa��I�[Ez}��׫�С������fov��{���`0�Eq������l�n��lT�T
��ĉ�DΥ�mfd�8����~�\��$�)9;9������|��ή��K�myﺫv0~���!Er\Jܐ�����*!E�*�E��.���4�����7YY�{�����*`�!kX�FWU�˟���sN/03?/6i��'O*h�K���;�9��N������:�e�(�ń������)�W��>���^r�,���0���	%�TG���!�����\�����'rGY�h61*1�&d���j�B�E�{SYC͖������y����C���rL�5D=���`������K;E]=|�vB[�GH�
s
��$�%���Ha}���զ�@()g�������2�d<�cϨQ�����q���rR�\{ ^�oX�I¢�W�v�A-�џ�q�;%�^�I�5P��$~�s:�,��<T�Z�i��ﯣ{�O�]�?�Ig
%~j��=�(˾�7�1I�_�D�m���jr�u.��^O�0���%�,���G�`�hA�Ο��s���ꄽ��=m�x�sw��b�d�-���2�ַnH�����ȓV�PM�Y򵰒u0#/����Í�i������b�8�Ɍ^�I� ��N�8F��Y���/qpx.�/�S�dzZ6_ސd�*p����8�i2S���Фs�R�-D�%��Q�H��&��8�f��kB}%kq��Sـ&����rE��ަ��8�4~����F۶����ڙ,�a�|1�rNrj��d�"�����>�wY�:
�`+�r���ѡ�e��� �T�S�[��V��q�]NFer��C7���mI&$@�e���*���MT��)�ç��:l��O+#%	-6�$��C����)K^��6I��\�3l�_ ����fs�X��(Z�B^�,�etK�U�5��0+^M~)�S�Q�t��PPo�����.��c����W|��Q8�e�r*�.�DeD#T�>�"�1�����d
�~��T���xǧ-<}���mi9��f���%�D����8���ސ�]<�w�p�T�9ä3R����~���+|�0���	�oi�%z�S��^���X�CF��^����,��B�^�q|��[�|����*����y�J�<�=x�bއ��U,�L� qW���G�x����~���m���Э��Π���U��=nʝ�u��Y;A�8��3J��W��Bh���%,����ʲ�IvL2Ƶ!ɉ����1�t)���p�r]x�rFI�N}9�hR�_l�X���Ż_��D#������<>��Hu���$@)k׋��LN����U[!��.\�)���	����|߁���ϐ�(�I����������	~�ͅ�Ҷx�YЦ8X��ģttQ~����;��d$�Hb\��[���ك^��`�(�x,�����gb�\;R��s�QE<���%\k,�ɋ-���v禊�s�����JIu�ˋx��Z��q��$@(J�V1\C�jd^txG93ɹ[�Z�6BZz��L��*�"��΅吵 CF_����*�L�U���I�;�w��0��_�KY��H4�a�Գeg�W�*f65@�����&2r����{8<�JRT�Y��e����A�O���73L&��T��0G�Z&�)J _F�^�2�3�DWο�P��c�}�����<_D�J���v�X �~}7�3�����������HV��u|��)	z��$�����z�:��W��}$g�*	��Wߜ��OJ��?�Ke��L���~󷿇�������>�������f��S��� �R�Fp�Q3Ap�Y���U����Y,�&�S���3����^��ۆ#�b��������)�ܒ\���X,���0v�
�x�������a|f
m�����+�P���������>�>����n�&^�d�$(��E_�і��b���A_��R�S:��_(�Ԁ7ZC�S[RW�^\�����ܜ$M��>�i���8�-���jT���]�vW���3c@<����QI�f�V��Ɲ�vN�T�$�YZ���Ey��/$v"����t-�-3?&�Sg�lG��k�\����q���9^�KS� �)t�v�L�E$;$A�ܔx&J��M�����d+}Iz�m�Fb+r�c�wb��μ����F������Kyɰ��$��R�s&�IDX4�M�p�K,��x�����A]0d���"���t|��n�#
zS�+�;Wt@,V����i,�OH� w<��W����8�΍�X�>��yO�n�`X�k��LM����i��'וq{�nܘ��g�����*�rp���T��g�,���N͞�3
����7>B�[FvJm�3n�$j}��W��b/��^�M���d2���m&+(;f��ma��K
����y$.�g������U�qf*�ӳ��fb��#��劍�E�!�λ�wM�(���u��+�����nS��II�,�!B{��TƳW{sZjCxI�ӔX�T�+��{�ĲBevך��(�ѯ�$FQ�]�<fv�w�3vM񵧭"s#�$ڀ��i�yj�.����YyI��=g@�c:�:�"����[�L�w{ƻ�}>MY��)���4苀נ�lw=�����ɡ�����6��r���`�qA4�ȲR����<�(��	-�C��{�X�����c� DiWz��(���M�N�{�kD	:�x=l��XC!.����q�#XZ�&_�+���'[*�`E���t ے !���S�������˸uk�Z�g'��EֱJ��d��gb�*�ʦz6�U���m�*���1rn�Sm��+������)=`�<�D8��a1��� �1	��zY:w��(�ĭn8G�6�ԗ���鉡>ք��Ҕ$����x�����z8	y�\��h�#�*���BL6��\0R��aqW�
ݖ,vL8sh{b�,R��&1�B*�Z�f��Կ��9�@��7��"Y�����%	��0�����C^���D���_�ܱT��k%"f[e	��(�{��K@���>��=��#5���LcueV���h_�MX�{��ǃ��=,J"M#2���6:�Eb�#l��J6OV/h0��K�L+��9���p2e>�9�ǖ�N�8�6�ي���M(��	����.W؅h�FQK�/��S����&���V�6O�吕Ѿ�վB9��M�sh��A�F�!A��P&t���ii�$(ASϩ2���QW3]a%R0��s��j������!d� t�=<}�JXu�q<�<�cy�nW���v���@�쀞�8�W=1Z���'�y���H@�5������w�x��8U�|}	Т�Z�����|�*�Pe)�*F�Ɩ��}�3�7 \��ije�%�h�Z���Ⱥ1�`��kطL�P����Ct���O��a���(,I
9C��C<x����s�mbto\��w޹!�ђ���ͭ�XU�Ĵ(�3�(�~O~O�!�a��pC*�Wk�I�X��|*	J�#"K]�6�LY�j�AZq�9i9s�zI5/�AB^���^ܽ��k���c�dr������Pl��t�7o'p��?��3c�!WmW�f�����7ޞ����K@d�U��"��8���j�*>z���E|��7�Β`��q	b�B��m+ܗ{ǲeO��r�䙛%�[uZ�D
����*I�t�b�,��\��tp�%W"��l�����xC��eB��ܩ�갚j4�5�\ɳݹ�,�!����	�_=���n�����G���X:�[KY���P�g�c��6qV2��$��h�K�>���N�]{S-tQ+f�Y���Α���Q�LH6%M�i���d�Գ��!��0&���xP�HKKi�/#���H���r����:�����(�5�Qy���=���[��7n�O��)�ƿ��s~�㟠*�z��k:ް��������z��Q�ܖ��� ��9c<�,��V)3��'��b���L�UG�B��:�$� �{1`��2�DZ�4���J(ݿ��ڟ������P4�F��:jUZ�=I��hPb����|� �������"6v�rZ��"IDS�j�\�&�B���]=��Æ=��� ��UU�L�(�G�m�p��l�Ͳ���7��BjC�P4�.��V�Y\���3)�LN���+a��A<�hc/�ǩ�Ӊ�fof��7���=�#l͈���;,~�;���IL���$jL��$��<�C-D��s�bc�����oab&���7���e�D�c�0,��&eM�� k&�AAe�	�c�Ä7�*�ɧl���iF�)�a2.�,�R�m#���/h*�Mɰ��>���^��c�I���u^W~=F�&�mI/��X��wy�L�����h[�MAa�:��n5��y9E]Gw��r��Y�Z��o���6x�|����,6W%�m�{�;112������2�����&|�{��BCM�����������W��b�D�w_ǲ��z��q�oJT6��f5Y�~����٤vb+񝱄�0q��
(԰��bb&P�x���nW<Yhd7��*A����Ŀڍ�9	Ez�Va�D]�hǸʫ�%�yj�]v�Mb��G5�$���qy����^>���(�^��{�R���PK�=X��ݖ[Rs�W|>J��4G��u���|3�ڒ��d�8K�2���M%G1�3�����A�Q_�ܥ��y)��cو��1�k~�X�ȑ�嬍���⡐�F[mgLA�wDΡG���qE�b�SS*�R.��=!slPmZ,��3�Ŗ�&*0��(�����d�sKJ��v��pu%^�B�"N�n�{&���1	SR4�
#�A�G3w��:YhI(��9�I��2���^�pTb3O�,	}����Um+�6�΍�@�&}^�CmOs���xT5+ �.�d<���3B��z����ٲ%;M�
�v  ��IDAT�f6q|v��t�{�ؕ 1˪�h��Ӓ���V�����i3s@ղ8�L&���t�1|뫫b�G4y�*SX��X�;��EM�w��	�T	����&�F���N�v(�m8���!�»�H9�R�M�vq]��Ab:C��|q`� @迤V�J����{��E��Zݰ\�f� �ymN�����Ŭ�*e=5y�^9d�>R��ߥ�����v��G6�K�`�d_����܇e��9���|~D��^/�|���q�>9୪�i`7�y�&��X��IG�����aiu_� �s�%u�
�S���9y/il�������u�/�K#��$����H3�q���X�������R��)y%��Q��: �S���8�W*foP���U�Le�㔷mtl�˼�;#-�宖m�w`���ڏ��w���Y�d��@�E	�*���(O���#%+��4.k���$ ��&�j*I���3@e��x��T�S�L�n���nk̜m=S^��#���X[��I�k���}N�g$���^Jp�LK2�#'	|�(��w^��������b�.�HK�ʍU�y�u�{�ϟ>W��o~�ʒ���>|�Z����E|�w��� ITk��]y��`B�'��%ӭ��;�ǙǱ�˻��/�gȍ��7l�d���G����ZN��MY1��u��23�Z]� .�׉Hr�y$8�$�0&����QL$�x�ʋ͵�G�XXY�Dz����N8Z�s&*n'v\�˚#WBC���<J��:R�8OI�a�j�V5d%�MD�27��Sb[�H$%�j��b�,�8�>
�h�I�م��pb~V��$��I	j�:�)D��B��rq\��nܺ�pEJ�$���w�ǝ�7��ļ��EUOO��%!�63��c��@�\$�fU�v�3�'g�(IO:;��z�*�C;�{��2���RYێD�5d�t'LT^��������cD�
��SɌ$[�%��~m	���}��n�o���.�?��G��Sc��|K��i;X�͎2�m]%�y.��i���1�qJ���!q�^�G%�l�w�TVm��?z�q� �cuqo�Y��d�cF��0g���S����"/�㓵�*�X��A�(Q���p\g>h�b��b{�tL��M-�|��b����l�"Iu$�ko����
]
ƣb��h����n�O;w�ԛcRؔ���5=	X@��όY���%���yn΄28��a��
��B�o4�=��{����?��~�`˵�$�ɪ��ے؎�2��;�(�:��~_4$	�oiߡ�m�^5����	��Q�Pڕ���Zȶϡ�}�K�U��V�M<;��-�h���9�`��O[՞G�|6�ks˘�`qZ���N�������K�PZy�M�%����<z��̴����ѫ7��u�&٨��N���r�,�J�cq¶��P�+A�w]�wDa��7 �k�>�<gKe+�s�rǋ�(痉�����L�/�1��	$��/��f���SQ�ӫP�:��N����`~Cao��7�x�*�aj2��;�����ݹ�����<[O�qF&�8��q�jI�d>c�ad�|����	�2��W��N��"�M��*��a*��3�d6��t�@%%�;������I��$8ݐ��8<���$�q����%��Z$��#;� ���Ɲ��t��?1���e��%!n�.���$�&��Q�o��̠���o�|�W;�^�9�+��*:��85���>��կH=[���m���L���C,��+�S�'�k"J���0�[N����E��Al˞���!�(� ,�p��$FF�x%q?��G�'���ɫSS����nTe����hy�jB:3�.#,};k}e��j���dJ4:�֛{��j�����QL��0����')6Ԓ��?]CQ�}�̔<s6�G�>C���z�D.Q�{V����Q��r�jH&�Z�&�O�x���!]���oal$��-轑�� "-����X��=e���(�� e��T�~��zɽ��$�"A�+o�D�4?�0�y^SyA�D̀��1{�vK93�l������TDg�v�t_VFU[���ã"��$�f���W���V�2���!䄚������r������U�4Q��ٔ�7��ޒ�Տd*).#�VL��<r^/�H����15�!� ��r��T�qn~��~��'��V1*N����o�}��B]עI��sTG��&�&j9�9p�4�t=����+����Ei,ܦ��IX%��^�A��p�9�2�Z��ğ�kd�k)��� �IP��H�4n���a��ۯ�xR��ª�Θ8��2v)�F���P�N������m�v���ך��!�h *"�?+{���(�p�PS�kŠ��z��Y'�� ����Vd�2��X�9�Gku~���q�!�%�葃�����(\�ި"��7~��pf�b����~����O w^��-�g�2����?���R�-Rd˙�4�קƀ�F��G�Oj�#�p�M"tM�������IĪ�0��n��f�W��wXW6��,�ǠPj����v"�T���$�ees�����n�����Y���[{g���P�i8G�\}g��5 0�/���s�@<CAz�B��8�y��>��r�d��ZD4Afl�l��ハ_�����&{xrV���m�g$��+A��X�����+_}/�?�`rzf;�����!��$���>9@�������v�IpQn���F�@�Sk{�Xq=������YB�%x�(+�L@H����ݴ�ʚ���_)�h�������]�LPC[�%d �9È���!�cllL%S����S	�N��o���yC!�Ֆ�}{��o0�N�b;t�
����ڶa�e��r�E=��X.�����μ'_�Ӫ��i����}}#��$H�����53��:��e�Il$%v1.Id]�����&��_×�zk�e�͏~�����k_G6������?��-��-������&~��K���׿�6�%a���2�#s��Q����kuP+�;:B� 6_޳Gl�?��sؒ�w/.�{�!?���똞�UT߳&ﴻLV!���7�>��c��}�{���g9	9��7�l߸�����RW��6~�����Ƒ��p�6! kˎG�m��\�@5(F�8��Ξь:�#���3l��d���_+k����7�I��Y<�T�u��^G��G���R5�a�{��JRֱ^�`g���V���?���������{��m�~+��#�M9��)l�1}`�_��_-��?����ct"��>=��g���$ �&Y�U�]ր4��V����>e���'
��|�V���h#�����uѢ>~��{Ouvo0�B�|ƾ:�o�ur��	���$��Q����:���q��;Ȍ������xD�� 	��y�a�6�oE]�ys���8;���ԋP�|�Y�1�K�K�ܭ#+���edd/G�M�8/��t�)qʽ�>S9�j��� �(R��(�n۸�� ��d]I���;�X\�{���J|֙�nǃ����oI�v���}M�����K���SU��?��`Q��@P)�9řˊ�-B����N��ؕs�`ynaN��1I���t���sX�N�ia��sWƊd<�V���kU\�B���yuo��L�1�#�����x��[��~��Oqpx���{I%���MH-�O�����+�_�9A�5Lv�bC�������*�l4dauqo]� f�m���3E+���ЬK��u��녵�N-�^��͝C,N^Ǜo.`������~,ܼ����m�˺3x>�屽�Í[�l$��Ѯ���|�:�1�ϵ	�E5Y�U�Y�	���Bވ��s�Nsj?+Œ$�5Y3�J����`n�$|#
��l%I�Xs4R=��k�9O_Gc]��U�'��״KH�!'c6��J\>"�D�Sqٷ�
�G�	I�(J�K��>�H���:�ڰ��:��/��=����P�^�c�otB����Q��(emIN=�%m��1]���q�e��\HB��Oi2��$�s3���U�<���}��.�6�0��<��/(	����=�9YR$b�/eO<F��D9��!a�%��E����I�o�������B��%�u(7�1���A,PFmT����G	GC�/������~ނ^=��`i�A�iTny�V��0��	$�a���"÷��,�ͩl^��!K�L|%+l�lҍ��@�G&�49W�sjN���Cv�(��?������fg1>��ak��(H�҃���$k;�����^�/F��9|��/��k�w���K���������m�l�7����u�t�8-��0��[j��Ƞ�?&V��j[��t.�î�$y=�̜����*���;�x�/�B$� ;/%q��VP+:`I4 F4�+�q_���^_~�V%�=/�X�����1���o�n��XP4�&�}�ta��*��t 		��k@g>�e�d�2�� �^������hT���8���\��(V�u�=�� +oR�g�~<{�'�SIxZM.���'ѮP+�Q��o|dT��LH+@�g� Ƽ:o�n1���yT�ݰ��*�Mg�p��D�Zn�k��H��,�4���S���dG�J���!^�p(�D��N~>��Ӕ7I���V���g��̛�X�t���E�J�c��.���'X������{r�k�������0S��A�6-��U�;��x7��`�^r��.բ���d�u���2|�+S�},`4�õ�L�'��b|zL+�;G�����[o�qɞ�%`���O_�������zF˥SY��V��
=Ji���f��Ȍ����������@P�v�Y]R)	�D���(�� �|^@��v�){Ǣ���H�d�Q�d��gMߝ�7p����
Sء!t���ٴ�w�7ɩ�Ѡ&����ؘz��Ý�^�ů�g�:�����x�ݯ���"6ֶ��s9��n2�w
�}�lQ�C����3/h"-�a\��&q�<�ǂ��,�jX�|�����ԴqZl��|lz�ˢ��6+Z�N�G/�w�b|6��]I\Y�==�`e����m�6O��Qk��P����	�(v=�`���O��B���х�ڤ�5��I���
��r(�s��$�J�gRL�Oa�.�
�R��{hHb����$U�z��1�����z�I�Tm����j�����w:�<��̌��>�����My�vc�����?�֝�w,u����z�n�������mc+h�y����b��e�ps��]C·��؞��ф������ûo&1����W�;x�|'<�r/g�L*�V�X����YuO_�cr�+�]�
��?ؖ`��%�{��G���$�I	PIP��{O��W$q�%>nww������`u(pdL��9#���QdM�ԛ& �\�$���9��=9WӘ[�7bƍ�)�ȝU���W}x\��ὰ�	���&0x
ʿ�����K���;h���T���[��m�K�e�X�r>y���~�r��9}�U>�+����]0�۫(��i�����S�A��xM����ײ�IZ���g���xu��B�!�Ф�Z��2�!��ѓ-|��E\�m���񧘞�����8/N�b5Ci��=���-��� �˙�p������2^��V��x"�C2�R󤄵K�΀��B�vྰ�vq&���	%IN*UL�W�tmE_�ɓ;�e�S�����RAdX){�D0��F��a'y3s�
񖤰Ѩ��ھ$��X����_<[U���x�֎� �q�����F�������A�Ȇv��:b���`D|H���/��1-���F��M��t������;˄���x�����c�L�APk����<���������㤼ߚ�n;�O���5Q&���Ξ$U��Kr�l�%��@��b�A�I��ڿ�QS'�Tu-	%�Eb�V*�/
��X��۷062Oo��8���A7��Mm�}�ir�z��S�-G�L38��P$�����S��qE��(�],J�!��✜w?��y&i9�NW�-���gXP2C6LKY>{��ʝ�1)�*,����%qI`n*�lʯs�����'x�QC��8��B��#J�nXu������ħr��:�e���e߻���`r:��[2fSz�M��D��>�� ������-��x�R�N�����hD�h|W$=9=չ=6BL���� �g���
N�v� �nfjIB|x�Y+3#�~i'�%}�C��{����j}d�	|��_���5�z�J�8Ʀf�-�����p�a���+��7�#UsK5c�ӲQ�˘��`#A��"��8�#l�<E�_!	,�A
&�r�?x���I��7�Z|�_}	ׯ�㣏�i�m�j���5Eu5��$[ݞa"g�$�t���2S�d_��7�5F'*��q�ϣ&�����u���%�?�0WrA�����*�W��F�)1�d��M�m�s�yl�o�mI���M|�h/��x��w0;;.�׶��N��tU����$�m�[nR�0��]���k�zb ���Ks��x03��0�~���$��g���>#�w��s�&���ܪa﬊x&���	H�b���t�֊8��m���S�,W������7��g���k�;�կ���l��"5d_
�c���k*�JU�j)_@Y^�%A�Gy�r��I[C��Q}��#	���F������J�8>w��"�(�����*��7dC����Bpo��$���9����xp��s�rB��d�����g.�ri�a9X{gN'^�bٴ�X�$���z����
���+�gun!_�Jۯ�qt�T��wv�Ȇ=��#�Hplw�p�ƴ��J�5	f�iܸ%�u2�q �*)���|q�[�~����>��%���0+�����F��/$�l"�ᑤ��3%���P������˦�Vg���^E�$@ǧ���1!瑕O:U���no]I�U�!��3tyW��]v�(�bv�;����ϸ�ZB!a���5˘���o�s��пK0�ۨ�VB�$��Ņ阤~`*��KX���c�|�����p_�ڙl#��/�[_�2��ϕA��ǅ2�KE���!;6-�P	�R�>^��a�ZI����^ ���(�.�{b֩�����I�r��z=�ɐK��z��3V^?���B$\:$�7.Ζ�*=�r69��h4���eK�U��p���	I�2�yĉ{���T���!�E��{:8�&+�8�v9�/6�0˗��$��a?�kW�}?��%��)��G	*T|�k�Rd�c"��Q��x`� �k欠�Ė�n����Y~;�uv)kQ�v���dc�$��X}�W����љǞ$'�+� ��2:�٠vO�
�����pYa	0�	��~�цFTJ,���X�9嬳���O�Pv(��������UZ���G����)=95V+u	�x�J����("3a�2	�KГg��X��Ʀ9,@M�����lC�����_��ګa��Y7S�	�s9j7�FTT�6#XTΙ�	��`�%0���GM�s�e�嬕�B.�r��+��KL�x�|bG�e%B��5�S6cJ8�����1I�굊ئ�*�w7��Ƚ$k�$,�t$�}�Y@��<��J_��A���G�s�u/����i=����(7:�]�ے���ŧ6q"�z��@\~�0C�M��K��¥Y@��8�s��,�g�p�L�\�X����>a��Q�_{�������`0L�L�n�%���P ]ź�Z�V��w
O5�U���V>��HPI�66ױ�r+��ʭ�B��}����+�i޿��?�ӎVO��7���6�a�1{G'�0��J`�A@��������r^�B�cey�%�P���G�b��9���,AI��b�k��7�=��Y�[²�a���3�*mR6�74:��Z�'3�;��eK�h,���EB���K>��C<��CIT,^ '�d��H�GAg��|�u���Jl�&_W}�I0�Iw�.��-��~����6lٿ��K��cL���<�Q�W%��HL�GI�+}*�s��3��܄�y��� ��A�"�W7��Q�����JI�G&Ӹ~#)g֒3�.�>6w�q�/%�&6Rɇ�9<�����?��������\�TQ����Vt��wr.ژ�K�Nk�:A6���$�������@�'k��[:�<�ĉ�W�y<�&�Og1�5�!���[xr�S�go޼)�<����CoF������W}0�!�-4�58�U*����0=>��zGGǈF"��2/q|/_ɝ��8�?�|~�� قa��)ۛa4J��Z��A6�E6��HB�E1'oSپ�r��;8�W
�i|�9����),]��zHJ΋Mg'��0%�+��p��\�S��w�^D�mc{�@�_��x���/6�H+Ҁ�0�԰� 10kJ�W�KVgV� j��:8�(�Z6��D2#AAR�m����'�S�����۠/t�!#樁"��7��X:?2N�$�[�O����I =�N�#����EK�:�M���ņݼ��<huENsY�
/�8�B�i��^�I~lf��UO��\��R�6��ߺ���vc�W�k�8�BAg�Z_�{qB�졭:n��|�v�w߸��5��/jX�=�KG|dRd� ��R��[{�L1�0��bg��.?˅����m�\!%���9���v�vo���$��%�cr�=��%�g��=9���d�9�<�� ���Ү�Wf=���n�$.��ܴ�')LZp1$�n����x��nI�T��|�A¿��������<G�\D<�RI\蜟a�yy�\(��Zf�SV�M��{�u��V�,㝷g��З`bG���g�p7pV��a�Ii"O �\�r��<|�Ý�S����{����p]��v���`Cۈ�}|]_��k�������?IF�x�jSa9��j6�����|Q���$-����k2�R��@Ul@�,��rG���/�^G4���.�D�WQ�W�z���:C�{����r��1.:��
�F#�`M�����������������������q�ψ��=�����5�Ih�U�\;����A��lр��5йV��B�)�Cc�����X����[��/6s(K�x,���$t'�Cr/Cbc�P�P���.&���ŌpP�[�Ǚ�%l@�$C�L��Swf�l"u�t���!)7�&������A��(^2*����<�`�0�9E�3���j�����r7��L
1��ch;� ���7�M����xp��]\_���&._H+��G����>_B��&Ff4��<��u:~��PB�KH�휭�C�B���s$V�m�8�O��q������S�ycS���J@��F����}I�rȗ����
�<���t�sVF�ב;0*�M'��`3Ӓ Xr��H�L)IA���A]�5�/3�Ԏ	~���F�o�C}~S�HXk����IyF큊43�MgF���x����f.���/��mzaNY���O�.�?��w`�WG4�?�od�K�`I��������0��T������k8��=�-k�����;ϥ�w�����3���<ٵ=*���&(~�A/�l�X�W��a�|��r� �0fF�X�����yW�MB�������:O�w�@(&qH8�:�k{U�u9'r�	4[�OZ��ܯ�ܝ�)�I�txV��Y�;��DbJ�Z�)v5��XV	E'�4�ha�,w��g��+3c,Ds�>�`�#8����p��aow_�7�ѩ	��̬_M�Ĭ��'�%��YG����53���v'!T	����YϬ��&�ft��?�@�a�A�DX���Z=#��&D���y�������V�4�8��c�"1�E9�El��HK$1>���X�aI�zO�Qe����ا��p��W�DTMc;	�V�h�E([F�c�N|ь�@�%���`Q��vF�����z��9�(y�i�\;��^Jȿ�8C�p;p�Yt�PNF��l=�k�կ}U��������'C��oN!U�q]g�5���"0R�N3�!L��!�@%p�Բc��^�Yn�ɂ󊽁#w5�\B���'$����*Ξ��G쵧��6}�l��^q�F5Kbnzq�;5Kɿ��*�����v㕵*�X�9D�-���}��c�%$�ηO��J���8)���7!�X|�Ǐ�u?Ȫ��䵃����	�B,��0���|}v����������P_>~���IP)�P���Qہh_�7��DP���U�[��*!�b�%�:?ñ+�2M�$���8}���H�JS��4��ޠW� ��p޹3��IJ'�$b{}Mu�j���J��,:�La�F[]{G�r��NO^��WC0��[�^ú;��B0�R*��T���_Y��ES���8�?ߓ����1���,8�A�egű*	��d���(L�+r��4�C�^1>cK��!�a�{`*���iv��|Y}��|����X6�]����'�9���H�����=�����6w��Ku`~	*�ݾj|�w�;R.Y���y� ��\�ޅ� .�-��Mn�.;E}�.��5d,
�L�m��h#I\sk�A<�)xI���V���:o��'qTh�DI1�O6��j�Ӓ&�P�C	���Ky��(�[�mɚ��
JULL-j��V�����&5����J&%��]���J��D���(�jE��ޞdO/-�0'�<_��m��2]鞚6��[p�[���1!�C����Q	\����䂋s�`�:5�3�b��899D�֐�B'�d�T�\�{HVd�UW��5��#��q无]b�Ij	��%���hx�hu��������Q5�W�%�Mal��>,N�'��G�������Ŷ"���}<Y/I� Aj��h|R��7����f~	����9�U����3�Z�(�E�m���$��yrE%�iS�O�`VͰ/h��;-��QOIBy�Z�3i'��+�H��*d������0vo��a@�{l`��AV�9������ $>�-���-�&�*^(�t�_�^H��ux.�4��8�!���i_1��P�	��8몼�IiSzN�� �]2([�>5�x����X(7�!����]�Őߜ�ĵ�iy�Y��$)�e�]���k��]x����I$%ɱHJ#��&�<QT��a�y�`�"]�
�3����P�w5���H�w���t����a�{��[��j��dQ�{
�f��"�6��(K J����������Y3��?%y�����6	�}��c+L��T��H�u������:��`q�������a���f���{�UZ�/���$@E���80�z��K�=����dб�FD�ޫ"�a�C��F]��؟bM��2>{�	�P��0?���YI#x{iAk>�?�`�@��fG|CԂ�Ζ$ ��"��Lw���~?�����ܙ$�R��1��t<%�)A�Md� @�%8$��%��N��dT�XhO���A��q� ��Z"vw�є3y"��$�dLlM�hf����}hҠ��~�_��;c
&�n�D _zwU��~�x]��#ٌ$��[��Q;�3T��M��K��kG5s����48�Oy�=	@)�CKۖ��������V�v�hg%��&�%��D|Qp� ��]�O&15��Ԥ$~�K���N�P����\g��m�E��$�#�$��$J�X\���>��!4����	�����~C�@�LΔ<Aey�X�Ϊ�/�zEA��CJ��l�,z���啟a!��3�R�/J8><�5�(\&��v��k���04~���#2�}�l�iٶ�l0)˦�x��l��/��-�h���1^n�I��{�	����(�A��pm�ۃ��3y0�,[�/�,#�M":�>(�_�!׵�3��G�l�N0%wzVmn��f1��p&~��#H��Q�;K���y$X�k�/�w��F6�w3B�3)kOv�p(*w����5��N*T6�2;or�9o���I=�}7���Z����Q|����pC���=�\����a�õ__�d�0Q]1%�s%[3$4��Xp&r�%�Ǹmai�����X��3Dmj��E�l"���S�sL�.;��xZ�C��#�z�K�|2���Ȓ�ע_�l��f#�RK'$�X��A�9�b�ϐ�ܠT�P��U��'�XʣX,ha�c+잟q��O��ʲ�8�/��!�sp\��B��rM� ,�$�>)���\����gL������ľ#��S�*c���<���?�����RJ荻�����ڪ/��&)�]�}�9�Ɛ��v�Z�$�o�ÄaK����O��ׄ3ʩ�(
�.~�o�v�)��U��Z��_U$`9��ő$0��I�F�#p�A��d䤍�&ٽҺ����">��-�gR.p-IC��,�]��QY6S��؈&����O�T��{���9�Uj�xr\M�f��.��ٙb�{:�D:���$����sE��f����c4+UX7n"#�
�sd�����έnC+p�C�b[W�2��@���3�
�$w�_~x�݉�<�;������F�A.�T3�?�aE�6l7Y���iw�Q�����;,����M-���zL C8 +����`��W:c�:��@}__Y��Uqv�Sz��"�Ϫ�p��7(��P$
�U�����=I(QK �Q���Ӓ�ڊ�FPY#9K��Zj�ޖK��>��Y���% j��0������s���>�t��%D�a;��^3��K�H��@�Q�g�#�?=�+޾�%a�P��r;���t�Ϸ�,�%�i�`!1L8(�����
����0���i���ɏ�*��H��!?)�"��>�7��]�����s�{�a���-��2dt4���Am?�?[�E>�x�Ƣ$�KKx��]	z�Cx&	���9΋MI �b(%��d>�W��rS����S�##S�Ur(?�P���	Tۖ����u��ŁB�����[J�ʪo�ޑ`5&�h�BY��&*�dZ��$����z[IGbay-9?��_��f��dsK�;��>��r�5.|�)����Og-'�w���3$��ʶm4߮ݘ���s3�OIx{N��Ӎ-	��D&�Љ]A���������E�ӣЏ���1�h����l{�V9[��Z�!���D�*
�����^nbR֮֐���-x�)�I�<:�3�d�����uZ	"**�N�J���o�9�Ox�~ѐ�͆&���e Ed7Q���td�:]�;����x��w�W�!�,�q'�\wH�y��`sw}M;�:��5�s&X1w�~�{���c���|�۝18���QY�B����㒤����K<�����$&FƐ�3���o�y[�2W��L��30�LD��	�ӝ�tϑ;���z�r{u�2.�S���˽�*�H���T�$-�1ɗ ��:>}�D�y?&'�ځ#ʂsHA&���%��i�jќ��+Rh�����ɝ���F�SL�ڲ�dÓ�C�����9.�U�Đ��h��������R�#H鞐ve�q���	�'&����+v5��y�Ʉ�������/~����8����YW�Ύ��<��,ҽ_|��~����I���7�tk���ы#��d���(�Ŏ�b��c�ֹ��w%��_/�����7�>y�������I)vf|r����~��C\��1Y�t�c�XY�����:�� �N_�;�h�� @������Y�XX5V)�NI&1�x\Y�	!e5�ov�H%� !��E�����DJg�) �"�50�H:���)�$�my�D�$���G�QY����H\C�����+wx���R�Hl�v^��'�ǆ�pv�`0�2�iL`F$�%���Α��Q7xzr�ݼ�	����B���7�� ��ʀI�9t~�L������b-����P�sC� 출�O�켅�l���/�P�!�hblngݐ����\׈�e�X�vSʊ����0�� o��ޜ����f��^-+��1���YP�a�����M�� ٖ�4�513d#!�-��HL��	%��D�������_��u�ԅ��z������?0���,�q��W2���B��ٓ��MA�����Inb�Q,7���U�UCrh
z��$t8O�X�+cr@�Slo� 4<&FR�o�f'�
g�.=���qI��gb�{$v�b��5�X]�m4��5�)ٹ�l��It9�����u"�4��G�x@�]���ߣ��h�pup_�.��at��ɛ^��zֶ#��Q&,�3a'qiQU76�����N�hD�⬓�?~��;���0������ϵ�)�g�g,�Y�Z�H����J��6��?5����M�J���"_�Ç;������t7＆;o,�ի�,���a�BK>J[��ŕB�P�KPӆW.D��U6V1<<2�Wq�lE3H��x�TE�e���`JE1����#�9�5��o�q�	�8D���xF�5���832��bS�5���+�9B�����ju���g����t�_rX]z{�<O�����A��I1Irl,,�"W�`w�T��	xL�����P�5n:}u,J�/�>0�@�G�=�1Uy(aYFjC��̀����yö
z6��M��z�$��cf!���F�Yc�(&��Zݨ����L�|9�q1L%Ij���5���!i��܈��{f���Ę&;d��ة����S�0J�	'%p"|5��C/��U`U���ls�s`9議Xq䣒���K���uu"љ-�8��+�C����
���Cz<n�긛����7��&�6�~��7�88�����'U1F���8*:��8� K%U�l�e@�n�n��9�v߈��)<O�/K���Q�h�^��ơ/���9*���R��I��2����<<�����@�+JS!��! ��lx�XL�e��A�o�c���RJ�tq~!	hP���FE�g��,b��K�$1��LƓ���rF|0�b�t���99��G����9���KP[�$�pQ�v�>�쓊np�e��R� �����eN���!���`ճ*A��x��� dUTH|`E��x�?��k'����P����u4�:���v�i7K����d�UV$y�x"��_v0��J-�]u~_�FS�YP	��`F=Wꭺ��8��q�Ŧպ~�^���J�Q)�%�����v�r~�D�r��r�Ii�!ϜҘ�X�����QS|�,�]O[�o|�7h��֠�OY��ay�`X<�ٵ`�B
����4��҄Qs:�VW�4쑵q���|���m߾$��8���(�"/�֤�V���^_�3r�<��yH&B}��ګM�H�����2�={� 3�9�E�"�t�L������n�]YCy�*�[�ucK�qZ�zK�?+�ɊlS)ڽL��&7Y�� �0���`؃����)�i<� �U����]H��K>�P��ڵkU�c���8JPGT��ŗA����2C6�UԊy���ԧP���F�kīv7�΃�6�M�!?��Q��#[�B$şt�`�o
T�3wbl��C	/�J�>+@�����z�'�ư�ʵt���4]=�I�></r&I8���������2��'�{/
��������̢�����)�)�b��@�X�W--&-p�p:$�#�q���,����3�����Nz!w����Y	ٓ���Ox�>P���gH�hs%-吝��'Sr��f�/�IEl"Q+^�sj�v��Kgj{:��Hz��$3L2H��%�����my>v,HB�qȫ��!`!*�#I�-�����M�� ��s�$�7Ư+�]����%��5Պ���$�y�*�Ės�^6�&1�H��,�����d����$�!����<f���o�ׅw��(s���w\@�����U�ŧ(%��a���a�·l�K�XT|�O�i2)qE:�ֈ�5�K��c�[�Yd��`R�J�td�i�Z�o2���K�5Z����"1��[#�FHr��ܙ�%���**�~��l�)�*!�nQ�v�.��-��qb?&���Q4�v$�8��;�%��:0�\t�{p�.�1�[�Qp(m�ό�P�.���RO�w���+�"1�w_�4ܸ{�(>>�N�1�S�ؗ�,d{]�m���vn]%p";5��,��Dh��C�d��K̔/��y������ز�c	dG��*�|�֢NH|���#"yXPc&wd:����*ֹ�.y$y�� @��G*:SO93�jڍ�H��,m����w	}UF���2�v[]�!1j��S����}n��vq����;},���� _/�ωE�Z��*���r�� O�077!vj{��8��m	�S�l庿n��`+k��10��[�$�|������Xڇ��(&g3� &���Y�O��@2��|X^������&|�T��1������1�)�K�C�7�U�F����!Ӛ&@���Akb')7�����O�A�%ˈ����F��q|x���R�4f��hv{=����?�=�j�-�cg]J8����T�T9q�W�7搎�3y�Z�)Nzo����bmOq�*2juԹZj�IG�f3���Ĭ��ߺ��%�A�,#T;P�z9�츉#QFA�E����>������'0'�9,����_;*n�KP"��������SaCŃ�7��+�4T��:K-v�$�������A�I���ju|�ð�΄ɒ�ϡ������LZW�\N�r��и���,��x�e9�l^�k2&*˜8U�ϯD���p1����H.l)�FftT�2cK�x���Ʈ��w>��g]���
go�CY��ɠ����8��}#�\ojP�n}&���Mi�
Z�v����J��d_de��3=1��b�h��@���a	�Y�����Uu
I9M#ƹ�p(�{&��|/�˩����ոR��Cf>j���mտS�Y7�B1Q�j��P_�L��ߢ���h$Z�	���&�8&����9�C8�e������ߖ`+췆U�q	J:m����km9;)����ر	���;��uxd]=����U ��T�=�yt��Vfxə��q�����|#���)u��,]_S}�p4�"�v�M�6%��+Kp/��@����(���L��n��lIN+-$�M/����=�]U$��rb��k�徳���Ā��c8��*�o,9�w��;!�;�,�>B��]#�Mt ��A�礡�����]�~�@��j�+!������Fu(��O|茭1u�Q !JW�+_���H�=�ZE�s"���^h���Ih��uPf&I��*��h��M����t�����Fvm�k�#y)�Ir�$3�FcX�;"�f6W6@~��<���:��m�$�7��ͮ�}d0
�zRG�_�s�Z��2��'*��9���Ղ��4[r������[�<~�\�M���$��Y�w*A�L窼���@��P�&]y�,�lȺ��AB-�n�ϙu��V�s:s�A���չ-n�١��b%w����,&���|�Jg_j�ި�J��ƩO��]���^�pa�
e�\7�?���:�'��{��
�M����.��1��}I����\��h2�a�1P�[�h2��ݬ����݋Gp�/ ��#DK��d�*$Ɂ�7�	+�uv���٩e}]���eOx�,����^�0�ِ�%�B����
�"k�Fh.m�jx:Za$:�F�M?��5��rF[ղ���C�t��v�Ѕ���zw]�O���Y�)����Ȅ��%�����toٍ�����u�o��e:��n4m�K0N���t�ݒ�p_1z�L��<�kW�����όc~��g콟$��+��^zo�{��w�0 )�RRH��"��F�R�� mȄv�\� �$� 㧧�}wuwy���޿��|����@ '*���*�w����Ι�5	�zR��-�aL|Yg�%�{��I��x�^��^S;���PUa�C���Ó��O��v(U��%i��ծ5$q��ůrP�g��ǝ[�����������j&~�4qXȋE5�V�&RBa�j�B�H�3�!k6���~�҂7�+;�ʓ��;�c�IB��F58g�݌[�ӢiM�����8�<J��r��8��q,�2񴯡���P8j��uO�C&�
�
�ѲY�1�?���P�Qe%�z��%Nt=��Y�qR�gd�*�N��@�~g��،V;�(.G%Gd�F���:%��-ę�(�i��vOg�h�<��a�Uu��V���s��9��(c}@ס��iOkrH��xZ�l+TS�3:6V9>���@������߿��#8	�\��V##�0��sDI��ʸ�&��FNH���x	3�*�Gi	3��Q��!�Q4%��A)̼��7����GpRꢲ�/�HH�#��(L��A�� �34;�e!�*�V�AI B��aC���ą���:"�ȨK�gI�v�tHX�$az�>
W)�C
%�&��
�U	J�%	�h�ĩ9�������t���lx:�<J�LO��P��΋�t��_~&������*./�����6|<|��T�ս2Zmv;�&��cN�~9}��Eۗe�SBK�B)KIf7����vF�J��5O�3� ��#N�t�+�t^0*�c[	b:�m%�3�nH�E_�B��� �{@(EZoWQ���hL���,&!��,�q3�`%�M��C�ؖ�
w�>u�#�q3:�ĉ��.a7���c"�و.�s��?����r�3�'ո��w�:B�(���h4$)������(���Zg�%ᗠtqi/��Pi�58	E����"Q�����C�Z��FZy���}�ô�L�Ƅ*��Z����0@�d��a��C�Ձ
�>zv$ơ��[��k��!��'N��N
���(T&"BFԐ�Eǣ��ьuN��n���'!&�����ׄ��)��,1:!�Zf��Ud�5�10�M�L�tZ	���$�)�t=p(6!�c^��j����Sq��J`�l;X�<����0�����[x�[�a��
>}�+�~�$!ay��ms�������t�B><5���q�=:��Xz�o)ayv�zsV!d,%�2)_Τ�D	�����YI�$�U��{1�(���0U�&1ԥ�%�y�"
�����_�S���r޸�th�¨ء��������g$�=D<�afjN�Xha����kL�
���!�c$y؅"�T�D|ֲ��C�L;�}eA6�wڗ��5W�3�5�kl�?ZO=���'%!�W+��_��r�ӿ{/,a{kG�z�K�Tˋ�]�:-��̨����cu�ᘪ�
Dǽ!��b��H��?{.��D?����9])�Z�Tx�<zǳF���&�`Տs��:���� �m�M$�`Hy�.+��s���[W��?��hX�k��د�'>+�n���L!'vZlT�����И)���M�0X��#J�S��E&d����YC�}s"����eQ��ZRMu�)��_C?<�A`p�&J��nMȜM���(�Z$�L��(������w�᝷�qc��kWpt">=ɀ'���z,IE9D�<�t�<�V�V��W����ɠk$��d#�
6�g����	��&��o_�BQlT���rO1��+�×�bks^�|W���W?��y,���n��!3G����Ĭg����k��=Jh)�h�T"�T4���e��A�ސd�0�I�L8��܎HB���X�78[�NOOӡ�|�&/ �dtC�(�;;'H�<� Ѧ-�V��nUMa�]�Ox�AOY�7_ma�E������ nom�Y�i�7�9�f_���pL��o������f���J�Sx��<-vstX�:7<��s8?���Q	m�����z��i�M���~ӓ�b'eO�[�*��<M�FSb6_�d	�[;;��7佚�P_;���.PƋ�lHb̴��y<���P�������?u�ƣ�ty� ��Hc��Ǣa��bێ��w!�P��%A��5;�|��-�s�!-0�����.��E,H�8���&G`$��񫭊=�&��mL��/<������<�ɟ܋���K��� ��!ո:�IJ�>>��ʘ$����Mx�>Vb��Ҟ��Y�F�GN�l�<FB�6���ޣ�Ǩ���	O�n��#s�I%tľ�@kBL�F揦3n:�s�>�9�5|?��ڂ�Bƌ$�<��3~{������u;���ZpvI�ǔۃh�tQ)h���(�M$��C��`�!���8O�z9O�Lx����J��H����e!�8�Db�=4]�L��Y4�aH��w,]q��� q��~K7��1��B�|*9�k��^���<Oj���޼�d%~ܳ�bq��=�)7j(��X��r�c���5b�}����c�ƿ�
�Ι.u���q/5�!ubE���r��F[ŀOH�<A�S[r��������sx�v�P6B|�^�$�9A:�[�W�HL(,�7�?�T��#S�L}�%Jp�qQ���c,ٔg��		�}4�B��t��<'��+4�k�]>V���W�j���x�b��H��&!?O�K��{6)�f�e�@[~V�_"����vZ�'T6�=j0��~���3J���Qa5<\�d^�e��Y����O�g�֙ʋcZ�JpAv9B���3�gPo�pauo��w��q��/�z�:&fǴ��if�Td~���>G@c?wd0�����|+�10YK:��8�B:%��AJ�0��Y�:���Ɏ\�A�:���fXI�M��ٹ0�; 7�4�N]�#g!Du�r6����$*������w����Lv\~>&� ��Da���f�����7sY&�$��� Ͱ�1���mJ�DX�g+Z_��Z<�<�зue��.�2a��~�g��ӧk�|u�v�p� ۛ��zc�|���Vg1�xs�º����7��\q�^��#du�l�ˮ?�&�.m�p��=z�daLgQX�1��3�A���ʀ�*b��3��簲pY���j3�%�.��H�M���Q�^�O��R+��o_��s��t5G���8<*cv�Í�9I�����qL]OI�'�~��B���_����F�dK���~�6�1fna�'5�4�����R��;%=�C� ���JX{��u��O?ݔĵ�����tq7�M�\�Ɩ�'/v����Rk[}<gDCa��C�� [0s�F-�?d����T��(+�X���O���1%�%�*�Ju�G�"���EI���t�g��M�P�����$����r����d�L�D�����������່ȵs�TE|�y����buqI��>��!:�8���dY���3M�m���(�9�v�	�GI�� (d�B�׈���$�e���g�J�J��o���!�]���-��O^bkW$�'�B6����O�����u�OE��v:��HO��i$�(u�� `�>�<�P?W�j�9$��Х3i��k��Ei���}$�c�ů���&�GhT*XY�ӹMfG]� r)fe�u��6%�x~n^	��ռڹ��ee�,$171'v���K���ygZ|�/If�ON�I�NK�gpa�2=�*�����͇�XmoOJ�m�H,���d���k��|�f�H�������l�ς����fV�g2){����K|8,����7�Z��k��]�D�q|�����C�h��-j�s�;B��m$ߠ��`˂�@�F�3~d�����2|��$%Һv.d�6�e\��@��Ό�Kf��_�:�l6�sm=��1��4Ҝ�����e	/��d�q�5~CZ\g��%�,'吧�ҨV��Ww�}��Cb��g۶��,�E%Өm+�5&ke���"�h��4�^����y\g�91�YR.ϒ��ܲh�����d<��O�gO|,��0�U)�G�9D���gO���,#��W����,�J�?�G�h'۔��m�_k�������N�9�c�l�B�w�He�b�(n�g%4��Zv)Sf��\Z�~fwd*m1�h75����p�A󤫰b���"�'I�K��`���l~H�)�\g��d�T�Z�"�x��e2��w&���$�LG���-i�L���@�Cq��qT���)���%�/$��6��ԑJ�])��Ǿ�Z�p8�Ԓ��Ӥ$�t(:�1)��A{:Π��'`O)�	O`��)�ZG1���#����L7lO�l�dL魫mBAC�F'^��ݐ\�.d�d�1�4&����	:��h�T�Æu��{-S��b�]'�HP�/Fwo�xe2h&���(�K!U*�`���wG�M&�#ঁ�ڤ��Iv��;<:ƕ�Eܹskk�4��t<qpk�y盘�A�f��{Z��P,�h2P��Ǫ�����>��Y��U�7�kt��Y"^95�$����W0U� iw���ˈ_���7*q.*�^�숡lJ "�#�ʠS��0b;<3�������^�Y���=�5]{VhX��L����8������p���k7	�z��ϲg(�;ji;���0}�\��q06.ɠ�V4��z�ҽ�:���XY{5p����r+D�[��}c?��w���
��*r�Jg��ıwP7�˖��L�1��I�EH�&AP���̞✡��]'΅r�!����N����x��$ؤة�(��ݨ��i����5�_�+�{�T���N���~Q��]��L��ͭ`jz�G��>4�>�Ґ30��GO�阇o���g���iG�P;2X��"��agT-��	��y.�j9R�@%���t
����Ɛ��hH;�쀄�Zb��wv7���ğ���^�ǳ��hJ�B��sWe��t>L�1?�UIU����U��(1{��k��A;�R�H#���4�D���z>\G��Dnl
'�$�W*G����g�(RgSh"!�[qs�9\��#��, ����8��cIpSH%�F�����BE�A/k��+K�8	���ϱ�����#-�%��m*�-qt.�Re����,��>�;Vj%q� 4g�2�b$�q�Q'�H~�"����3^|����T���t1%A����x~���X�����$���q���/�_�Y$�k�2�#hܩ��K�#&�¹�8gH���Le�'{���!�,�t��Fs��;��~�2K&3�G��'ϯ%N:.>t<�GQ�e�UE]�Y:�s\�8��iI�d�5N|�>�!��F����^
k*X<н@��\.�)I��ž$q�8��"˝���*���B�VO��#�9O*�S�.�_&�C��p�0L>�$S1�|�vT���d��%#�ǱE�Ӏ�'����Ľs�Λ�\�����{Wu�2�q���,4ddMb���[�m���x742O�I��˨�ng�:D�zr]�>%��g�b^_�*��4% �TƇ����4Z������KI0�`�66/'��M(l/W���y\�䨶2mV���|L��$cZ�൤gvaz�V9�6T�I;Z*uTs4%6���#Ŏ�&�Vk0��uf���ݒ�]��:-r
�%�q4Ab��sa�5\;�� �2�2go�R3竄�LS��ša�e����lm[�d��i9�crn2�)�xS|Ʀ�')-��P��tm��v�g��$@���U��zѮ�}�>�	ZJ�E�J�m�J���]��I������ϕ��A��%������qP�s�s�F_c�!���r��.�m����0���&�=���b;�����PDΒ_�����VH��ds�4��[��N[�od�LK�����]���}j�1J��xř� B��g���%:<<���֟�^�$�N'�,�:T>.I�<�q�k;�A1۳��AqA2x��M���+c���i[��CrJ�8v�AB�;wQ:���}.����*�5IZ����7�E�ِgC6�Dq"�k�=��ߡ,�DQ~_���q��H.Q�����ʘ�W}%�!?J2���j''ql�:o��lP��#	U\��D����M�_�̒ȁ9K���(�R���}��+H���:��N߷g!�L:��=��hh�7��ceeA�N��U|��FW��[��?�
kԦU�|LD��l?� _��Λ����ЋSɰk͎a����p�m���Շ/4���]1H�cD�dW�͓C�4�4�*�s/��pXmيEG��݆Iq��ͦ�8�����>6�rx��'q	�`S�0�RJ�B���84�����a.Ȅ��5��i�F�K|J�~���⏜J�Tr6�4%zѿ�����P�����z��Vo�߿��Ws�ۭ�t\WXk!U����Y��(\20ԧIf����:>��T#�!xP��wY��	:v��y�?7�Ӑ��@�Y\�o�O9���ꄝ���UMNPЙsJ����lh9y1�䠟���իӸz>��|��@��Z����.,�#73S�j��ܸ�E7�Sx�ӧ���I�E�D̒h��4M�=�&�v>��VםwF!TB6I���_߱]\�Y���H��	D�t��U��.�f��w b~� ����\�ÅK�P>�4��/��A�=R�(<�EC���: &�`�zԮ�d��^�� �q�Ae�9,/Jp������ĸϮ��>�O}M�	q	����"/�}���uLI��FK����.\���tR�!v�j:ϳ47����l���W6�-�-`{���Ba~��#���
��6��ku��YQ��i��[=N�`�.0��"�9U��1���3���5��i��53�j��d���n?���3x�/��?��:�c>i�?��D9�~:�L|<��T��~]��{KWP#3�S
u!��c��=;�u��ew�痨ʥ�%L�Ϣ1kН��!�DBe�K���?��>)�˰��ǟ<�G��b��Eh؀;�:4�[-2�����}��������cRF�#��B��V��chB&�DQlP��d�ͣ[{,~ .��V��f���ڜ�Pd���zDT�Ɲ�'e�Rb8�gB������W�����$ڑ�7=��~p�K�xx�S-p|�ɧ�7>@J����gP��� j�f���(g�I_��#�a;5sh��h%Lm*���Dn���0�&�h"=�D��V�)XU����E,/�P�s�oyZ�x��'�����W��	&H��<�4���e�ٱ���>���&����gC��d�><b�4����U�+@鸌�Ĕ�{J�A�Za�(�I����0*����(#�����+?^�b�
t�-����e���S�h��w��:5�p��UmVI_��o���~g
/�ʽ����5�g��Y�$I�*^�%ƈ ���51�{3a1�OSr�8��ãn��{���$����(��7g�h����L������ƵC�D��7!�gT���\�	��k�8�$�B����,�kM�GO�
\�H☠����;h��贎�.��L����I�n��<�ݐ�ф��N�X���[�]+���0$Dv��W�@�����U�PP��P�xBü|������h|���|�9�dQ%�g����>�rN�ak/��ѓ��11q����+��OE�D��0`ar�hA}<�H˿���:@f�����g`L_ܖ8�$	�;0���5W��D���{�tV��ydrae�e�з\_|��F�$��[r�?��*	y<��'�ŚJ��@���!g��	{A8���M��L��ea�on�!�s���,=l\xf2"��aLC��l*�G;+	,�T�?4��4-��N�+欚��=RI}ΠF$a�,lB�$����zu�Z�Pb����5��'&1>1.���;X��&��)B�m�Zh1���1��!{Dv��wS�9�����yԁ".8���S�_=��_3�	bK��*�f��q�5;=Y�r�4n^��"<g�#�����3���#9KU.?�K��P�ɡ���v�[�#;D`��������d[�̙���b�A�y�eϦ�������2YEט��G��Y������b�kJ�4>O��|H֤R9��9�X,-	pVd���=�(}E�P6gM$b�Y�}U�eY$���%�����!M���25���%��K2�I��F&$�ɦ�G�v$��K��1��C����6pP.���p��%�b=�/3�����tZ�d������������#�*�� �ݫ�i��������*t�7b���i-�3�X,?�3sGɉ:5��)�a�"enV�㝽���v���.����X�+a�n{b��~�\�A����N��h��gѳ�x~���{A�t'-L�qFUp�1	'�e.���Ow��/�O�'V��e�07�1�5DyL-&�SﵑΤp��<��K#6$�&��vuq�]Y�ى"޾u?=�X!��tT�s�'��_��So���?!Ni?]��g�~��X% �R�<M=\�oŁM��0����zn��p�
f�y%|9��sIg��qZe=gs�a=�:0{E�(M0+d3��7�+��'T���+�wk�P֖�uA٪�**_��o��Z)tmB�B3�ף�8eu&��!
A��=x�!��ь5����|�
�d?��J /��k�,\\�x�{;��C|=�8﵋�t	t"�e����;�L�pqA���	I��љ�Z�,�e ?/�]�e84D�^F6Mm��K� &@ԁq���Iq��K��@ai��a�hqI���8�9s:�1#�;0{����/&�3w�����011����(�C(�T���+	��4@�z=9�	y��.�;hS��~��Ӗui#�C�X�3�C{h����_���`o�<�Ǔ�qq�ַѮ�iI����޺u]X��1 ySN��IY����12�v�	I�2��\q�6�ٯ!6�SM* ح^ZY��T��
�;<>��W�hV�
��a���V�B[ZͲ˼t&���1-L����K�eMf3��@T�AC� �vtȚ;Zѯ�Kߞ��� {�]=�Ɔ}3{��M�;��|n^썃��[��=D�9��2�����'Z�fa�3@$%�����?
�����V���ɮ+ġ��%{���8��b�b!��}�Uś7�η�������Q����8�8%IMݶ��6}�_��M�Q,��@A��X^�\�~/7��Y?Fnlcc�hWk8�Wğ��ʅ9�%aW�[��'(�����-���'Q�DD����		�{ht��s<b�,5w	�
��A�(�����w��rϞv�<���M��<?�n��i3�vvGW�P�U^��}I�(G�F1>>���Օ�jnHP6�2/�'���+>������Oaq��k53��ѵ�3��4��p�=�Y���d�����l*gy��ۑ5i ��y�L>Mv����q�����c�:lI���3���	j�cI�)�N�;�nP"�K.H�ۗ8��>���}���&#���֌�@B��DHEe�'ǵ�FS���$U�HE��haX�Y�d<�PMl`Nwv2@�NOK�U��g��G�gfϔ��k����j�6�ǡ!�т
;�rsa����e�;x��j|X.��`��c��E8Q�I�q�PcF��.-m��ž��?�G���dG��z�wy��|�Oq\����k+X_��Pւ,��T
����q_;�v[������ʴ��ژ��`<� �!�k�K�%1:��y]��p	;41->oElP.g�ԙ�����մ�V) 5���5�亰�~�̖y�Mk��Cf��U�'ɇ�ȯ��*P�wʀ|F���sz-B�zMڶP(�I&I¸�dr?7�F2��ye?=<��R�$ljZlS��J��rgٹV��l׌�p�����s�V@Ȱ�:&�bh#aV�S�D.�I�Q��$΢Ga�H]t$�����Q��2�r_u;�'�����jt�o��Jjd�'
��ZK�I��gq3���>	-�l�<�z��P�z�F�V>�B2�V*UEwQ��(2��D� ��3����������́ekf\e�����bW=�xBɾ]l�|i���՘M��#3����Y�9G`h;\���Io@<*M�$�F���K��d*#0d QN�F��hL�!���NL�ӄ���)\\�P'���,���L��~5��r�;�$��censQ%%Q�L��v����S1�V��os Z@�m�{�}�|L��P'
c1 ef�{);j[+�dԙ��сZ�97��I-ԍ��Ŋˠg�C@ꥮih����8qx!��_����<z���)�0��q}����CyϤV�0�f��`�A#;�A��A���:���m5t�6���9���7l_d��9�]EP�v��ы�ё@�+�ۨ`q"&AgVߓ:7���$8}�E�=jç�fw��|Tn�<��rVX�.�'	�4����v�ʎơ�n���\ǉ����i�M��V�5q|!�&��Wj
%����}��������Q)�@r�(5%����P�H�/%2g�\:i[gõ���&�&�е�����+�$kX�u$cӳ'1C|��@|<"�#��D��=6pU�Y�7��A�lʯ{E;�03C�5-��Vg��^k�Б�k���=:ޓ�S���ýfO�4���;�I�U���{�D��jU��IJP���}�)\DU���g}kG�ꮬOY�eK~K�nA�®�{��$�qeP�WOP�gAppx�k�!2��V�,ۖ����B-����I����?�㵫��z8�
���4�wmw~�D��0����J�=K�>6>�wo���y��	=���^%X��,]����5��NZ��
��o�ؔ��.FS.\��)J�)�}�8J����y�V'Q�Ã�^n����}�vwem��Sbb�@�c��=�}����������pu��/d�4-v�1l�Ӯ���2�J ������/����լ�U���.�����q��ck����x\��������)���(3#2��i,H��C�$h�VG����ًL�}�l���g�5�RZVX%�9�F����RSls�O���hؽX���}����$�Ib���s9I��} ?|��s�{!�O�S����gf��w
,��uDWv4�tm<�=K'��uZlq>�Ck/噝�����%�;�ʇ�V7)	����
�$:.>��$�sXI-H�I�qiyQ�I\�ഐ#�tvo{���O7Qi$�$�^W�\������˵�B��=��g��k$Biy�!�V�&g$�ʉi���W���! �\��:�����@q��BI���Φ���T(�@,Y�2�����aqt�|v�s��CZj��͎�i|��]l<����y�v�*����8w9�v��#��jҶz�3�+�Ϡ����cab��oGS���XTZ����z��
"bQ�XzI<�*rz�x!�~�;b�qp\�309^�T�"n�*"�w�_<�.OL���
#[�?��bR����=8C	�=l���j�g)����\��'(����ծIl��e��l���*�΀E/���Y9_�{�O�.m�6�A�{d�VM��v|�@��}H5�C&a�TP4��BgfϘ`��Ϭ���̹�D� �F�H���@���D0�[0^`�%�����NZ|���!}�9����[���1ڗq�A@l���?!%����F��e���Զq��n\Zƍ[�r����E��SB���.Ju�o�YMn�������0�����۬��A�4Ǳ8�W/��ujʒ��
.��kRUo���/όcv���O�4F6�P���a\|�Rt�����r� �MǛ�1$Q$�3Y�Y(�����ĸ�5�X�{DG��汃B��"j�/�����g��h!�%��?��A;�{��,`V���c�=$2	�0:6q�%��{�a~������ʺ
q���1�RFYV�"J�5�����>��թ�"f��TF�ٖ���]|�dqBr�q��8N�L�$��$�5�m�H8UGJ~?-�<a��L��Z�C�)D�Y#Ԩj�)l���R
�5T��D���f�v`�-�kt-��c;�����,�4��E�R���C�����0�`��nM�÷c%���3���O*T�g���;bD�M0�'Z�����=�3Zr�9/���p�GU2-��˱~5�f����u�/g
$��Iy�IqD�ŕC$��Z-�4�}p�VIn��=��f�}oO��^[��S�OZb��ٍ�d��1�
il$��O�����MfX�#旉L�^�Y�a8�s<\&ʼ>�;4]@��zd�#6Y1�a[a&�N+)�!�^�|V�(���}D��� �����o4F\�]3��f��Ϡ�m5j����7Q�\{��_��AM���qE!��FWY�ڍ���>7�ѻ!���d96<���A�M��(.5mH*A!ֈc�;F�x��@�������.b��XQU!�c�cXY���TO�U�h�{�1R<�'w���5��-�[�NJ�Ѡ�ɫ��d��Ȏ��Zǳ���ȳ-R�^>��a�xy6��6���rO���W?���RŴ$:r�=�;��Z��1�����&n�'A)����
%�!��̜yJ��J�ca���L;^D�JǏ��Mp yY�7R��}q�dQLK ��o�bY���+J�R�$C�rߒMa︁���I������� �U}�v�˘94�Bj�d���t@�t��,�h	3��{�I�7����#��d�$<n�ϔ&��<f&�{���Ouf%��������7;�E%�aw��
����#��@�0�ơԬ����f R�H�f�Hl:�6b��Bj��&�c��gt޷�m��'��S?l{�?��z=�k��	9{ٱ	'f��v-�և�M7ό�&�0]������bX�ϻ}�o)I����c��4�}�l�T�m �x�Fw���e<Y��M�nNЙ`���ϢK1u-����v�4����pH\�7�Pf+#2٘��Y��c���|���ҟ��!��˸su�/Ŷ�Ky����|�Oo��u���8�_Ǹ}�"޾�{[8|QS���lؙ�W�ru
�����&����7n�����>E���ʽ,����o�A������r!	Pg����d,)gr�aG��V��J��Q�i�L~�b�3��LR�����ae,��%��y]"��Nƹv۬�!G0P=��_'t��֞�gɠ�����8��$�5L%0�`"#A����Z��O�E���{"{�����5( ��_��<�5's }a��V@�cIp9�Օ{n��$���J�K�֫H�,N��?����/���dӊx�q���v�����<})	?G�"q�b�r)���ݐ���2�7=���b"�ޛ���_����+\�q��_\@�8����op\:P�]���/(�̟����FL�
B��bk#rf�f
b'�ؗ�$$�!�}�jfvtJ�E��<�����s�z
C򕅚Ɏ��@xz�L2-�"S��b�V��xRO�Ǹ�Q	P�'<�����뫗����[XZ���n�C�W6��W��? �/M���0�*���0!��N0���gB� T��>&���K�S�+�?0B3����5�3w�/����.�$��N���[!=ߍn?��=<�-�n�0Ԋ=�y���̉9w$@�j��Bu������̎���/�V�q��ܸ9+�C�~$I��e���[��������#�C}�#��� �3�CBR�F�}��<%�f(�N_Q]dO%�(h�)�TA`�A�X�[/����T8������x�r+�Hj�)rƵڬ_~�/�=l�|�T",1��r~q1l��}T�M�Y�a2H�c�;ԙ;��ظʵ�8�S@�$�pSZ���ސ�Wg��a��Dg�6Nd�6qqic�;�T���{�-	�a�'h��E�qx���b���)����4�gW�'{iZ�	��s<��!�ϝǭ�bGK=|���Q:>�sۖ3u��u�~����_<SQ�^ˑ��".?3��Xڋ���*>��7�#
n�_�Nk��T�����*��|�#)���i�[Fv�r-\ېgyJ���ϟ��l���t�r�2�����l\b�0j���k&���"��Pԇ�X�{�լ���-��K�d���Aw�uOd?P��!��+�{�2oސXK�v�٤��
�[( �K�అ�RIc4���=8���D|�d9��Ċuėvڞ�35��krnZ>_���������5g`bG�G���\�ϓ������r�:U_Qffo�.1	aD���CrV*Bv}��cc��2��"��49�f�A�Z�a�?���	��)��E�0���o�ndo��	$��Om��[������|��n�*?����g���ۉCs�I�����s{;�k��+��\�k�%�,���+:�ɅeU=I�l�Wϟb�WC��A�BJ�� ����"��$�"�NS�g�6J8�� FL6!3{һ��(��S���nӰ#�A�W�Gb��M+\�
sH�'�)�ޟV�9�)�,&.�=b�Y���d���Lv�le�4�NA�*v�� @�Q��@�x�X�7���'p �`��X����Y1��X|rW��ɉ<��h���t��T T3�7ݫ��g3|�RCs�ܠ�mi�U�A���VY�%kr� �� �;1LLOJ��@s^��2N�_���ja��+����U�z�吓�v�����4���Z���\�Ĳ�W�G6�L1����JjB!�xfL��~�H]p6�2=�30#Tϳ6D=���^W��x1�+p�����Ȟgh�N�~�%gf.��}Ԇ�,��]<v���GK67v;�[[��D��/g{�Ƌ
�t���r&��Z�#�.vB
o�.�㎠nl��M��F�l���������r�y�M<��P���&&��nv�ҪB�6^m+�'6x{7<����0/מO�̨��=��<.7Q��K�U�`jrF��e,�gEc�=I��I���<~�������BZ!'���䤒���eM�xFYEV�2�qV�O����&�Ƅ$-�䋤4$���m 0��5�����M�`�b����D��G�r-�S�U��V����x��F+ˋ������ؕsm<[?ֹ BEI�O� �bʐ�44;grdH��~Hưu�X�i���--��:�-Ϛ?S%q�$�x�d���0� AZ��b�Ku�U�SH"���=֡>a!�b.���>~��_�`cC����f/�����ے��]�5LQ~�ՐD�3�:�F�y+��ﴍ�.�'�3��}�{�2��������j42�ʽ�ņsf�v�K��n��_�N��aHg'�6y?ո^Zı� ��4�7,њ�Iම8�;��cQ���DL�����M���O���:J'C̯ܖ"�Fh�|�ԸW�0����a�
i�T�ϒb�U�j�:�}�@�W��M� IXe����L���	!��_�Hp��"��U�5G���
����5Y������S([ȍ�~��w����0U��3	�8+9�u��QI��_�@��W$��ܼ$n��'�䨲�r��'>�ԐL%�(�ͪ���"<�v�L��"ş-�����l��)��HG�����LZ��8@�6�Sx�� ��˷5KW|��*����������Nư���ݯ>�{|��Z2���v��h8)kѵ#�$�C��2W��4[��W�Jy��Q1� �GJ�5��$y}��^/w�
;9Ncy!�tV�j�}�H����N��~Kmt����Kc�;|���#���W�O�����W'��"��RKݎ����GO��{��<E$Y� ����W�arf��%����n��DN�j	G�N��G;���k���%.#qF&��VȦ�Az���b�A4�l�0,��6V?~p�=�+�8�*b��-S ��/#���
�͊�J2��w7����"d�zzE҄-���B~p5A�c:�f�_,�F51�1 W�ȡj��%��K����{���ή�$+�T�Cޗ�/�e?�S�|�eog�ؗ >�Ob2�A�L�M9c���d�����/�S=�}J��D���D�Xo��7��e\�>�N��>C2�G���P{z�;3Tx�o�e�0��].ʳ��Yh��{d�+��f�C�c���I-Ù5�� ���SG�*���\���5߾�*v&.qDF�'���]��P���e�ymNN�P�*�ױ�߰A��V'ó#@0��e��3�c�r�|�~_>���	��=76��TH��6�C>^���S�_�'�Gd��������I�9D�t,�����Nk>;���*�����*Qt�¼ܼ��'O$��$�unJ�z�¢v�w��H�~���ϐEM�*�D�k_�u�ɺ|$�J��Pt����4��rb�Q-�7�hߪ����H}�hlcG1XXg���f�Cy�Ⱥ<�VQ;9T����U�+�h5{�ٮ('@(96B�����D��2U��� ���JCt�|�������� �,�V�b�f��P ;פ�#	�X.-��*.-�aJH�(�CU��f��ul�K��#� ����[7p�ܔ$q%Z���?j���	�m���n��(*/�U���V۲�(��i�*Q��<+�$� ~�Ud�RbׂǰvT�Ϊ��2OqFFj��d"`L��`�B�}�����l�0ƋYܺu7n_����Ka|��nVc;��ŀ��u�۪�v
g�W_��W���~�ׯ�>C�͋�(�����h�=�$XJ�H$\	v���:���U�_�uW�7.-����ɶ܋lpq\y��\wn��5j����Fm᭷n�{߾�^� /�G�3е�1�rE�	��ڡ��f[�Ž��`؁q��������Tq	���¥"�ݘ2�0�Ҫ+,��n�-��<� �b�����
{Sy	i1�/Q���<�J��M٫$�Y����$������c�����U�Ji��H��hr-�t��Ӵ^a�H�&p�A"�1�Db�/���������Ҽ��=M�C��4�����=۔�YԮT�Q�����[�5�Mzh��<p:�ǵ�8>��>�l]�^�|��~}Q~��W�֔�ig�W.a~aI;����!vJ���Б�प:��l���R��S`.;4�h+9O�W�I2��=�.sTg]��Y�0J���c��
6S�3
��0,eD�M�|nI������z�%����`���7-WZ�R��h��L���0,�c!33����HX)s淍$�K���+9Պ�ka��\F�+b#�{5�+�mJ�6�NnN2�� �DXa5$b�K���u�wߘ���W��,]IZ��܌�O�W_<�Y�O`�����p[������
�ay���c|�B��ؘ"N\I�X����f���YXj�pLϏ+,�!�<�O�([C���؉P<d�}f��84
G,���·۞����{_���۞�PA�x-d�	��$o�U2c{k�'������2.\��7޾���ʪ�I�ԏ��u="�Gs�C?Ш���9|�ҧ��g�ɹv�TL׈/v��Ēb��/��5���Ld��*�s6�Ą$�3���A�e�j�����x��w%�7��7�[�_�V��r��d�ڊ}���*�\.`r��gbg�X`HGpT	�Wߗ�'���Dv�<O�Ў��8�,a�9Y���Gm-���g�����yv��7I��D+`�<QBޙ8������E��{ct^=	�|vf{�P�)���d	j`ց\!���I��m\*L�O��~��5�ݸ�)%q����$f��7h+����E����B�2X�ԅE*v:�n��P."�7qX:���>��zŒh��b�~_|S8�p2�h�v�S�mO�𨎋K9-��:%�z��?69����$�<{I%<�-5P�����,�]V���6s�uivZ~���ڂ��9Pڜݍc��M�E�ȍ�5�6���8L�#ʶN�:v����]c��Q��m=�a����^ɳ��vH�X���0�|L�U_�7<�ѕ�-�~�Δ>_�jcs_�{�W[�:f�.L#�ɉ�0�
bHP�N&����^��;˳��CkLLId87�KR������P�%㲶ء��rFHhkLxtx��C��Ļ�~ClB[�L��G��������ݗX��r��5�3}E�p�����}<}���3���s��Ay.�5_S:6�LI�%v����k�CQ�b[\~��Feu£�\�)6 4�5�"��k	�8�i�j���O(3�P�OI�=NMp��$aS$)��8*����)6!�dvn��]tlvg��G��m8-��
R���f<˽1��R! 1��$�ia&�\6�NZ��VW�������Q!���Ϊ'�)R"/6nwsϾ�}I�(o�����7����I����n7#�r���ה=�	9m���*��Rq��.Z=ϰ�;�&}�oC{.Y<!���P�\+�NOO�Z�M�	�|>�l"h:�#�ekG24`a�.[��4�EG��=�����dRa,/�G�XD<3�ra�4%Al�Vn��j�k�2���|�Q2H�Hl��Tq�,FE����'�C�͘Å�I��D�Q!s+�O��dɡO�1$Ý���o��9Y�#|Ԑ�p���KX����=ս��/�ƭX���֫x�hM��b�����KZ���$OєV�xq���a*lf�T��t�tfi�ٹ��&�,
�)�I"L�Hf�4f���<���2t��vХ�3<,���*����V�r�z��{�����%e�b28>.�&�S=������1��1j�N�V��:�΍1J��Y���r�Ӫ�%H��ڙ��$-H�DA3�I$�Lg�`�@vk����jm/��$����~�0�ba!����?*8N�tB%���ÿ�sL̍���'ʠ���Ž���ѯ~)����C�Z���Lb��e�/Zߨ(��%�@�1���E#L�S�Lv�l�!tH�S"���x$�]�v���<�%j1�?�"�fOx�����g% x(�����U��o}�mL�Jx���W/���匐d"����%�8#�EO�8:Hƌ��-�YAf�И5�9�T> �^��>x�R����*��!5��VIa��;]��HN�CS~/9�z�����|�R�~����N�AY#,I������ߺ��7q\>Q���I���_J��k��(��x������_1��G�Q���f�A��!��:95��1�0sb�rΒ���>i��<����5[�����3�*A�q��c�4�M��+),�i_�!?n����"����X]�C1�������=ܕ�Jf��0*�cJ�9�VK�N@	M8S�:�f`W$����#v��,��]X�o%Y�N���QΖ6�`L��K7nbn��|:��(��W{�x�q���.B���}��'��Wq��V��5$ّ��t\�����dC�/��$:'{��㏰�<-�w�,kG�\�b��/_�"��ajvI��J��Մ�]8*c�Q��Ǖ��<�f�l���$¸Y��9Ǌ���{
�?�3R9A���?M+L��|����F�Lv%�}��9����'�(�r��x��<^{�k�/I����_��ṡ�+Y��7m�=�eE��so�*{@�zrn�yQƻHDE��3a���pƥWG�.�\/e���{��G�	<���J/_l�_{"�ƛZ��s{��������w�s��\T}O>�z���A���k�%d%8U&��g�\���"�$eW��k��.6v*X��'���@!�ԅ$t��Ak�C*S�R<��;-IBW�?yB,��HdF�S�XE�)R��&#��<C��au�]���gՊ�}�g����?�g9
�XZX@R����$J)��$���/qrR����@����wg���{�m�3���"G�m����q�l��&C�JR�料2g�bW$��B�j7�DxVڻ��=�J'P9��çk��/���x��M��rf_�@�#���N(e�ĳ�]�ŏ^87�[7/�d�ۼ�r=���P�3�guvI��u�D�T�Z�vZ����I8r�q���>g���D��| !���uU���uF8c�� y��3��n��%�|�+(�$�PΤX����igkl,+Ϫ��I��f$P%��A��{����ȵR��0P+$6����	F+����Թ:>�j�خU���07�����v��9Z ������x��/�qR�H"T@$-�m_>蠽��d>n!�윉kU�Wn(�-���B�{�ņ��=�M)U��b���'��	�ԩ�p�6��W��$����B$��IK�KO�I�j����΅�$�O�.I�;�ۮU��M<���1�J�p? ���Ԧ��:��+��ѣ�(Wv��ONpl� �H�7�l[y!��#��l���p�f��̀j|6�'!�/�^�$0��㹻w����y�I.���m�7"o��KR��5���ֶ�2ARl3�Z��&��R�&�hm0IrT��^Y�l���;��z�d̗Ȍ�Zsf��C�Q�p����e�>C�鐳y�8!�%��{fvPGx���خ�E��v|�ѳ�yB��.8�@s�CaqƁ"
�p�ڌ���GJ=���awkO�Д��b'�ο�?8p^��&��GY+/vgG6A���7�lTGu\l�5$�8G"A]/���^������iT�K�����b�Cb8�J%|�o�O~�VW�%x��p��4^<,������l�پ��w��k�%qX�ǟ<��'vZq�)	�'�Q��-I)�X ���.Y�y^k*����0�Զ�Ԝ��k���-�&�^V��|�g�Ae�a�(��l�\._��d����ƕ���ں8�}���V�����V�8"M��a5��J��{����Q^e����i:s��>�X�#	~��2������k�	vhȢy	��Y��AZe2+�Z��N�Ѩjr��g19;�T>����ES\�cl�fP����͟��2�=�j�秕�Vk����ᵒ�3 �9np7d���X���3�18u1�$���lY �e�0��̩AM��y�\��%��k%Gጒ0�Y�t��I0=�V�2���!^�o�&A���e��<��*�@�ư�V}���#������.�)�I?,m3t�7�� p���6�w_a�p.R"w)t��D�!ɏ�fd}f��j���V`�P�r�̼v_	 H��'Cv3H~�fP������K~C�VFާ�XXq��$�Ĺ(
�꽈�<V�
�EhZ2�Jh��؂����n�V�%p�]%ar8�u�C�PhJ�t��/�R�G�9}$��Kr��4����f���I�/��>�Շ�:8�4�j�,���~�R�kW��9e{���F1�˞�@8X;����z
�`�7Ԥ7�LU���x�u�$ L��H'}[�q0ۤ��8Ƌ9|z�J-�;M�^>�kLb�pϞ�S	�z�!k:��'ǵ�EId1	�[����"NĞ~����iO�hQ�*&	|�dN������11�]ey����[R&��a�uil)g�郞كY���3����v3�r����6��a F,c�`���
���Ca�4̣!y�h���� ��O�9/���$��..\�(��D�	/��x
��=�����7�e߲]F�i�5�����M������I7F��G�����2��s�x����K��N���E�'3��G���h��$I~8kJ6%i}��?x�r�c��}�yd�!�)�Cx���ׯ���s���I�v�]ue��&�P�g�${�&�ȅsm���&��%0�j�.8�_CG���`�,zNT	b�ɔ&t�c��,)�Y��4�)�g�4g^h8��5�J.�	6�����e�Z\���#��y뭷����� ?���$Z�e�=����$I���f�	tu��Ī�n�?�s?�*Rǵr>��)�4h��>�b~2��/�M�"Wp�@N�_��m_>z��ۻ%���!�P�㗟�Wt�kjǞ#=:���d���ƣd���Ͽ��gq�N�KM4*5�tPflZ��N�nI�R0�U?-��&v�s�q�sχ�q�Q�҇�q�QY�U-�����3�ƞE�`u�`��)�D!��*d�%"�X/�]���{hUU�mrJb-�%�WV05;&~�,�\���P�M�i4ww��F�`A]p4{�r.Hqm�Du�K����s����K��(����k5�З�M�rbC�:����'�N��dT�������������&n(!�"��b��y+�Ǧ�*x1�����-[gD�(����$�y��	'�ޠO�=�ze?ؘG��:��!�-g�U�N��$a�fv�3�QǢ�`H�`���}S�1f�1vK�o�6f�L�'�9IpTJ�a��ww�����03��ʱ�1L�O�m/�Y����
�˺뼜o�B�����Ps�e��z�BB9���Q��uħp6_�.��|Q�v%���v9��q�+�Z�"�?��	֞m`V���/#quj��&,���[���O�Ϧe���0��$�)ft��'�mg��um��	��!��nK��R�ez�GJ�wMιWW3���z�5a-4��!���p[$vFf��D�|G�р'��}�8	y:�db��%v
���Q�k��$v�e���ı0�׹����U���F� X�����P).tU���zK�xv�+䆴՝~B��9y��v
�PT�"gB�x���=�0���E�_��`�љ%B��
��$�)���[Wq��"�1��K��5!ؗEb����
�=���5�}9Ȝ�ŵ#��?�o�2� &CV����P�7��,C��5ǐ��r�2������h�t�
��|f���x��+XYt���|����<x�R����Uq�e�d�Hɦ�{��M��A��CS��_&l��){��:��Jl�'焜$A0v7������FI#��#M���I婲��a��)��aT.�mY���n�V���L�9���_ﵟ� ����q�l88��^;��~�x�����&���b�3`2�'�w=b�ؗ�E8TX �B��3���T��T_�3�V�X�*)C��+	�t�..�J�Z-��S�Ȍ��[[����&��v���2&U��Y*�/#��65�<�O��>��ojk	�f��ErH<,WO������VQ�	",��az�O���:DBY���%�!@�ds��"���~��Ȉ�YL�S��h[;Y�^�o@Q��a�<�����IB�ϊ�VRS}6�8�<驳f[eUb�V_k�U�n�u��aUC�9�/��$����e�}i~��|�Ʋ6�|]1�u|����{%x������R8�8�b魖!,Z�����m짳p�����U�U����fC�Jj-�]`�;ΪN��
`Uy�
X,#�A��ꓩ�wѯ�k��ji0�49Y�����I��QRnVq�d�v^9�$�y�`k�Tx�F0<4�����H~*AT�����̃b���Cb\{:<o��tN�m���3#*���H�i#3]��4�}"��9�Y��u��������B �k9�X_C��x>V=N%0;=���&�<z��p$�V���＃���vu��U}�ۻ	R��Ce�eE`hxH��´�~J�������>�}h#'{�9�R�"�CA`��V=�0�x��WC��ݬ�w�%_Ί���o<ӝ��Vu��쇛����h�L����9�Y'42�������y�E�r���ОԳ�*�Az_|�v�2�X4���V���]k�宄�e�)l����vB����b�F�f�͹s<�b�*��*�QY��N���.&R.l���ruM�)]�dEaa�g'����񟾗���R�pp0��������#w�n���-�엖״JO�N���y,����?����&�}����g.��)
�s)��
���+:Lp�	��:��i�0�,���`�ۡM%y̐��?���B�x�?��"����:U�7v�=m�k�ȀK��/]��ܴ�4tT�����˻pŶ����EP�s��HA'��`t���u::���,2�
]F`�{��d�����]���L�41�Uf����Ź)\97��d U9ƅ\ː�Ȟ�<O��2�;�*�Eb��� �,.`aƃ�Q/�CvW��%�f�S������ŋK8� ��̤Q)�y��TQ����Az�	���B�.6&�:���ab��'{���^A�SQ�G�!m��u�0�BK�l[�s��Np�o8t�5�l��O1�).�k�g&��h�x�^��^d6%`.J`�}t����\q3�'M����zV��7zyE���;�������-�H��(K�Ջc:W������Kv,���>����D
��(^�ڔ��Q&�PdA9ɀC���;u:ndJr���~�|���DT�j�hW/y�>;����,���k�����&ic��:_α�<?	-�������
�41�rdۺ�s�ǂ�:���[Gg����r��hI�l3�r�S�R\adl'��RɊdb ɨ_�ޔ�Il������y]��j"��1
��-�u�h8Ԣ�W���aO��8���V�c��򀛄/e���MN�1��^��(�2�^��5`��Z� �k�'v�\("#�sXo꼷�^7�:˧��i�Y#30�{sGY<�Ov����^�}��u8&��ߣ�a�N09�3�|@�o�c:6�u;E2ڢ �03��ZUpG�����'�dS0���	l���NB�����v9�����2������.�*��E%�*9��U�������Ӥ��VI���m95����#H%��/�����B�C�=��Fo���(�ҹi����Z�f��%`�Tf`��k������O?������>6�,b���x��<yy�hl�b�ɂ$�A��p�� !$������B�G*WK��r�C��+i����ZZr�z]���;/�[N��V���ɜY}�g��g5d�=���*ۙ^ʁ�ɆX>e<z���Gc���W/�����^}����"�v�>Oo�}�B����I��T��+�eD�fB�ԋ�f�c�\
lmp���NZ�,�l!���Fn�X���CZ���V��;
���l�����	TR�"����xx׫��c��(_R��DjV���)V��}�lt�N{]CaNP�s�)�h�V|�����duq/�!2�������>��I����L�3lG�����pwV��A�z���g�pɔ_G�f@�;�=��zZup��t����r�瀙�lZ���ўQVF���#�׫��La��Y,�	hI�`y|
Ҷ����7���.��	���2�ٲs���(�Ȳ�t]ݞ���&�sb\��PQj�q�kcgwS����T1�	�K�R�9<a1�!���ϥ��A�}��Y!����$�1�,�L+�V��Yr�VΞ����߫���q0h�W�tX˱�7�e��qPh24�{�ׄ�R�[�G`�Cg&���;�T���5�İb?15����-u�b?����
�������q�Y_�Lx�d^���iOc`���S�������#ILM�Է���
�%R�s|��E��й�����pn~�t.�"k�����ss��ޒ ��:�)4qT�`/#`tm�L/W�8�������f$�=��x��ĞZrN�/�����M��Xj��fjMU�셸��!ƒ>L�0�����Kk�y�� >xA�{@i¡ Ԑ#zU3�r��q>�lO?�ujF�o}��8��`b4�}���$�}�#Ò��¯?���O^���~�����	Mp0����l'+ΙA�-u�f>��h|��`����3lA�6a��x�� .��o���_}�\��+$�{�rU���ڛbs�ؐ�F:�]|��Ό�p��y&`uC�X�3S����>�EyOM7r�:��?��q?޼���߾.����`Ŧ-�qO��oh�Z�Z�h�5fkma��B�>9_`�湏9y�WkGHآ�H�k�l�N�1r�ʝ:��~l�$���|@2޹i�Y�(�Ć��ח�P� ��.3#q��0�<:���k�	�w����
�u�,�ѫ�5��s��n��ϵ���8RS]y�eޑR�\Zi�ꧥ����ɐ��ɘ�޾�'k[Z�x��ɝ��OI�v�݋�|iV�m�BA��Z�!�>���0�>� >	�r����7rp�Õ+]�a�R�BH�祥Et	�SdK�#]��m���=04[^���~	&��Z?�%��V���VHH�S�O�g���U�z�T�m�]��rZ�l��}��	���m�??�	IH�.�V�z:�C��3���bhP�	n��.^�ob}m�隬�IV@�����P�L����>_��M7L��㴩i��*`fh���Wi�w���$���~�v���p��^�C��Q��_��;�&�����q����y�⚒�?��)�,<�Je5����x�{�S�h�WclzR��8���宜��R$.��ڨ�l�Gi���PB"	�%1?5�AbE�I^~.[*�\г Q���LUHWé��Z����X&5�e�q��`���~�����V�ԥ}��8���~9O62Ţ؄��.�5#ǝg�Ǯgf��׶�8��{_Y��|�,��H[G,b���)L��ct�/_�\S�2�����A�/��gr9�"A	�SX\��s�FA0)gy������3?	�H�$~?!�Ҥ���!��,��G��2�-��׸^���[�3\��Z,�Y�|���f��CɈ�������Ye�N�JI�ޤ�nZ���U�����B����o�vY93�h�X�\��Mk4g�i�:��u)+��kɽ��ɝH(���߇}�E.L�C�����B-\8�o��\K�C�^���U�n'��׷�c����D4 Q:����r{ey�]���A	�H�˨�a�&5�x��/cE/)���I�^�A֐�J ��bFC��VRf���d5$��)z��L+@^�lk��n�Ҙ������s$w~���Kf��2�}����]VD��r��_'B�* +Xb�3�,�6^����+閇���c��@"�������l��M��V��}�K$N�a��:���wS�5I�@������Yܸ<����B%'�ۧ�(���O#J�%@bS�?g�CQ\�0��Q�+�8��A1W�C]�<J[MxA�9:���/˹���7�Qp::<�Xįd&弶�p�~e�y�U>�kHi8ߦ�Zr�}����q�r�����uy�4C�8���q(靜U_3�,f��V��~&ǡ�d�m�Y"VKܚ�� )��Ⱦf�"�?�G��Qm�c�G�E�	
�=���~�`�\�c�����f��>{���W���RD�n]�>�+'快(fsb(MBbx؏T2��C�c�P׀:!_���F"-������C5��-K OV߁�)�o��|�:޹1���7q��]��k�X,�z�#	e�#��Θ�h4:�dG�g�E�d2���$N�D7q3=:r�۩8���t�l�R��vU(��]��e��ZFYV5H�;3[	�$๨��E��-�M ��F�\54IQ�V��7���G1�Y��rӅX4�UV:���B�i�^��M�U���F���/��\�Aԭ4�]����*g��l�\C4l��C�o�!5�({U
� Y"��x���LË��!-�<0>�t:����������6�8{v�řj=��jd
:�t��][�_��?�^Ư���'��G7$Pg�V���R��>e;z��;Jހ�j�ʹq\^����Z!k=U|�p]� Y]Fl8���s���=����v�8����z<����)$������ �p�,~��kH�L�����#��	�"hRX�	�:�|��iE�9-�ܿN'�2(lU��s(��>�/�y��=��Ocj`D+�}�<	KWŠ&P�Ԩe���������o����݇�q�������W_ྫྷ��w�J�}
���b{��4��`���曇�oTy|~�k��=���Τ�������Oa7+@ue��1��s4�~��e�[�"��Ύ���0f&HF\�#nsS�x���_� ���+����f�[ˏ�����������n�+[z�l��TnhB :�Y��-$ba	P����XZ�� ǋgԃ��a;�C$�.���ɥ<�&bH�@�%9�9q�t!o�*sò�Q�z9��r#������ޓg(�:�D1�taԱ��
�3S��k%G���m<����n^����_T����إs�0�BUl�ݵ
V6��5�������6����2�~���F14>���n,oE��Yf\>���yhR��3Eņ���GP�����F'�Fգ�-k*�K|f�Ջ.%~B&I�2��oб��$l���
��Z�$���-\!V�[=��e���������x�,l{��i��1̉�z�Zƽ�/q��aX��	�n�id���T�
7��z����1��S�t\hW"m���C�Ih7$����\�<��'r T�QUl0�Σz�}�NK�VJ��Q�$Y$ �1�0�qO˯�,���Sr*[ɢxaA��K�VAg&(Tή��F�>�c�����Ҏ	2t��Fq�� &�B������Sc1d*	����~��|
r���ː��B��r.3nD�\�q��-���\�%XQnn
2�ӯ�"��'�����6�>�UB����=?�p,�W�q��gP�(�qt�Nk�٧����M���w���i��l�u��M�cvf�Zw�D)_4d^:��ұ���y�[��1"��G��>7j�jxNOOaA�l�RE�PBY��zۖ?-�e�����gd�5���,�u��t�%A0���Jh�AӉ�s���q`뺇�mDRQ���3{��ݐ 4 �Rl�����&��C��j���i��x��L�����0���w�;�159��Y���v��9��42LH������=�п����?�0��F[υ�x�am�;��"[V�����8�SSx��������8Rb��q���]l��bC]]��̢,�g t��花�p��\�P;�El@RR��lb����4�lwQ�Y�k��,=($����ʦ+e����j
����@�����]2*��14*/@-?V+X+��)F�*��;�ɶ��q{fO	nj������Ȩ2\
Y�Z_ǋ���_b�uv���������1��u�i��F�v������C�8��Ο�E2j���#�-�� �a���Ƈp��Y��r��%��փG�G9u���&P���Yl�Q�`�B��B]m� -��B"$F��LN�
��kПB���#�
1�U9G!���6�[����� ��(�k�f��}�Y���a�th�t�g� ��-��0M�x���xM���T��!v���g����|��l� �0v����ƣ�U|�:�����}�MS[n�F����+Jf��8`u���5DL@��^gg0���]�`��^.o��P.zǧ�=l���p�꒜'7�| ���>���̨3��qii{�Yv?8j�X��0[����Q�y���I�����:�:ۭj-$�:�t�m�TwZ��)�M`&{���JR�(�e�bg'�ڋOǽsP��8���D{�AgH���~��a�d�)e`:�iu��Ke˵��4�N�����/V�Ά� ��g%���k����N����W���9����� B�	yƖ
�zIP �[E]B�0�Cl����e�Tϐ3;&�q��z���CAly#����CF8Z������8*␙�d4�h�|ll��8��%/�E�)���!�@!S��� OvcQ�7��iG�E���=���R���r6rd������Y_��� 	TQ�p�I����f�Dʑ8�7�-���H@m#�S��/6��Pgt���䣫��?���ؕ����B��`�->~4*MmY#!��k���`Emtϙn�q.���q6�k�%�~�173�'���g��_�p\��w�ཏ��շ��{����F֏��m�޼��e*��%�s��v�0�J6h� ,MR���²�D\�%+i�����e��e�|E�dJΐ���-�^9?� y��hB�dY�j"�`̫{9>�`6��Ѐ>�`2�o�	(p(�@2���F@\�vCj�2����&�|�9+~�><��euL-!D�I�5�?c8{��m7��~�b6�� ���כ?�?�x�����w	�o��g.j�"����z�	+��s�d�hgn�S6���p�"�:�A��Z�Q
~o��ŷ����o�o�ƽ�˸v�m,\8��b�V>	~HE	�@У��ԋ����o4!Q��^�gZ��̾l!#�HC�M�3����a���o쬐{��o�k�{#א��3�
�#��T g	�B�c�΂]/i����X��Q*��ͣ�yZ�����Tbjq�UIs���GG��ة���E�\�$g�����{��u�N�x-WB���$�y'[�
\ͲnܸtW.Du�@p/ZIzX��=�J�y�U92��(���Z��6)"I�S��X��茵�R�ʟJs��gXF�tI�g�Ij�iU4q631�3h������M	)���ˋ�Д�/�E9��h��H�c����d��8X��x3�7���`��t\�P�U�{�z|��:���Z=���ey^Y�(L���e	�GqE�X�LZ�#Tѹۚ�I�ɡ�FS�]��D��3�Ю���yu�eD�h���쏅�sS�s������>����4c���jh �3eZ��h���a��M�������چ�j @�f$ù���XпB���
�6Ɛ��	rMR�T��r��[���:#N�I��t�)�@|A�A�CB@������W���'8��ܚ��VcS����DX0Ī�v�����l�_;�ǉ�84:�^�>JF�.u�n8��n?f�cr���]����lj`H�=�̧L���
~��Ĩ���n\�hU�Z����vK�2�ᑄ��8fόk�����g�/�d�-����q��GI��GJ6C��N=���7H�L܎�)��4lme%�U{ۑ�CB���tJj���[��g�)�A�퀩�;����g
�.븓�xƉ����eN�Y�k��J���b_F$_�F^�g�t0h<wn^�[+/�U.VD	ጯs�Q���9���Ы��P�8��8��&�Mx�ů�Ñڢ G*����g���ƍkb��᫯��'���h�0;;�3s	%P��q��l���um�X[y����ϟ�v�tZ�&�����X��3dX�8G�C���DL�3[L�bblT[I��Ǡ�����,]y�&'�9��2��^� �z�A�Rh_��V��ʝ��.���z)�_���)�Hb������<Z����pFd�0ev��z�uB^pLC������A������,�f�0I`!�m2��=�}pG~UVpT�c�Z>�&�n]���zb��\B����jf������%��AY����Q7��=|}kU�Eϟ=Ū\t��L�@����#�����KS�䝖�o㋯��ה��A[�������x7�U����8��� ��(��y���X� �6B��ήr��e܃�UBOٖx��B?^oB9���Ձ��=g�T�f����[����N�����ƍ7���Z��"10�T���g2�4��<�2=���}Z����٢��9�����pM����ξ��$8o8b�B�����07=�����q�Q`Y��X+߯��K3�����h��{��;�\"%��ܹ�"���{;x���e���i1$�{�x�M�I��S������RR�8A�I��Q9�5M�0 �u��\�t��&�0i�Z�)x�W���;���s���'F��Q�� ��[�g%@�N�C�u���-VW�5:\�mde��[�egSZ�r�޾qC�x�}��B�C����I}��/���	���ԣ:��6VY��6়���X���H��jw��&�3�ŗ�6f�ӯ��	��QA��2���������z��Os_�\Wg�_�*�"Hn�5����2m~�⬮��,�I*�6�U�h� ��~w0�f�����?g������O)ϋ�@����.q�.&d�sԂ���OZvS�+x�(���~�p�#����j�H$��Afa	`n~<' Z����N��aU*����LMPu�*7O���YV{�u�m�}D~
m����B�������������������B0<"pJ�A�C����X�tJ�$�$����~֪��|U@�O﬎J��~_M7���Fm���5\Y�������Z��V;���%r�C��?��x�¨�lMK@����B��?��Op�BR��[{=����_��O�cu[@DK��[���P?���r&�G'0�B���g_�ċ�m�����czL3��
�3�� ���Lx4p���#l�� +��y	*��C��`H��0��R�u���[Mٷ���{���y!��cXM~�p�o�5V��3
�N�*@��i9�?����CU���99�Y�ht��Lͳi�z
$զZ�)���ҳ3�<ӣ](^C�n��]=r� �qo�m��U&9��q�2�[�Y�Su2�%�J���KX��$!��j 
��z�2��OcF��1rÚ�Y}���CV���^�[.--��였հ��[|�"��ؓ��lmFʞ�Tی��z�m�l�Z�(���Vp��E\�����e<�O�������'c��8��sŮ��rv-�Vٞy��!{�V(��{�r�2���v��=�E����Jv����_Y	��GiL�T�(W������5�=$)a��3X��>JB�<���j-<����~�6l���X�0���z˯�qqq7�(v����^*�d{�����DV�КM�Rʚ���n�E\���3	誅�쿍�lG�hM�Fl�6�0*�6���=���GE	 wq(�c6G⽐�ǐ&����t�bL1F;�$*G�n�i�$���9E&�����R:���A�Ί����ةC�t�̏2��Jm�g�5�8�{�c�i�;�3��1�F�s�-�p	,���Li"�`���x�݄��ǭ�*X�2|z�z'l�lG&�v�>�h��L��5�����G��|�8ܫ����Q���X�	vc1�����W=�L�s���#Y��5��hr[^e���K5Ե0d��w2�=	ig^r0)>-���[;e�T5a��=�S�n+�fPjk����.^��r�����:���q���&�����F���e9����7s�v���o��E�L���.��vh�����!H�3<�~��졒Z%�	�7	��$�΢T� O�@�s��\��`���`���A�{�*]9[��d<X_;� ���lDR�g�n�hW�o�y����c�k����M,w���7��li]6ҏK�t�m�փ�.�@]��*^<h��~R�r.+����l_w�q��+Y�f�\:�	�>�fm�nI ���E,-c�,��᠞����J�?X�\�7<(�����+ƥ�,�ǡ}��P��\�t[���?�az��J�;=?���	�6�8w���#�\�pI������*b����Y����ٌ�S��[-U���g�_*Lɾ��;�.�㉀�~��]D,�%h�:Uk)[g0�l7�H��࿭3��(Σ%�Vobrd Ѥ�vM��9�RQ)���lMg��ߣ�r9|ؕKA���պ��d�_��a�%\�� �
�G%X��3�Mr�������O>Y��%|��=��)#j�����l+�8M�_���V��{9i���[/|�̽�j�$>��s���o���*-�p4���/brn��(^l��t������rv���=�ӣ����>R�Y&dX,�f+��`Ťf���تt��
�����DId*�"Zl��uTd�RP+N)��%͵ =u$�x�=����O6��g�atb7�{�rU�~	P�2znl����h�{I�d���r�t��kZ����9���!�;68�wnL�l�g_�#J�ڸ�r�E��G�e -+�mq~��9�.�f�L ��q;�c�2k;���W�2��S������w_�����/_Qِ������
`��<ɪ�3�j�@���v�[��~uL%�zfZ�v��_CU�8�)��H��ֽGb{.b�RS�0��}<x�!wgf&0< q�E<��Gy�PB+��hH�|H�e��2���Vy��W�=Q��� �j���d��K�JO��,�QÍ�NV�"񔜋�JqPh�"� Ŷ�%wʺeͫe�6w���w�����A�����_୷�$m��/)[�I|�luK�L�V���,-���J��+!B�������N[���h0�2��o�.�����ַ�J����ك{k�OoJp8+������IM��~�?(?c+z�w�<�c�	(�Z�wk��|z=Z�T�W�b�W+�\/W/�͍]|���
(��|����(��:�#�q�{c#a~��u�iq�#�����0�а������ܫ���PF��|o����H�-w$����W�֑�U֩T��}���$
���{���u��	�(������k\�����o?��tF����t�|W�7�?�=&�*U�:�|��#��K&h���Ұ^�]��5V��3uf-%�����+�8:���W��/"t��z�̼��ŋ�Е`�DY�VW��\F��yN%�i�E��dt�l�����Y"�ߝ��S�I�1&�\J^�U}���-�S����p������� mOi�Ͽ��o��o~�)g.�~�%�sbd�|4)���9�$:��H�A&�PrW4 �hS�A�{gI����m�Rk�ًm"����4`���ɋ��I�$��Y׊�+�6ъ����J���Tˠ%�<+�@��쨰]*�����m��0�D׏cQ��8wO��zFW��u[uM���x�{N'S�Z�i������3�K�����llb}}K��^oC}�2�
8��[j������:?���]S�rN�zQc��l�U��^m�X�S}[J�y���(lw
�{m���a�(wx �PX�-��B�P@�(���]T+-FtH�(@��b[��
�O�W�:t�͡X,��w��b�S�˴|���.��Le�R�-9�2<g�x��7�l�m\�|F���L
Քѧv����	M:�B:3�iȾjEf��r��H�r9�j����sXd` Ր�62+���%�J��w���E�<�-��O�	3��s*��R��O0��U�3�bP����A��,�(��AKpz)��D㵫�8���US�乗.���d\� u�+b+�ڥ������12�R�;o0�J��m���,Jb˪��ԌO�bN�H,�>���}X��,J���u����+~���l�5�d@�!�an~�'b��<��s�!	��|�&&'úv޴�r9�prD�٩�@L�#��5�a�'��)�a�̀p��԰$��HΌV�g��a�i;���<�l�{_R��H$Qh��N�p2��o��6�"3ā�ߴ�K�Pْh�-*̎4�m��%bp��uR�B&�a�h"��$�B�3$����)�!`�b�A�l�L��O ��XD��z�f�8��k$l��l�[:SD��ճE���� �~k^[AW��i��H<�����3�P篾|,-��B�%�}Ƈr��Ɵ
k.�! df�vv)��Vџ��o�c14�l���E�̝õ7����#�9`u��D��62y�HC{����%�-~,�S�7@�r	������r��<��6\@�aF�x���H%"�u����P�kd(���i���S� �a����a������H���"s���������8�C1z����0#�] O ���1���ٺ���m�b��K���b�}��n�� �έ�P���W(�$���)��e�vyT�5�Q5���t�g�1���*�}̈��A��ק瘗��2®�@�P.[A���v�$]��������0;3�����~�l��h������3(|��N������g�I�{s���6&&S�|�"663(d��x�M��Ֆ��M�̌(�ET��j�Bs��M��	(>#��F栉G/v�0Q-7UJcp8�ɔ��Ie���ajf+ki�Z�����~�C14:�Ύ�}a�l�e+C��ߩ�q1���?�V��D#A*u�I }�ڿ����J��r^���+~�]9ޞl�]�j�#y��(c��Q&p������0��}�<ωӘ���3z����V�U���afv��+=&�k��9�L�e��c8�載��4X�8mXy��av&�/��dO/6VQ��e-��������&A��X]a��:J�:B��J�p����6wXԑ)V�z�i@�]f2["k\����*����#w�)v��ɩ�6S���L0��VT9�Jp�Yk�Ǖ��7�;}шr��`��_�\����y�?. N���C���_��/4�A%yo$�`�h������h@lK�,g����C9�Q4
GL(ĳ�Z�=CE��>���Uǝ;�h'qiag��:�900�������-��4
�".�P�zZ!��3q���P��:	HB!���1-�Z�䜍���/�AH�H@-�cy�[�nK�}p������ʬsJ�ɡ �_H�r��CT�Aq�Ch�ʧ���OQ���{�b� ;��he˒���m��h�j��ӆ ���N1ȥ��L'P�U�-���*d��L�CCCr�w�ןޖ�x�]cb~��cL-�A������jCE���=�*��bv$�[uj�)�f�6L�m�^�S���e��5�Iٓ��Q����?����l���[�.|��9�N� )���:g�J$�$cL MK�Oؘ�n��t��nM��qv��(>�d�k��4�=��em;'�'�sC���H ����*)35��p�6*�g��;{�x��.�ϰ�I�"������:�����k��ʝ��"�߭	��K����gG⻊���G�ږ�!�f��@a�\Ҿ�xZ��DM���V����%�[�_��H�=���"��������p��y�.l��h�*�){e�+�t��ܑ}fe�Eٔ�������m�3�]��֎��!��W�#<�[�ia||�)���18:��q�æ�@���i��Ū]<�y���߇pl'A�Ut��>���1d��ە�
I PH���WXY���|!���%~��+�z�u����A�k�[+Bw�l�l�E���ϣbObx��;ۑ�����f�ʹ�X��jQ�c�Q�1A�h9Mb_����ڤ�v��" Qz�g����0]��BAbx�hYeD��$��+��=-j@�]p�ߥ4Kj �RH��W�IO�XAgOU��2zs�5g���2=3Bý��#����ܟ�ȳ��jW��`��޻�+�clr�e�{nY']����qvьO��:̢f\����`-W�x�����Ν����W���?���8bq�;e�z��U�`$�c]C�HXb[�]ɉOM���R�)�]���D\<���M��d��֔(�R�)������4� �F;��{9d7u|�X�Ԑs�`hl�ܑ�^QaѤYU?�N�j�8�="��$Й�Q]\�@8!zQ�;�e��9��R�ж���`:rE�*M�/Q��t\�����x��q��ޜ�b�h�u�,�	H����T,�buH����>�31�Ų<d�(o��W�p�ʜ������R3��p�
�8?1�b���1�e���]�&)�)���`P ڴD�זbL"D
V1~��~��2�wK�|���e9��A���-ոJy���~��o�8�U���1����+����u�������$�[�+�S���3��Z�3��[?D��������V�[��Jb}m_}��5��}O���e-�R��x�m*��r�6G˙��G�����󻙵�i�Uǽ�k�y}�|xM[	���lmk	 ����0�����;�	��5��/-M����Q�K����,��ZU��	�]!$�C��b魳�����׷p��8EH�_ mO��X>0[<5��PK��yt�J�C�X��uVN�sᥙ_��A	^����u�=J����U5
WK)�{F�2����@���?׋3C��a$ą��;�# �狠����Ǝa�{
��<��S3hv�ܰK�Ew�����f:_�Z�+��Gy/U	J/o��~�Û�[�}{�RF�����v]�.����َ��F�ѩ|��%�Jm<~Y����\����š���<W ���᩹y�wsR����6��x�b]_�|E�é�f"����7��e�Z�hk6Yj6_F�ƙ���=�Ӈ�
��mw���A@�p\��%w��AMtH�.����6g�ón�9kd�Y� R�H����'+��J���G?���я��=�����M"��`���A���X8���g	X`��v�T�,+ʘ�Ѭw�� όǐ4��tw�H��j�� �؀�U���`8 v�&�l^֪��[eet�����i�?/�1W)���iB.��g`�,��<
����+��;f�m����^193���9�6��wj�F`�3+�KT~Fn��̖�ɗ�*��
s[���ʾ���x����R��/���&�'G�\Ɔȳ� 17=$�Ņ�ί~�H���W��9�3�Ӄ�Ԧ�����o�:V]̇ ��\��~�o�_���U ���gO����XOk"�Hԝ��>>+}���6I<۰g�ڰ���Dv*��4s���Y��Ae���:/_)��l�����Y#�F�V��k��!H��P��l���æ�)y}	Z�&fUǰN&Wv���e�Z,8��W�6��a��A���yX%�u�ʽD�Jϯ��v�9h�U�P�@�c���7_>ē'Aվ�k��W�u��� ��:�#�����B*�RQh_؍��\YUR��v���SImX\ǌ�̰5��~�{x��9��ç�x��/6:,6�z�Ie���b�� 9�r�̘���1�۩�%�3�۴�r��R��攼�]!h!�2[ߛ�
���r4ѐ��������J&D[ד{ѓ��`+��7�����I�/�%��]p*e};���.V�=�a	�(#A����2fu��z�d�kռ�	&{����r.�@4;���I-�x5I�S�P ����I���x����F$�r�`p@�Zk�V���+?OR�.��m���
+Y�W�E���;�q����D��{=M�3`�-ϓ�8C�.g�/�"�*�IBD�,Ud?$�'a^(����rt�3y�<�j�s�_#·�3�ñ�����mNu�Bb�⺶u	�f��0����h�����1�?�S,�"2cG�nQ���3!��<GG�JG�,g�Tb�k4;��5��X�=k5L7�E���@��d�{�uw�*6I>|���_�d�!�91�sW Aև8��C&s(�>�%��#{��I�Mh[����B���	�����T��z�et�u��c��}�����ݿ�B�xP�%vl���nJ�ZB:c|�V��^�il�IȾ�c���!ѩ ������z�JeG��VY��VWw�(�o�G�~딥kW��FV��ٌ<o�X[��7�s�[�%l��j���C}F���8�$l��P�;���J0�ge�o����iVW5`���GY ��x��KMZ�_�	�������������J0��� �r�7G�癄>8<0$W�F�xU.�d~u��nwP[\���􎙴�VʵM�\bdy���1-�>�`�k@ΰW�	L�����	=c�|^�9�#�a
F��G�Ω`�γcCk��K"�,�Q�xa�/Mȹ���T��'#:+xn>.� ����t(���葉��!�k��s���9���(%
+ۑ�r�f���[��d�e|woY���<eٸ�T6Q��/Q?���#y
C2PH&B8s�v�6d�BX�pVM����Rֶ;5��)�p8�d��@5eѸ��Vf}��2���x��V�d��y�'��g��c���..�>	s�>�@��� �U����I�}�m�N��XS��&zj��e|�]g�do-?�g�����$��g�:3<.e�[�K��Z���.*����-��r�/7q�iHP��}qzP�Kp��%�2Ɣe��k�<��G�ڊ����LI����ȍJ�f��e�T��&�ɸ�ߝ����ko���L{q����1���?U-��>� elm�(���9�4'%BĘW�U�@l��K�ϡrV�;�����`kQ��ѵ���(�8::���Ź��A��e�Z8{fВ3���efO��}8�q�f�����S	���6ٷ�>�4�Ưq�+F滇O�-���X:7���d�����10$ �]�7�3���{� �$Х����ǫlg���F񨁮��������Ւ�7[X�ʠ!�po[����}V��+#7<��G�V[��}�TIGMr2�qv�.띌S�1���������E,]�����_˽��=���N�k�,a{�E��FYqC�G�'�qY/^��h&Ͷ��)��+�]'��j�0S7�>�&	4B~�[~�� �I�A��
�O~�SL��������f�����qv�n'jdI\ǳ�.�RȯiK�1ȹ��3.#&�jAT��=�"Qв�������>�����'�$H����j3�����`l)맥�X"���E�t�H���HpP��E���]��t0��3  ����:�T;�����8,/��%�v��n�4��L�#�s���2�&���LD10WfȉQ	f}����侏NYX](�S�6I=�h|�,Cu�c�1�v$���8Mz�k�p��ݹ�o��N+?����/�zXcS%`�П�Q 9�$/�2�C�(I��F3��T'8�jZڼ��,#Ѱ�:�v*K��&�١�z�F'�q��Ye+���L�jGوI�D	�5�oL��Y����Vz���ztv�zf��Aw��f�,��f��X1$�AS�[1}��H�cG���ER~W���$� �~&��(�8z�F,&�<2�W�i���{<;6���&#�M!�:_�m��a!��6�^S�$��ԞK4󷬩c��~Z��&�A�YF1��'7.���7�����rF��pL�{n�/\U� �� N�qӚ�z�-W_ë�w��e���z�mtƩ����.�� �$(I��.wq�=� 4���8�g�Α�,���� ���Y�[�؞�j���]%��G����7lC%k#uU�р�^v�f\�
��U�f�J��Z�{"8��	k����$��9gƪ�������J���4p[�_x�QY�r�	o9���,���my&�A?�ǒ��{���
�]v6��T�u��P���cG��Q�e�u��we���a�-�U- ��/~yS�R���_�P!ʚ ��0[�7�A>�ab��6Qv�\`�zN�a�i��9�W�՜��9t!�|y^+����������.}�ū���n6f��=f�e�Xܰ]l�jE�h���-��FU%���b��2�\'vWY�4��q���R� �
��)h '{(8�%�	��~^	o��F05;��P,���@�0��-%;� ;q�Kn��P�-#7�3�k�N�dd�Y=�9\s&��&Ƨ��#{��ui���rx�tMp^�I�`��� O�sj��Te�:՞j�����Oe��c	PgR@���p�xJ�"w�*x���N1��_����2#6��#��0�Al7��9�����/�P̯���L6��Q�7�kU+c"(���²��;GA;��ڈrO9:��v,�o��%��ְ�lG�LL�#G%Z�ȫV���ɿ�ğ�1�����`�X2���GG-��f�T���	�qpH?٦����;�0�AB�r��=��/�f�H­���'�}�|���2ι�V<�"۱�0a�U�U�)�#��ސ�`��D�G�_�7��2�	(�5���=l�"Wh�k�46�5��`g���8G�a� ��\�b�	Ry��:*����9�z��RV"�b�\6qv>qV���wLː.+ef<^�8N�.�w�ٔp���Go��_�5�x��x��œ��d3|(�
�^�vDt*��ff ����BK`i�	~).�=>�'%r��׏33�����BЪ��� �%p8g�H��Ҭ��x��@f��>��6�dDz{�2�V�~U���8��in�к#���W�����(e$�'��?R0ȪГ�x���bY�4[�K��PrA6v�X{U�b���&fL����z��a���E�/n��U�e!%N���n�u]Ze��6/*g98 �l��$O��<�a����+��W9w>ĐT�'�ב>82���C9�1�6L*s,��t\ ��O��͈<پS�`�?�����l	�؎��i���'�x�]�022�� a��\�fv̄��w�9���H�nW=΅��Dm*u!e�r�Z4=[�A6S��� ���q�w���^^������t�C��ds��??P�Ӑׯ`7 H�˄�f�.��L�~.���Jp�&e/%ЏI���7��uf7az�Ի��b�� ���P*����g�P�j�*w��|qO���Cm}q1�-`��d\ژ�ٸ|����ʹ*�R��7��
��백�;��
.۳�~�����s��O?�o��bt(�k׮h��%./`ϒ��R��|e�jkf��>x�K
Ӷ��J� S�Xq�۪A�=iE��L�Y��OK��(Z_���>z'�/?�E�B��a��B���+^A�~���k@~/������YJ�����=�n#I&K9-��RCJ �h��Z�����3g����hyM^��h8�����P-�9�0�s�F�͓6$NR�65����zE�t�L$�x�"bQ�y	z�v�t�KlK�K"4�	U�f�8����k���	���
���&X�|�5�7+l^s7�</�"�EA�SAl�S�G���`}�$�UK3��L$��3�t*��@ԑ ����ϩ*뼙�?3(���U��~5*��Pk*�y��Qrj�}�v/_����� I6�zfX�d���Z�$�W����Wk400<�T��ʡ �� ���A�5��# ����"|jJΊ�6VT���yu�2����ڎv��.�F0ͤ[X�(x��7��Zu���p�&d�~w����#�(����*���
N�~y-&_<�,�S�a �����J��L�
��,���VG�p#�|����݋J���9�C<	 �ur{bO8���RlaV2���2�1FF�XsʪP$Hb	��?����{�=m)ѝ���LXȵ�fe%��zi��ᗟ�c����Q�a�[{������p�-��ʀMr�Vǭ-{����x59U��o*~>�(9+���c��ɸpԧ3��B:J��S&�.Br�u2ˊ�[�h��Fǰ�3!@�^��=�szC�L?36��HTGz"N�P�����w��RV�RB)����k��C�z'��M���{rv���я/#w8��4���f�Y��9��H�"��,ϩ����B��Ծ�N0h��U���L�Df����8��3E�.�Wz�"ǖV��-e\���K�x���VK�"}��SӹT�^��A�eCF�q�#X%Q��P����ݤ�)��u��g�/�9+8KX�ٲ`����r��#�l��!e�o��(&�]�����f�@�K2z�ueS�>��Y�u+A`[T�<&�c,�|��X����?JAy-�R�rS,��x�r����K�8�.�Y WBG�^2Yy��i#�9x}�L}�cO�8G�����}�W�z��ޓ��<񛹿��,��$Ι�X��ܔ�-66���rw|�%��J`��mk座U �)&���NL 2�Il�ʽ�ͳ!�ni���מe�<��ڞ۫	�yF\�0�]*��yz�EU7tOb�l�D�[=�\C����Hǵ�<(�btpLS�`@��a�M��:�T�q~G�u��j�2�w�KI"]�08$8�|(A��=Ι6[��L;��U��m���@�>Q$��u�B�V�R^�J��4��HJ+m�B۟~�xB��Ӷ�F7�;��p�[��M���:���}��a��f~�ɸj��Ph��/�G���WF-_Rpٵ��<����*C �P�)���tv��,�.'x�C�ˇ��X>>�Uf�wT�C����m�{���#��C)D)�,�(��ɱDnL�"�B�_�YF�db�9��Ke9�4�����P�mJ�A��D����g/���-\]Z�l|UkE}C���^G���N�2����lp|ɶ�}��<�����Z�u�Wͅ��\� j�:8f�U����y�*V$P��x�JC�G䙹j�]��F�@~�_�' ��(�/vR.�8Y���QĺI`�4t�,�sn��e%§��c�r�]ވ ј�n��P�b�>m[�8,/ �3��pk�.�v�H���4�X�Mkpp�|��&���ӳ��D��v��� v�(l���`o1yf�ѹ��*��螩�h��Qou5�G铁�mxO#�3��8�+���P`�������iir2.�a%�1m���t;���V6�.���5d)F�����@�ZC�V��Рfr����ta{�,�$�!	XK5�I����6���=�X,��GJo����)%AM�;��C�,n��ka&�ө��e������v�Д�㉫A�Z�;M���(��×�lhu�����ن&bb���G0<�R�ʹ3�I:M$=$|�����N�[ޛ�m4y4��A��F�B[2��vi��e
}������1V�/kKX��P�ª8��и@b��$bI%h1�/��Wg9�v,a��U��6Κ��=ت�g�͌�ef�ɖ���3qb�!����8�+��x�~0�e��AqVҋ�0d���V:�9��*�g�SA����1�\�$w�X�� ���\���|D^?/gx�¡�Q2��E���.#�K�<7@i��zx�(��^Y�����?������ZE���B@0��dWg����j��ݗ�`"]�_.���Z� J�z}a��,8�^����e����\Xl߄V�v�q�o|/E��!r���z�'��3K�ܛ����e�]�}��ɦ��c8�Վb���������H�Fh��XiW���}����( U(�By�U�}ޫ�|��pfG�h�L���Ϟ�����	���N2�Z^F�2�0�ȵS('�I��Ĕvv�������E�ڔ�R)u%`�����4)+sV���1�ބ}�39��Q��$�f��it@�l�CY��W���K�@�|�M���u$oI�x��<
��X\ZQt�W���~}�J��5ern�y�kʚ7k���b;)���r��'
(���?�wu� %ϡvY�y��ePٕ`�'����S������+h�ڒ��)�3����ztt(�sk��'%��ɺ�1:>���������AKѦ/��]o�Bu���z�c��I&i�8�W���@��~O�A�Ż,�����=Qy�3y?���w�K��J��m�]H�}��lU�l\�G?����.��m<�.K׮.��OvkyV����+2���zW��W��d��[w�kO�8�嚹u�%�#D�ݥ��T�b��!�μ�����֌I�]��XA^Oⷼ$�}I܂<�$���؈M]*u䌱P�*�S@������'�'r�aJ��(��Ui���P�PV�n�`�J���-�&�pY���c,�Br�z~E�8�z�4H�~73����t���<MK�h 3ɥ�ו���	��ښ���>Q�<��<>�kAB@m�#G�s��G�1�ZkOHFQ�Ua����b�H��s���pV�&�ǏC��.ꝣ�<�}���I�Kƹ�c�(,�-W�~{��������8�r	�W�r.��;����jr����R��Og)��x�AkI"6Ca�b��8F�]fD�����~��cdAE��'�q�J��%�����z�����at�A�����,S�e���H�"Z8Z�|^�Ye*��q,�=?!��;;[����I#�:[%��Q��r���|�᜺��(ae�麴-�SBG֞�)�%1$�kTB'�:�zM	�G�Bw=�c��j��G�!�G]-��A�~]�SA*����4r���-W�6�qH_���[��@D�9��L�~��N�4��
�C�˼Hb	{�ڴ���!���}�Xn�X��Z6�mqɟ(#Fdܠp���:M��u�P�`[���V���q+@�vI��QL��k0�tcO�P@���f�Y�!-uT+(*]t��ѕC�I�d���&���I��L;�9��=��w��є�!�!)}�B�������xL�A}c��7�n���Uy����ڑ`��#;5#�'�@4���8kn��59�ۦz�d���A���
51�4��VBi��Mq�}[/���$f����`myY�����x�t}��Y۔l!e�Rau%�X����Nag��h����aayliƒꥲ�vR���I!�}q��:����[�16���gh��J�v��#���u*������ݘ����8�"; ����JG���t��EЄ �זKG]�L:"KT�Q���s�g
I��/v[!�L�5I��c%���ZS�y^j�|�I�Q�Kan$��_�L	$b���j!��Ȉ��K���A����e`����,W�y2*�N�3(R��N���_���\5y����ء��Y�@����  ��IDAT���0r�!�m4wɈ����ٳ�8�c�׎�)��6�2��d�cr'B��Dr۩�#��3��y�kc���ao�$R��}wt=UG�:Y���}$�*1���hX��k����+s�%[�_��#{$g�+���0��89*i-.���:��#����صHm��l�'ki�ņ���qbG!dR)\�0��g
 @���L��$�����1��;8���ϥ�i3H���'B��HX��JC�I魔�I6#�peo�9���˲w��\u����{�����->G8)�Kϐ.m�d'RY�䞪x�R��u��N�R,Gr&�ȹv�9?�qu�I)]:M&��^:��7%��ɮ�R��-J���+���E��_����Ֆ׉��^�|�Ħ�h�Z;�{o��8yQzd���g*�]L������4�<���I۲��\K�س��g:(�t�8;9�	cc�9��o�M�Bb�B��!��Q�8r�|�N����-˝����B!:�sJ��	I<%H�EӚ��k�
�B ݮ�g�p�2���@A��diID���ÿ�w�Ϊ��Ff���[�H�����`RL��e�iig>i+�F_^�U��d�>��$T�I��s���>BZaf��X\���g
)O�(�$���0<>���:ƒ����S�/����$yQ՝SZt	J��h��&����d��2�WVuCN 禇1����=9�Y%�IP=*���o�1;����C�Pͻ�2�C�cL�k����-�l`v,����.��ң�r?j���. ��o�<54�8��L�[8a0)?�J�����TD(Vf@ߛ�Wn�0���L7��8[|2gm��C�Hfsx��`{g����J����������$�D���d�D�%�8���&t��yy�f��s?��X�����
��>�-���񵴋`�;:7�`���Rf�B�Bmŀ]P��7C�v�&L^���펒'�-I	2y��ɢ�Y3%�пwHE�e%lDB�$	��i���K��h{e	R�	�����VЧ�)7�De]]W�����V[�$1$���B&�t�E6ՙ�h�r;�|�A��'�vė��v�T��	��� s��?�#�h��#��2<�ثIU �=ܿw[����������TΏ¨�Gˎ��!+i�k�d%MY�����޴�=�նO��Z�2g�oėU+�ܳL_��Y�����*��%-��$�3�Ҿ�~�4���n�ln]�$�!��k!��1!gE)p��53U��OAv4#av#Ú��	%��S�Y3�PFlLѶ*������	�J�ٍ���xє�I���%o�ܥ`��!�J��z[�Mv�$I5F����g�2i����k)7 4�6,�]ܿ���\��h"���W��V�$��4(�c
�,ޱ˥m|���v����;X���uT�G��Ylc��l��O����2hֵ8[G��6����4.
���B�/�
��-��N�F��P��t��Ue��J�%;��R��jcٰ�������3��Д3�x�:Ӵ),�(H~�"MY`f�����l"����{�ʔ�"��������VO����d$N;��Y3��5����⥎���G���S�����D�3-����o��߮����.��U�x�cD��3(�@�H_2�m��ɫ�$��re-�x�OW��+�ʣ�K$�ݔd("�����Q�rl���RL*w�Ј��pR�v%��:�uk,F��rM�j�%A@�T�&[fՆ�r-~�R%A��ú���H����$.ώ�$�Ʉz�p�l<��2�Ѭ.IglV���,��V�s������y0��M���*뫯.`bX�N�.�Y{eW��Nc�ht�ت���-�iPN(�����R��])k�z��q�*٠
�X�SJa��7e�f�'�����M���D�ZǕ��t�,�yK&�n�d��F+%��6���h�]қ7�X5�B\\���<����2j��1(�%�)d�V���34���z����'�'�y��J�E��^�t��3�K�`04"�~�bdɒEf/i�ùT]#�j�k�ꦙU2�cG�=����|��Q,����Z��"��N�΃]<|�L�\By>l�f�'dg3p ��A����VMR�A������J����Maؒd� ������!qG!!�ymi���a ��c���-o�H�0�����\����2��s�7Л�c��8��CqXuy��v�c����2pf��Rȭ$�rf������� Bh^>�G8��ɘKhH�.A�u�c�� �v�`�=�����\,�1P�F"��7Ob�\Ш�P��Q:�	I�d�%��56����<�����<R�-BC����Ğ_V�� Dh{�r���t�pv�B�>[���LJ��#*�'�=�$p�˛xt?"�bV��%�|]�PAB��)8	�����F��T��������r�&w��t�|c.��<�� v]�tQ<� LW�hSx��"�ͣ�$-XhǌG�#g@�竗�0�fB;�������VFR��V-�d,�����ݺ7e%v�¨$<�aM!�v���X'W�����:�o��RR�s�魷�a�����b���Df���~Y|�ȸ�rr���J�s�a#��=-��x��|�~�����[���Q�k�݀��]�eFU��3��>�W�^}����8�~P_+*߳��"�z�tN!?Z�&�Nϕ��$d�~�XRlmH!�de�D��K5Q�V$�O���k��q#��M����v�i�Bz�lN>�c�0IT�n��JQlh	�\o^���/��xG��OM,>~,�g�cC����~~P��'��\�g&��Qs�H:��Bv(}]ӽ��LĬ/��-Do��1���$k��_ywo��5ܼy��m%1�Ue�hH�wX�D��T~k%����!�3�6�ծI tą�mХ`q�2�!�Z�_U��a�@Ѕ��s^��$�Y�?M��q���I��'�� Ѿ��Z&|J.D[���|#L��q3Kli������HD,�sc��&0�m���Z\)�,�.�+��/��3��IMM>��g�isP���t4 �rR�m'�G�wGhʝ�w��߮H R�����f�RC;ڄ�9�)^��וu�8&��D%_r�����}Ѳ��	�g�#eRb�5���g[Ed3E��(��x34/6?,�}B�m�)vN$�°)���)�
�f�5�r;}��鼽�̌��/����9���-��:�+����r�*��nYFނڂk5z���d��E�vuF8���H\�L(����m�$�dG�ݪv�g� UY_�ݖ$��D#���l�GB^"�f��o�$�(���$��4��6���W�����pb��	�Xb�ʕTj���f�����W&���zl�ʖ�+��W���J�Gd��,�c)Y��XǇg�����ϵ�"�{�N�o	6|J�g8��13��>J��e����GO6�ĭ�i�j��5�uV�0�3�e(�bឺ��?SUfϠ�DZul��J�Pc�ئ��,��A�u��ь��i $���If(!��_�*�uc�c�>F�m
Y�b~����;Q$���;$v�s�}�G�*<��|B�ã��cd��ո~��Q�s����R�	a�rgmI-�1Na��y3���wMW~�i��c��U�,[Qk$*�u,��wG␒���G:/��w�U_߯y��k`�j�a
.�38�y���_�l�CɬT�1�	6�� �fq���V&Ǟk�����ohW�Dd���ݳՁ��}vU �}���v�'��Ur��sӈK�hiC�d�T����Kq�9�,�%�?]n/���	m�Q�vng�B�5\�X"����SG��ןO#����0�2s#9�c7����@�ݘ�N*��1�O#?�µ8�U9�1	Z���n��'Jt�zULC%j�L�"D�]��&�/���}��ԙ�	�$�/�i����}5�P����+z1�[�)��ݠ|cItV[.m�L�]&y>���^G�!g z]� �r��V�r�"&�>:�م�&lK�ٯ��UB@�{��C�v	ۑ$2 �H.)�[��cq�a�r֗�!�&�A����FW��t<�j��Ws}�<������w��a9�pQ�u=WK�m�T��� �������Y��䑊�0;�E.���mM��8���� �I��D����(�Q�o�f���Yt5H��TV[C8&g�Evc)VN��
��}u��Y��[J�M�����t��aS���9S%k<��<g4jK��J0G����G�ً#�¯� �5���b%"� 1ic�Ɩ�&!�y~lB`�7���B.�v3zׁ㓲��h$�i�9��eɵ��d B4Ȥ�[j� m\�~��b�����.	Y>��c,=~���I��
H�	�K`n�P���N�p#r�G�3�uՎu�j��	��j۞��=�˜���t~��RW�Z�_�$`_�uS�9K��d�nM~FDx�hD��p�Q��N˳2��08���ЖD!!	?�^��3_|�~9�-n�?������*Ƨ/)[�~q_Z�TFL���K4�Ȁ�*a�a�V�:��d�~LdrJ�~2������G��m97�(J��ɧ���FƆ�N�"QD��j�vW5d��X������$~:�a��.6E����|�������O�������hu�o]Y�g�=VZ�8q�ֱR��ϙ9!3W6 ���O�bЀ�웼���j��pY�|V����9�ik�j�Db!d�ÒL�p�Uev1	dRa�QǰC��r�,G�rQ��Q}j|�Ѫ�t�(�L-I:	;;j6����o�I�B:���ԏ�rO����y��uyT9�l+Խ����ϭ�¿�r~�ƚ54+�@(
g�ʈ|i~D֭�n��f�ݨ6>��n�YQ�ʟN���v��6$�E�j�od�����_X��<�C��]$z�I�NH�-	������br2�|�}����K%�!U?�w��Q���S��!��z!|	�4N��0�s�~e6��x��:��$���<�a�S�(��ٻ�U�����^�HfӒ�(�Z�k�O�ɞ�����Iߧ�n��дt*-�SFU욎�D��+�v��EH����]�(X^g���R�Q��v��R|(񃴃�>I�(�.�{:B�3�aI�$���X����UKl�E-=Y���C�?ߗD��8�$���I���)pv ,����A��S�
׍�V�({�_Q=D{1@}��JN���L	Pة��(���ZFe"%�څ��K�B���}=��A�h6�ϥ��@��G?4J���&p�\A��`l$�:�DTȳm�UB"�A�^C&S�]"�-���c2�P�Y>9A<��J���ċu%Xsmv��>�A��W ��`��T�!2B7:-M�Xl#�(�2��T$���S�1y憼φ�����K�`?x��z��K�.�{R��v��"�S�̽����Lpli����%�4��}�#x��F"�@���[���9:V]}�����%�fA��KYf^�|�A*�2���=`��pw������8�i���3�Fˏ�p��P�2[�&Y���[Wϥv&��r�Fb��2��ݶ��&[�Z��'"��O
e$�0�e����u�[8O���Lfy�e1�ø>��\����(�'2G;γ����@���b`��B�SD��I;�{::M��&��5��i��;��l�k�0dk���p��9���I%�Ѳ�{ ����;�/L��fs����yV��+L,�\>^R�l�fh�&����!�琔EP�Y����
�OgĠzX=%Uhk�� �P!V1�=3��(�&�M���L��gP�t����fz<��Ҹ4��w�t8��z 3{�my��.&FG��%����F� ��	���H,�C!t�Y}�0��qhd�b@����9T�F���`y_�A���;d����� ��_��cD�A��'�%$�1~B�}h;N�t��aT���^��@j����4 �[/�-Z/a��u@�2�r"�7����l�\�>
zpI3͎^8b��l3����Ĉ�A[����Ѧ�����ڲo�j*2��k����2ʘ��$��0͝)��(�I�	�e"���$���`R!���7�Ύ˹K���'G����2Υ6�Ʌ
�u.�"��a�S{J�a��0AI�tR���V� �6�i�O+�}�p���l�R����:��>ER8m���<�x�R�ۄ�r��B��7X�]d3Ȅ�?�F���yP��(��A�ׂ�crM��g��	��f���oȝ)�({#�X�ZѠ=#͸��Q]2H���d��nː/q�C�Lb2�v����H%Rx��uLN�+�<*K|p Al�P��		�w�(ARR�����ێV����_��䨅��:��%�a��;6J0H���蓀i{�D���p�\<�݄P;�z���?��2K$�+�4�L29h-�X��,�ɳ-?�@`O��c5����&T<&�g��h`��1E�ܞ'0�ȷС��Ȉ��q��	!�8g��k�����ems$둠�3�7����k����/�[��ko\ƕ���Y���r��*�\\��P5���
(�}�:8bM	ٯ@�{�>:�GH�ל�}4��k���SE"��odl��J�L�>َ��i�Bώ�)~�.�O�tD��!�)�c�#�ji�.G���Q��cPv�ڨbqyM�-��l��J��8rٓ3�vAD�tF����j���Btދ�l�c��1�0���>]YG�h�H�衊1J%��#IlU���F1ydE���i����8��>���bo���c\�d.��i�=���KZ�5�i7�Y:Ǖ�3x�ٗ"�����n��&n�6�U���,�����B!I���x!�lj�;[Xy|s�J6<�ә���'���$S*�0z�]lo�*/a�l���ߗGcec'	:SY�Ӳ�7�DG�fՆt�V%+W�vB��:�=�u���L�2L`�@�%6E�����0;���"���;\������\SH�5x!G��S����&d��z߻����-�H�&�T;X� J�'��HhQ5�d�wN���)4C5v���k|*�0��l :���=S�"
Alci頋w�y�cq�_<�����u�.H2�BE���g{b��f�!�PlC.�[\B�| �%�N�x�ԖĽSoHBR�Y�g[xޫI�x �`R�Zp"A5��ʞ�S�(I�$s��%�QV�B�Õ�F?����>:,�K7��bE~NK�%?�T���*�6p��E�{f� �N���j��W+�xwP���x��*���'I�!k֒;��Xzt$�`gg�%�mb���D&�s���>�$#-�W�_U~��$��D��k�N�q�^�#�13�Z 2���R�].�`p�&���xׯM��l�+�J,����O�E*�8�Q��$�K+��ܝ(���I�C�u<_[�ر-� �gG%1 n���ދ�����F36�6���_Ըxtzs�b�z��9�I���M��&�y�%�W�"+�4�u�1��~bh.�41v�B� i�ց+�N�JQɆX�`q�-��ӥ�lh!^�t�Aw��@l#E���ւ[ߓJ`?�P`�1<Y��n��ޞ�鲐�L��P1�"�iNNe\׻w�i���;g�\]����~��^u�]��.yG�
��$�o*�kA��K &��TG�<����n6krF�&������q��{|Y�7��my���0Z�$ba#G�I�(A�&����cܑ$=!��Wn�D�v�!��o�S�_���<˨����5�=�ms�\��~��r<�ŝ[�G2��ǃJ�8H�A��ݼ�wάZ�wx��`����>�3�����.�Y֦����۞kЁ�����+L*��s���Z��=i�
f0�����-ܽ� ��!�%�S&9T�;������E<-;MhH��S���lGr��ͧ��Tm����˥#�zi\�v���n����������D.�e����Xp�r	f"� k
�yVd��ۮ`gg_�\ɜ�P��Nׯ��R;�Kr���e�(��P��S7F-����G���蠧�"�plEN�����N�I ?<��'O�sTCX�r����.�����;j 	�Հ��5$2�dҥeNG���yI���I�?����v�L����M�B���]�90{;������OF��Z[�4�����v=�+mgۈ5v�^RGv_}!I���je�a,7���TÍ:Ld�����R/�t�21A�,����lYr�#�$�L˾�1Z��\n�X�K/נ)��R	+��Ԕ �9J�����ذ��sC-;��`t����%vVC���&1�^|�����<]^QM.ή,�n�����D�blBj�:]��=�x�'��v=��A�m����`h^�mO��1B�����ْ������O�x���Ln��}��9��tT��}W�+)ln!&g-�$;%YA�J�aǢ:�F!Uy���M�w�}ҢC��m7q����(�Hփg�* O���uT���G]69Od��QAfԧ3��gq0��&I���3�]n�Ïo�`{���b����c�(�b5����p��=��)���oݞ����;�B~7����a�@�Yw���j"���v<���:d:O�'q*H��ӊ&��a=�����:���P7��D�5/��[o��U�/���d�����$��0%Z8�c�yI"�$����1<9�?�`N�n~r��7;8{�2�~�W��o��͇�zn��ob"n���yW�����k߸�d6��?��'7e�{E|�)i� J��+	�:��bח���$������!�L�y�]�H��tr�c3�$�t֙�Ϥ�mF	�ĩJM̈^0kzj�<���)�ʊ�������ՇL_��6�Ά�yL.�hW����4��m
+�z��O����0}��3���#��"��h��V=�;�1�a-:v��Twq����z���͵e��;x�ݷ���II�:���9�{��{Z �&��!��[7b���[9�[�Kb_�p}��f�E���e}e,\����),�N����ݻ�^�X�7��q��8��'�u/j��}�툝�Q��	�B��2H���J�N]=e���=�ca-��=K�EMP!3��iG��R�o$l�Vio	 ;�����*E���2�<�����jR��1�Q¦kh��KRI�P���1W����߻��=�t�33`�#�C��0c�,��/9{�,I�|�Wp��^W�d�x��Y��΄�s�����>��>��]	ʳ�8}�����Ӳ?qx������^A~H��&��~"I�b����K���X^z��v�{x�ƫ87?��u��S�%�Ҏu�K�z���B�G��h�8��~55!����@@^���MY8,I,tt�� ,gB���+�1&�o�!��;�7elw��D���oy�y.����[xrT��ں~gM��~��*�G4Y ��W"@�1�.�"�,�Wb�S=	S�ӹ{C�`>��yZ؎�������$XՓ���Ϟ�Ca*�GkE|��=K`|����p�V$?s�.]����	yC�����4RIJ9H{���JNcv�,���q��-��5�q~!�D8�Hl�޲ؾ���]{�
��<~����/H��*����#�9Xt�kQ��=
r~�C")9s��(v+���fVqZ���9 �0��x�ф#�i��a��f�H�t�6��(}��F��f����$B���Oa��xD��ItB�Z�M �qi�;��*�������U�^ft]3�e��KR���0�f�z6>X�vcG�ac懒8)5$�jȟ����d�N���Y,j�F��P>'��V���=�����R��o�w�M�ɚ��=��*d}e�l)����<r����G�HKr��B9#ٌB����O�'I�ĭ��'�]�4�w�!]K�n�L�5�`�,mP��`��e�c�˔N��%�Jw��|��|o� r&���?_��K� ��������L�=%�IeF��<F�����1e�cr{X,I�U�a�B:�D�R�3�Fi��=]\��h<�m�F���Q)�+E.�?��S>�cO;7,�ᰡ��s*����r�]Ӏ1.�^*�G\%�c�4�b����P4���=<\ڔ����r�#վ;�9���A������1�w��ƍƣ����@�kO����A>;�G���n��@I��'����|���F�Z�*,Ӵ�yx�:N�|�
�rN!��PQC�d�lo��s��d9m�����8�_�.���/�o`{iS155"��DC����$�U���$�Q	��f��RS����DH���A�hc�9�\Ғ���qI��xYx�h�8{�u�H$'����j��0�+4쐒��S7B���ծ��p���vF�B�Z]�;�8���w��� ��T�8����\Z��ۧs���djT�a�{��<�Z��������C�ma���@�z IUF�Y��S�}h<��4���%��9� �4�V� �ս�B���[�s��#���I�����Ve?c8{v��(�W�H��f��j[H�]��XF���F�ݒ�#�L2�]ò8��2�Z���ڐ�$A}]���_>9��Ci���H�44��$��d �@�%4����e�H��
(��J{����,,NT��ӌ��g�B��v랬<W���aq�rv*���Ki��RW���x�#�pB#��J����窞�~� �/(A )�	��HPĮԑؙ���;� ��I-m�.�O��̇R�ۆh�		�j�*pM;ܯD$�������*)2��̼R����痸��2�$>��ocz���~�?��_��w��?��W1;=��[k�4�N2��zx��� >��o��G�x�}��w����yl<{$�P�"q0}f�h7�=Ư?����-����.&&��o+��[]��D�mB�8������4�`1��?Q@��F�s+����Bx<��aI��7�6�����;͵j�8�i����]��Gm�-�B�zzC�ԕ	e5��mC����&���|��=�J����,�,��z��p��y��4�<����*�
EI܁T+脋��f%��D�c�����;v������nH`n�/����V�����x��nyK�Q5I�'Y�ksȧB�η�����bm}?�������#�y�I�V�ʢ4��-��(�ꕳ� �G?�����������~�%���}N#�R�*[� r�@�E�^�/����gydbdL@r.I�b;m��:�2����G�&��+���{�͸��#W0,A8Y_@�`��O_>�~�m/��bK�_�����f�Mp�V� Y\�s^R��o?|��g��&=9��=/w�~�h�7;H��ꩩn�O�}�}�ե�F��~�svf�.�`yyK�wX<��H_wA�ܹs�g$Y��1��>�-���,������8)r��$NZ���-��^��o��>\�'�U�/,$��[b�/`S����s�<�|�ƫׯ¹<���,+T0H(7G=����Nw��P�����G�A�d9�!�EU�a?�_ӱ�FE��Bv$/>2��D�a�{n��	-o�k U��+Lب(%�=���&�b���7�q�{n��r��7��NL��*g�����r.fV�	�a~n�v=^Xx�O�S��(�z�~����y�v��?/��+�݇kX�|����M��Z��{x��,A�0.^�!��I�r���u����s��4������q��m��ØK��?�Ն���S�hX��l!���YX|�㓣��U��J��D0�r0����HR��N����&댻c��
U�xO��E2�ܙ1-��e�E[�"MV��A�����2q���^r�zk�3O��s���QXdS�gJG]��i�;�`�M�Tۊ(�����'J�E}��!���i��q��6#/����C����79+�������aQ!󔲹~uJIW�/a8���bO�ZJ �1�0�y��ţ&�����J�195�ǫE��EEt�M���_b��w�ۛbCrV(M���ơ�.�y��~M���:�a�%�	;��s�պ]3���a>�\,�6����"��ј��6U��^��g�c��8�h����y;Ǉe-�������]����|��?����nޖ��Y3O�;�ˉA�СͿ��o���p��9q��p}�*�ܖ��Z
p�ͦ�M����*ƨ�Z�p�4
��'�ʆ�W"�$qY��,?�A�`0��*��Q�`��Ą�����!ta��g�pL�Q�
�;��b�ӒF"b�dtđIZ�D�uX�$��]I���LuC�p6���&�<���AW�����Z��6<!6$�9#���#�>��͠7��*��H���V��͆�N�cA%80�`_1�]�k�V��e�i��u���[��s��߮��ۦ�73���o_���1�E<\��p.���Y��ܸ2XY�byu�~��2Y�$�*dCx����:>ْDQ�W�0��΍�$g��O>A�,��p���I�6�GKےT�����c��8N�)=|t��d)%���<�V`(pJ'H�cΪ��q%,a���5��TJ^C�����u�UYGŰ���Pb�����^�3s_�k��������>��S���\���t���\E�	5��_C~�`����9W�ix3��No��L@�zI�&���䐁
�L���xe_{��\�"�6�c3;�û�ސ৅ziHū,���*+���o|�]T�,=���־2�͈Q<37&w��Ͼ����1������oJ��ժ��'O�)�q����w���Ïn�j���J.��\��x��4��[�*<*�4$��jzY�tHJo�bt�z=��&Ӥ�ϊ���V�H�)F�0�g�h��̈e��^b��Ա"3�'
ET_,󣸷���=���GE�&O�NG�Dzތ�I
mVO9wI�c<�dǐ�Dc1��7��V�
�e)E�Ŗ��r�6�tGJ�wO�DGl����܅	�.>���ߥ�UP[��4t�dZ��H���|]ٿ����=���?���D����Ƶ��bB����J����?x#g>����\�iA�۱�ȼ�ʶ�r����)"y�H��ɧw�����#;�C4S���$�A��ވ��{�^R�q2�P���b��A�B�}&��D_9�L����kV���s�OZ!<�����?3+�9�+�/�)�H��'�|8<�*��0J&�sN璼.6�ɓ(���8���xS�좎���ɑy�?��oG��h��1K��}��n(L���70V�q��!67v�~�w���e%�ɉm�bo[޷�r	���3�S�W���g?��ϰ�0�⽰��c����=��]9ki|��+�G�%>��K	FǑ�Nk�ԜdG�]o�S��슉wG~=Y;�I��5���%�JR(�jT�cfbT)�٭���Ξ�;���{��h[ф��0A�uː)�O���n�釭q� $XH�APȧܭ�������R���W�����Ut�.7$�g�Z5��So���<M����=ԑ�<��G�h��Ԯ7Da�k���/��V΀��}I�122"��+Jh����������
�gg�RA���M���PT���]�}���O>FP������ڦ�9_���V�̑�&�Jb���O��E�#�IB��`먮]yI�Z=ex�j���qU�ཱུ}7���"0�!�"B�Y �_#D5��9#gP��Xү>�O��	�I�'��ӱ����)IL�Q�E�\�$�+���Zőχ�.p�9+�|D�)T=�Ƣ����K� ��mX�tb��$�� ���������&�4���*\�r^�nUe�tr}��rw�L�0,��Ɏ�,�0�����:�ǖ��&�\R�}m���c�v�*r�6�?� �2pk���t%q���O�153�o}�Ēed�Q	�K�~��SE]�
�����tΠ�$x��)���L�-I��E|��;#�3�� �5Y O|i%�#\�q2-%M���Lh\ly\x!o���c�@z�a1&��Z�u���������,�ؙa����M����=|r��M�'~i�Z�<!4y�m��,C�����jS�h0�m9c��qy����M<^z���W_�d<�O>{����p�2f����8��?Q6ZN�e��\��s���*�7�q~a7.O�rT��ё�ƌ��� �kǒ���vp��EL�<گ*�+��sǲ�m��,n�Cq[;��t/Sr_u�>`&,T?כ��8IPadX���-��0������g>t��ꅌb�c����k(�ڃ�WŰP0��R����j���DHE"x�]����7dc>��e��AG�ZZ��}����g&� Y�-Nf����_��W���,��QR�_~��$b��:9:�ׯ�����_��Q���7��c���>Z��QQ.�_���9LMfp��<{������r�r#>����%���˞��z�
JB�Of�rWP��aЕ�ڊ��]�d#Z-G�dߊ�S�C$�K��{$1<�0]�q!�8q��3x���i��4����g�An�$�+�9	:�����+ �k�/.��A;�~3�e�&��цw^��]���]<����j`�6T��|S*��+p�������GؐKu��eI.�em��ѯ����p���*���8 vӘ�f�4��w�tΥ!�L>5�kWƱ�l	�K��\.��y5`##����E,=\�`id,���^���_~)9��슲�Џ���r`��������������7��4�6�����bH�p0�B6�*��2��%���[j;�F�h���"�+g��O6S�\�d:��'1��<@����Ȣ��j������EmI<8��
�m�^go��0�71���D�)����	����W��7��p��O�[l��������^E�Q�ǿ]�P&��fQ�5�����LH��K�(�2��/�{�<��oJ2��̌�k�&qx<�[�7�9J�LNJ"g������VW�%�	⃯�'�dO%pJ��NIP[���2�{���J좒�jq	n��.���:���?��NS�����ҡ��)l�L5�sJ����&�һ�x�G�P��v%�bb�c��>���Tr%I�`�x�PѶ١�Zb4���G�}T�KLB�T,z F��D�I��oYS&�����Ri9?iٓ��e	8�\���'%�B��Y�����$���8�3s�7,���Yo�h�CX|P�_���şT�_� ����^;sn=z��iã3H�}8X>��.�|�_�_�����Iď>�{,^#�;�W�����Z���a0�w���b��M�!�,pa~����������#��*�J��S!_��JFM�����BU��3�ѻ���H��y�ѡ�+��k�p��m�J�99���~�����<{I	��a�Voյ(�:���y>D����:ދ��0�Y2�bO=-6�~X,�>v��j'�]o�����g���%I����+8�y�:���b�\LL��^w�ޑ}_�3�O���&������������X��KSyk[�8ܽ�����_�w����\��rO����T������-�f��t���9�=?�ݭ)�d�� "+�yLIPSFT�Q�����ak���6��l��.!G�O�v��s=�� ���'����GZ���x		�j�R�S�19�6>����o��{_���d;��`��yZx1��zs����.N�+\�c�u���Ɍ�Q�vJ{ �6i��zF&'���H�DT�&�TO�"�D�q�~f!��w7q���bk�÷��*��CZ�L�,�vaX�#�2Ŗ�ڸ��m��u�v�,��6�0!A��n���k�
���nT��l��?�l�ͦ�ŕl��c)�d���1�CI��QeӜH�q&�@6:�~�G���;��s���/ۋ/��G�ml/�`�&�-�a+��˛��T�ի�$�͊=n*���Ԓ}�tKl���'�:b41��=ǋV�S$��AY�K�5!!J��OV��ߩM�*�?����&M #������ 'k���c�l����� TO^�v|"w���!	��)�r�'paaV;�����7�O*��� ��vQ��cww��(S�����ĮVm�-GP���L�/���aV	I���JETzM�[HG��I8�e�-A�('v�%CI#����6#K�O@� �̝��V�Z�;3�Ɠ���2��_d�,KB�GBl���g�f��F���g�X�ɋ���� e���2�Uo�D	%�$�����p��ۘ� @������.�w������)���J��m��J�����q{�;������3r�]�M�I�Ӓx&��6�
 �[+�%�*j��3�kOPktu���i2f\MX<k��to#qD����w$v
#��+�w�I��󒴸�?
u055���$cg�?�u���~*
�fd
��d��A�yEe�)��� ;�nGy}��ޔN�����Nbz<���
�%�ow�>+�����?���g(�{}#��_�>_|����EDĘ�;{V�H �Y���'�������`�IB@W�]E���x�d�x�:���KO�ӏJ�Ʒ��k�g$)�^fBx9	,�bxD|�yT�>�����]?���/�L`
0��
4:�]%���XG�g#��+�݀j;Qhו�&��0���1::����Br�"��!M�Z�������~a�i��m�djX�zD%0�L
�^����8��c[�����a11ʎ?�G+U��D'�{�:z��b�ɠD2�r��A�i��\S1�yxZt��B�a����i�Q6
I���͛����aA��?���\!r��2#	UJ	a,��g�b{�@�t�sIqBw��f<�˗�.�99Ѭ�5���<���o���(�S�+I��\�rCEܣ���+�>�eF�-%������b�q����lL|J��5���^�{��0'HE�zuì�M�U���2����Ջ�e{�k�/�YPK���Ⱦs8�m�v��J�V~��̰��yI B�W'5��T��u<��t�I��b�P��#�y���Ի
gh9���=f�T���m#�t��4Z�@:!��/�%�x��ܯs瑊���o��?�1.���+��%H_���e
��MK�CI�	�z�u��X�/�W�����_���4�ݽ�Uq\+O|�7/�܅i�����o�+AlZ#�X4j�-ҡI�L6�`"!I@�X�n}��|���XF�3�3*�$�l�
�B�.�ü$�\V�3�ܻ���Ώfx��2J��j��9;&@�|���p���αm`N�B7j=n+4g~a��D�VF��H� �g�ڒ`nу��U!�H�,���TL籫b�L ������u�ba�Qt�4&˯��YW�¨���M�����H�����=~$�ᬼ'W��]��0�����+x����	53���
�g�$a�9�r�����Z<#��Zw��?��g��ht��ه{���&G�x[�wő���� �Pe$}�%k��E�#�P�����[���q��rq$�~��d0;9�ᡸvwR,M	�Ͱ4�j�U%�X\q�x��}3�����0[�����ޚ⧭�S���%��������D8���.�_���>��S��=�uEkH�Y��뼱�>}b�߭VW�K �|���)U��V�QGp^�ek����;�����)	WS�����	��A���� .\��ӧGx����r	����@ҏ??TvL��Ųc���"��S��Mc{���-⒈���<����ޑ�1$�&��!v�?��׊�}��_��˛��)�k(V�|:�rP)�k5�!;�G��)<�T�,�E��d��fŶfpav�_�?$������!�Hxѱ͆����հ"�)WX��RĞ�;y���Z���8Dd�V�J�S5Y����u�|���!>��~��ǒxM!�$SJ@c+��U([���ο�U3	�v�>��+�Y�[���5��Tz2svY��$��a��u\:Qgχ�I�Ofq��,v�;���/�cu�X�c���{x��Zޕ �#��#��V�a]΍�����$?�}�	@�x�Η{x��P����-T�x�t[u9O	&3HF�د��Ƒ
EǒÒ�P�!"�bO���ZUɖb	�����SRW�v܄%w3*��0=�|"l������y�hЧ��<���萞HL;�/�E� ʬ0�P�Uk&��#��fÀ�sI�\ �luyj��.Pz���ۘo]���������ϡm����ǘ���8���O��u����&�H��1@X�MD����Ή٘����=	���01!wh'���%�EYv�6֟Ip���ׯʡm�/����fg]-���<S.���eI�b�I:���)6���$}Ń-�Ƕju�
q�s�T2-���sl�QeZ�&waxD|���|]>�>�z�di�R�D9T@��!�*�<����>��/	p��.;�Z�,RpnT	:�Ic��\E3p&�>�&7,	�D�^ʋ���+���h%��||�H�:�
d�B�<��wz�4�=�����jxCӮE7E^yPmE��}J��rF�����jx�1���X�\�xU�S�se%���sWն���cα}�W䮞;K��U��鰹Y��3���E�'���>���9����$�`��r�U������瑕)(����Vg�\�����$_�w4��H45^@*RΏ�$�II����L�iC!K�����\?`d5�%�$��w@�|�����f��Q[�wgg�j���gU�Gw�J���Ϋ�"z�[�_�������{A C6�7���IyjVy*�k���_>�ald�3i�y������hJ -�JjX�.!A�l��'�$a8��~�8��VB(�~n>����q\;Ą�Ԛ���M��֫������^��:K�h����͠��ݗ����+	!0���aedhD�C>G����qqzB�]��IJC�!8l��b��ړ��P��iI�b �����O�����+SY�:1.[���b(���s3hT���"7���-!�S��6̕�\T�g��P�E���A�6ا�
/�6}J�%|�l��]]�'R<�
T�T���\����΍c��)�nU����!�������nX�L`��kX^]��~�k��7��H.dh�+F�b�dʇ/no���}�ܸ���1b~��c�L�j]W+m���Ⱥ\.2[iatk���-��������K ��=�$��`Z���$�>IB����P9�C? ��]�c7@�r��{�Z�&�ݫv��HF�F?��gH�㈼��$�6w���w1��C��{B6��Ԣ�*7��$W�}_B8��=v�ӽ4���GM9�2�FK���z�)�� Ǹ2>]ZR�ː�ခ�p&D���'������|�կ�O��=IH�>��\�v;r�e3� N�����8����W�������fI���G�h�
!I$�
=�9Vz�������V���_�U�;R�_�Ŵ$�R������f��k�煻��U߫������ݪ�f�Z�t=X�!�pt.�]͛�`K�w&�F>8���u	�wp��5��} y����>��4�e�c�L
��3��Sv@�#�	ڄ��|��v��s�W�dp��y�����}	X�I!3���F?���`m�3箈��b����>�y�
���񿓤�9n��T�H	:)���I����������?�=��|��/q^�^A����8�0�F���$�r�T�F\[ۈ����������I�$`��K��\���ݾR�����!����fS���}	Z?]��$��OE
Ow��q��f�v�bpAL�s��m�y����c���<�y������z�������W12�Gw��=�#	e�~�T= ;1��|��Ȯ m���cG�ޔ �*I�#�嘥	�I�;$P�~��&~"k�_[�,��Ϸ��<ľX򱡈{���H�M�k	���uW��|��������xQ�iW��yIh��I�A*7�ՍuL�i���ه��u�W^S����
�(lQR���+)�'�U����AD�%���rfz�_���SH�-�J:A�x�]�I٣���2�T$Q�a��D��-�9���/6��m�p��n��]�@��'���d�݉X2��Z��ur��W�o������⥳��sh��^���5RR���<�_cM�KU�3D��m�a ��[���[]��Ƣ��V2�׋�[{��l �Ώ�O��uMh%�ǃ�u��=wM"���b�����ؾZ�����'X��Ɵ}��(��㗿��T�/_ã�5이�^���,�g���/�൷���ϟac����GK�N�^�St})ճ�7%���U�=	jͧE�z-��X����ȧć��U����5�T�o�J�߬��Ֆ�m�k<?8�^���mr>��v'�#�S���Gi
1
u̞*LMY���cڝ���k����`G���#�cC�b�#�h2��3�NN���`�x��K�H��6�BeW����~O��:*��"�-D�I����C7%a�=��d�����T6��m��?PkX|�ۭ��7���������w$I�TY �bxT��VtH,ƌ�X	;e
��{x�ɾa;f!��^|�ZP��ݘ�+�,Ν��KrK4����|C�zG������S�L��U�D�Jr��ʝ�ć_!�_g�!c�t��"�\S`��Dg��?�������;7�Էs��6lH 	��h��e�d�e�Tv��\e�?���R�lY��-� Lj���b���������nߜ��s��{{�EuU������x�s�-]c
W�{(۱���,��w���'�%����y6O���h8rR[�u�����{�̴�&4�����O&	�����r�Wx����Gǌ?�p���8���y� ��2�k/c�lw�.1��"_`.�5OG�������1z�:�Uʘ�Θ�yk�4p�M��;��B�g/��q����g����I�9�^�F�}00y�m<gK���Z��ڱ��h8���6)��"x�yq�G��>l�`��NJ���`5����`��x6J�_�p�� ������Q3I��t�Ìɚ�{UP�T1��7F����j��1N.�d����������:�q� ��CU��^ZP�.�O��{C������E#���hzZ�a�ƻ����Yǟ�������;F��v�2F�w5�ܪ��VsB��t���|>x0��i�o>�/^�O�&��n�R� ^G��l<س*��4���4���Q~2�dd�٩�9�l&e�G�;ҝ��#�aͱ�,�����>�"t�5L*��(`�[�u1���wn�~D�4�h�5;���6��[�(�:I��͏�)����4�T�C��f��E�7�f��P�幁1���o�u�K�Z�KeT����5�&���K����[&v���|W_8��=����4��x�-lm?�g_�x!��ҕ�y���#|����U���G6X]����?����g�
2�����~l�� �@ʁ�C��Ҫr�B�`Ա
L�Nk��U���II8h�X�h��̋�E0�AW� x�0�o���Q��`6a��n�hz��e�M�����4��cX9{)��3!3Z�������穀3��L����+��%�9�眈��pQ�_����dNc�{o"9�#�L������_�����9<ݮ۝�������zт�ͧ[Q�&2�=]?��������#Ԏ_42���5<~��3yO�rtH\�l��F,Z�����.^�S�}�{�>�vĊ5m�tA	��2P��x~7��18�y���o�$/������M�p4h�Ym�:g#$
����DC?����\��5o`��2��d�-�H���]Qg_	"��W_B�0�3&����Sx����B�)�,LX&Up���
��P��b2�������99A-#�ӊ�XFE��:�����m��)6wV�N���7���M��ԝ����'6�[j��.�8�U�C^�
�r��uuae/��kh��5?��+/"wc�ܼgso3i\[�b�I�XI���;o-0��c�Ax���?��OQi7��
�ZoGtl��i�|��k���W/dLd\p���D2�s	�KG���pT��ȿvv��d��&�`�!A��f���O[?	,�Ӧ�蹹�ङ/ˍ��R�q�k&X'�|v�d��L��>v��㰡NڣF���ACJh�=ϟ�}�z΂ڧ��iW~��R+��
~���)̎c�d0!R���G8�9o�	f��j��x�^��#VJ�O�r���t�JJ��|�׮�������L$V��E&$-Իm��w��?��'L���O�L�cPS���/M�ynF�U��~��)������;���h>PP�.����٪H��>>7�ճQ��ѭ1Y�5�?m�&�9�"YD�#���Ul�����9+�ÎI2%2SV�Ѽ~��OC>�������t��T*S�4����b�u���gȦc���Fb�v�|����3���T�I��γ�N���k�TwK�6W��������©L���\�q0��`�9&=u]b1���	n�\����V����hO�C,`��	>�b�%x�����|�|��υ�(���f�����O���/��{'���d;����"Þi4��X[[��W�p��Ǚ�9��z��h�IK�~0l���drb�ٔ�j~�����'�H�0�O�DC�ȭ�7&��6�Ck��lz�>�o>�3�?�6�a,����Ys�c�[���7v!��,Wp3MǠ�l���c���G8���ʍ�m�{� ����o�Q��H�NE�c&؛%��K��8������Q��?ɖ���Oɜ����3hWG���&n�nX�b�g��t��k�Tq넿0"���H��م,�)���;��������2�!�z�<��G�����9e&}x7������9ƹcO��	��#&X�/Q�e�w5O?t!Y�v)a(䒘����7���,�1ͫZgbإ/8)հ�D�t�����B$�E��p�� W�+�bHGH�:�I�H�Z�<�:3�o����O��0�h5y6*��z�&��l!芼f/��L^"h3�����BH��N��#DQ�'��6��x�k�2ńpސ<��ν����9�����XE��1�>��f\���WWi�Mª\92��H\�C�laUe���0�+/ I��N�  O�ٷy�LB���#Ǒ,Wg`�Jz��Ӿ)=c�b9�t6��4S����m��k3���NDb6����^�K� r�*����H�ր:mrM�Y����%�"]�%M��#l���y?�z��\����Ύ�޳���_��٥N���;�������:�r��熫%��wc���{�`6�~�������͹�ŕ5��o��N㳛�VŊ$2�$|q�+���"W��!��/�^����Eܿ~��>4�J��ܸ�5/�
��x�d�����%:� ���?=�ä1 ����	¦%���GU<F&�L��ñd3;9nn�Ið�.�`���m�։�o�װ[�aa��ĩ�y;e�F�o��鑇�VrUK��t�}:hk�y��D��Ɠ�C:�$ʵ*:� ��y�� Ř��)��x�W�'�����Jw����J؀p�f�$���A�����{�ob���իWp��2mMG-<���F4�W_���s|��>�w>0�Ey̤"h�_���3͹H�̓��[F�N|a~�� ?��Wx��+x������h�3L�OL{�ӇD�k�l81�O|p����k�	Cj1���ՕY΂?eyYy�<�Qe��^5�2�0�������5�w8�����sa88����͐)���κ�j�{R���1]�7�}�r�޼�������ū���+��r���GƮ ܾQ�nc����c�m &�_#����7��+W���:9��`��KLW��m=�<�7>�
J�^}�u&�Q|q��G7lV#�*08�'?�o�r������+��?2��˗q��}c-N/��x��O~��{�����'���_O�mT��P�'�	��YI&:fG,�b��?�;8��ǥ�&��2n�}�V՚A��(J|�Qcg��`�zO��a�<��Q��Ъ���3gA_�X�$�1�۠�����na�w27u7�����Z������������t-h5Ӏ�|2 ��xnNiґ���[ӒCn�s�'�t�[��XR�9&s���m�8���*�C6���c�):t�&��a��[����;g�y����?�������+ظ��������έ�_��O��O�[ﯡr��?���'��@����������r\��#�}y!m���P�G��p��}��Z��HeCHœ������>��Q�w6��������br
+�_Yf��#&?M>�γ�C�����Y@�\#�,��������6�,"�Y��5��'�!w+o	��_9�!�^�����L�3��M���j7&��
���4Ϸ4Dp�5�Wu3��a��ЬU��?����L�2����B�I���C���D��gs�3��U̯��g��?���c����������g���˿���g��������g��G�����❷߶���ƆϬ�����>6NA��>TTS7]0tu��'-���4��Q�p-�0�i�`�"hsKܻ�m�=�u&��z�l���4.];ϳ5�/�>��IIZ*�H�́�����|N��͗��Dv���I���Q)c
������+�}��Y�cYC��Y\��~G>0r3���K����~�W�Ďi�i&>���	��&FP|JG{�㽟 �i|�gKv=f]�M&�GUڿB��Yt����)�o���!�����m��{y���ڧx���������~���7߸�T2��?�W_���K���&����ի��	��m&���,<�[���y4���,P�>��8'���9�]�zm�Ǳ�.u5���|U���J[G�6��'�(������'B�� �K����%�Ɠ�w���P�t�%_�.��{��|ZC��Ե��A`�,FՕb@>X���"�X�ur�'0��ώ��>������t3U~��
m>��'2�i����Ǉ�c-��e�r���b>��L֪��/���E3�B��s)�h��/$T��&��RK5?��[�(��������1�<�3fm��.[���l�2���+"��L���76�X�ٷ&Qxu��7V[���/���L#!�L�?�E�Z2���X9r���x�|�-����+P�01%0�כL KՈ���x�ǻ�p���R�f�G�+�R����$ƇO�4�Mp��U怊�����:�?a��X/I[ޡ�:A��FG���}��:j�������"Ξ��9�z��s�W��<��{���o\Ý;{�S�5��(�Ъ0qb���+��Ƽ��W���&G��I���Z6Ea0α%�K39��'O�Ju�<g]bŦ�W=ھR�w�Dc|�f�Д]u��){�!�d��z�~<�V��_� bDe���H���Ov+��Q�o<<n�\n!1�?��M�ճl�]�_ٖ�i\s�&*���x;�����T�|�܋��/���͇L���z��&NCp�O��Ǎ��Oc� ��˗���I|ׯ��Pj�2�΅*>[�pa<~�����7�2n���t������r����D�*ʸ'�И���T*��.\��\���S9�z|/�[����X*� ?è	5WiHw�����P�3�
���/�Q�����@�v�$���a[<�G�.��^���?��/�8����,�����lnf�uN������b�s96�k�$�9H.m�ƿ��er�>��y9����*p�}AC?��Kx:���*�&�y�gּ�׷�+����[L�-XR��l����Y�s!^���#3y&�C,2�S�J#��+���.����t\ް���Ѿu>���-�Lڂ��%K����!K���
ⵗW�X�6ܯq��H\�ܧ(��8j��!�
�f�t��ܥ��
|p�\�������l�i��Z3����i��[�����ĕ)�x��.������;x��א/�pkg���K%����D��Bsr��0�H ��`��鉡�L.��[(�H0(:دࣟ�C畳9g�l�����:<�>�����}� �e��r���e�1S���R�˫:.�C+���7���ocg�d3�o�y��s_��sX��+�8�u����]���_���>}N�R�v�к/Ϣ�8�M{��^��P�s�t#Lt�,r�2QA124�Q��9`�z((*���!>ޡ3.|T�Ґ����|�05 Gn�g�C��������7������;�G%f�:��rSt�c�HTE����a_�̘�$�+v�n��:��Ng���Ds0"�2����D�v&{gWg���2�}���ٔ�zbV�	��:�Y.b��r�?��dPIr{]ڵ��_�m�Y^C,8���gQ`Pb�Q-u�O����~�3q��믣A��λ��L�ai�AP	�"�7�7{N��b`�gSS�X�OL���O]���3\%ڔ;�����A�;DKȏЀ�7���)\]:���3�=���]O>a�����}�j���;>�Hb��J5�g��)��6ka����#�$�&�"6�Z*�����
E��Q�`Y��_����S�#7�O�a�O�O���lZυ�ֱ���x���禱�����t2f�wQ��4�*8�`����<~���j����=���������9���/���cs�ۛ�x�L���>N���7��_¯��6VW�1���gn H�����J�Hî��2B:�ĈwoܗT�'�Q�w8�@��)(ڍ[��xk��eZ-t��3L gp~�VV�L	���apb��o���5��32��C�X+��y��O�ݓx�9� /���3 �_ͮժ|�}nB�H��KEZu��j��Dw�LN����9��DP!�)� �=т��غ*A����dyz��D�	|�L��&�Ȏ��L�Bx�t���v�,x��I.�6~���3F�����ρ��Q���눉�9	�V�g��Dl>W2A��- ��1�1�y�j<{FE/Ē!�`Q�/��G��T�f���b@�e`[n�yҝ}�#�U>�H8��8��������_	��6�9�:3�N��!���)�.�I?!n	v�Ii��e\ѣ�#�]D�>�������̢�%5[>rR'"�ss�#�ן�����������6��o�r�Y'����].�	��$�DF6��������w��u��6�e�bߓR������*_�|���������"���a���3G�Lhe&��߼�����S�ncs{�tӌs�C�2v#<cύ7�;��g>b��kD�ΘIl��r�\5�wȘJpu�^��?�r9�-."͵�e �Hǌ>��z�LL=�qGp�I�>hp|�ކ�:-j�Ψ�*�4��˔��)��fS3�����߬�X%�`��g��u��-��P���3��;O�����m2�)a{��N@(���%#�6-1��-�H�b
%���s(N'�ˏ��ݯ�~�7p�w���]�FW.���ͧ��==�7f܃�=�l?�=�1���R�����}k�\7З��G�(Q���_"���#�@�~���yJu:�je�KUTy/*�&c���܉�`:[� �i��K3�X�����5E��X�I脭��@�?Vb���8>'*�q��\�g}l�v���̘��>��8M�%t�=�fvL�����L'���cF=el���a�F��G��B�3��$h��!w�V33��|`���x�5��AR^z�"fx�47!V�W^~�Wgq�	D���.,�������Y�����q�K0��{�E�Mj#Og��峸����AU�PZ��錉�*0�����xJC�utb~�R�QCt�}�f� f���ѵ�[Ȍ��+�uV�	#�+p#J����0W@��~����S���Ea9�ĩŠI�����`֦�&}���ap��U�m
8�}�zfLx>��ؚ�G&c,j1L�����6j|�l:�J�j��������I\"ic�4�:�ٹ9�ڷ����-|�3i?�>x��c�����ߠc��~�caa�s/;tB7>�ª a�~��:.^�����u{��8�r�D"i�0����H��4��| �18A���$p��6��4<�=�z�A��A�vdc"�)�h��|���82�I3�u�lq�@՝�c���U1�b�\�����-bj!��,��ǘ��b�[�����?CA� 
b<
�����E�5d|�\��3��<����̢^>���c�{L��dP ����\̍7��,�H0$,}ۜ����0Io�N���EÙ�������?��G����Kx����O���k���W.�T����	j\�j�e��&�w����\N8��p�L�����	T�ViYs��D�8�G�^��L���ΧZ`c�	�6�8ium�'û^(fi'��F�O���{<���1��}
r�GVU6����^�w�����%�ť�8nz��O��yr�+�s�VmvD�Nd�$&|�B�O��>�&L3i��ؓ�T2��[��7���a�uv�F�ߢ#+����\W����T��� �"?t)j���sξ��O~�}�u������◿����<�,ײ��7���G$��/~y��^er��Y�|���̔Q�4���Ve/0In	o�s���>I��5J��I���9ڞJ�@l���;�-w��'�)L�ʹ,/d�F1�L`:Y@2�����d�=G5!p��δ�&�� |⃉.g��Vdw��s�ڽ�����#���o�Q� �x6s*��3�u�]dwO\-&�̠�����1����^gI��ńp�����t�<��^U�1�w ��z��<3���U��?^�j�7��:�|p����g�ʚpw{-����Y����S|��Wpau''e������ב�����N��f��J�g�k�AN�o����*��j�2Fh�0�Sop��}�o�1)�ݝ�Ǖ+�pve����(R���R���V�ȟ$K�Z�<�� }'5��;A+,L�0=���O��z�@81�S�H[���+h>g`_�ֹQo�,N�s4힟�d4�$
&��I�ᴋ�'��G32b)��}��~.�o���ΐ~c�t!dcFP�s��Yc%2p��Ԍ�8���瓇��za����]Q<}�d����`C�~���6���Kז����-)�Fr���]<�x��U�Ǧ����Jզ��փ����Q@�aul��b�#6�%馟r��4�Xot��=WdⲰ�i&��|q~��x��~b�
bx��l�>D�f��H��Bm��*6�X�6Ս�\��(zp;�c�1&j4V�2�-"�DȞA�f�ݛ4�N�͹�I|t\��5�G���,V�E$K�DF4���$(_���f�|Ҫ��GGpJ��f/��k	w��}�ְq����F���XZZB2;E��Ũs�x8�~������972"$�Ɠ={o)��AФ��|O���%!֝������F�"�l--���JcPLh���[\�L!��hR^��e����z*fQ3�:����[u0[�2��I�*�D��1����;��#��L��!�G�CE5&��x6�k���%-q���e,�����5@������i�R�5��J8�|Q�M��l\"�}�ب�sӞ��3%қ��)Ɯ�l�2Ϙs��mP�}v�������"��u\d���W�������%e�i^���'��Սcitf��Bc!'�8n3G:����\b~�@�y�H.s�F&���P̡���p�~���I�'-'g;d�u"QG�#%<k�C�I�ܥ�$I�`�?�����i,j-����0h(���X�&�*#1��B��R��d/�E��S�Ѷ��S��S�z'������~��Dk��^2m��~�S��η�������u^�.]�hǷ���Ýu_:����G(d�(LM��೤X�eg10�A��MX�Ө1K�����B����x��}�б���t�������7�3����lq�L�N������kؑ��%��t�?ԩ\*µ	��=nb���}8)m�n?<Ɠ��u;��UB��o3!��
%r���0�J�_���9ܵ��^��i��nq;
�F]c/��)�y�(�S�Me����&��9j�)��6��8d�.�[����o�\�cqqdT�1X���� qT�p2ɔ]8u���W��,0�ߺ��\~�#H�������R�9SiE��`�}�_��ۍ�۬#�˛�iT�8)7Q>�2�9���R��/A ���`~m	�.���#|yw���X�s"��;�g}��1�����u�u��̪�:���;�d2��3M���;1���9��-{P�	|9�W���i���g'���Ip��Ub=�ܬ��1�t&g�M�\1A?��	`��>V0�C��萛��md蜅��E�,EU)�d
��Lzx��k4,װ0?�d��$b�J��2�������5���:y����C��(ª��C	)m�y��F�����q$i�٩)L�dqaigVd8Ӹy����OP.�H�lF=䒬�9�l�,<���Y�;c��ݝm�t'
��=��m��]��9�&�1�:���ר"9a�����9���3�O��*h�{�W�&s���+@��"�͸��4:�{_���G���0D2��D$�Po�Q팹/�ni�ܺ����C��.�%X}��)&�o��*^x�]�/_ƃ��6�\���h�CL��pt�cO�������/��16�>�r >`;h�.�����*���6���
�R��hc���������l��m�ʞg�@�gP��s�! �ұ���hҥ�?���H��ƩȐ��M/����eM�7hVUڮ�A�l�^����j�$�������+�y>�;:�p,�0b��%1�D�x�6/k�a��	mg$���?��m�M#�PATA�H��"D����_��♕3��������gn� �b#௼������ŗ��ޱ�x���`s7?��X]*�����[��u,�]���E<=h����q��`td4�"����r���Ub���yhh���#��tSk��]���"V�ӘɅ�z�s�3�	��i��S�fd��0���΍�=]籛�r�n$u�p�Hk��#�0��Pg�9�RѬ���&s�³��I�b�%JC���O,����[������9*��X�T�Q2������d�����C���8���%6KςF��D�w�F,F����9�u{�	ys�8�cܿ����5�̯Y�%N��~y{�FF4� ��J�	v�����bz|�ov#&zz=oH���Lx�DDD�N�t
#�%�;/t0n��bgw
��K2&y��(fs�ڞ��,6ꍹƣ�h�Q�뒰�W��`�s���K�z���Ҧ��#�Iz� n`ƓIR*����~��+R��8�/dp�pԳsx�e��O�	�aܞo&�]vچpjuNfAIW��dP��W���m���+���"J�qn"��9L�F�tA�A�%ѱ����\�D�����E.1��Gᴓ�kr�����FNv��+ȧ�d�f����JD�yCK|4��Τ�y���E�� ��>�O�}HFFX��tvy�?��&n�]�~�b� Ċ�pc���
S����׼vq��b)�8D_#M>������
m�hIGQvO�4��.��=�G�u~��f�]�$�P�=i~(��І+�I����#����� �� s�t�3�M"�؋�0��bN�����c\:����EƉ'�������i!��ݪ������x������򼴱�x�f��Ǎ>��op�!�;hs��o�HU���ֱ��Ų�ݤ�9<�`��[+&��.�]=c~�PH,_�&��TQ2���"�>������ֺٹ����bՐ�[��D(8����i6	
c]n9$�7ِI|���+lmϘ���ˠ�`��(���f
�ֳ)#|�"��n)(]�]d�S�������2�5���7ޠ3�d,t��׮^3���N�(�E�p��#,.��w��"^鉭t�J'lm���4¼�=���i�VXW�1�XA�y��G�4�~:7i��=�yz�*���
jU�\����b������,�xé~������<��'��&�y𻂞/	a,�o�M&�p�r�2�
����=G�"ܼ6b(���|�Hk������Y	�%�J7�n�Lɗ�R��~��HJ�#�H/������<>x�͏��0����AOP�Y���e�o=d� �ZC\���s @�˫������g3x �^���|����2��C�Ҧ�{��_[Ɵ���6�n�(��D騁Z��J{L���$G9�Q�ܒg�t�(�m�3����ƭ;���GGd�.G�P@��[d/ũ,т�b��txtz>�݆	L4`Ne4�RC3��6�@&,��qW�zH��h�4G6�5�g��� ��gL�g��`]�������[
M�jAK�0v�Y�ެ`v:��ߺ�Y���%,�Q��A��F�3)���;Jh����8ڸ�h/_������>�� O6�P�=}��~�	���x?�g�
���C����ʿ���<>(㣏>3�͝C1�h������J\=h�;B����>�CE�"��mk���3��-,��crZ���O�rf��=��\�֦۩� 9�)_X�u��av�:;�0��]%W���~�<QW�c0���/�-�+ڰ��1`��#+p؟�����7;F8&�m� ��k��|�U�U����Z]v��#4���7}/�Wk|�`ݺx��n3!w�*�(�f���gН5g,f��j�Ȃs%�o�Ϳ�����2��`�S���:�pU�7m��,��7?x�����ߛTm,n,�B�NU�N��8�C8�
�����$r�{�拗����̚�pv�.�vå��Дo��HRF�z=�y��
���y�c;?kع[�9��XB�I��+ ������)q`�YCzKՊ���jw���GOӡ�K4v�@�2:�P��0������u��)�I�a
�&
�1d�Es��VmbD�7"��s%�mD���S���m��c?��h�R9&�a<:*c��Ǹ� v��?��.�\C��M׍ȫ�l[��������y\�:�{��a�w����c��!cH��0�
�$2��n�|i��ϵے�I"��y����HY�J�~�0��Q-�PAZq<���Q�Gn�5��BblG�����j ��+X��Tb�����o6Wl�:3��cODZ�塈����&Rɴ6�cG�Z��[�g�T��XL�D7���n)`3�~� pD]�ft��6ȡ����?��bͽ�=�6�^����3f�鏢֝SA�|�ሉ`�wm�^~�H���d������'����C��}=�"���<�x���%"����٭(�TmFS]���y�k9��W1b�4h��h�=1�B�3�e�v��]X�B�:[�.�p�{6�P�;!ml��!}Nq.��"�_KZ"!6���/�x.)�A�e�@�/4�Ψ`c�wu!�o�Ϩ�$�=�Z��\p�u�]5"�I9���������'L΂JsO��ndS�+
uڴz׍?�i��<k�Qc=�I�������+�sL�"������-~�Ux�N���|�gqk��/�.afV3���	L�fQ�Tp��}��yA;���$ھVr�k{�7P󃚱o�G*wI���f�� {��3��!�}�{����|��cv�L���.9mh�����n�W>���!6Tdէ`��4\�؈�<g�-!���s�F&�J��T��
��}�o׌�&�X:iw�-Z*ձ��ivEqp���F���2�j���u/�Gņ�=��z�,����V�\�i4+h~���'��cC���B'̣07�Q8`�͵j�O0c�p�g��a���#q���ud�:j�iw����H�c$��[��,��ߝ���z'�a��
�Ȅ�7.�IK��M�s�]���JW$�L�O�0����a�_>���f�ށ�?Ą�>��C�����%D�O}�fq��
�q�NCi+��}罳=��~	�q�+,�Rj�����������L3��?)�@���m�ⳛ_[�6���p_�	�7vh<��*�<�.���
�L���+�Xв��h��P�r8��� �Ý>���w:w]ˋs�p9�䘚ʙ ��,
Z;bn	�F��,`@�����s����O��uȝ�
:!m�H0e� �Ւ\GƧ��,���#� o�:����h�ž5��pFP� ����B6uJ��$��ƌ�Q9_��oj���ʕe�4����f�����h�������Z�ň�������L�vp�LΆn�޹�����.#ԉ�Fh�fPe�����&W0���vw�x��M�wޘ��[VݑԄ.�*�l2T�v�b��a�Um�:JW(h�B��[���:��������)d�LS)�:4�{�2tH-�q/��#�����{֡��
9I$䆬�-�@/��ީ�"�~й肙X�ص���d����FgJ���,8�O��6&1���ͼ�h���
�h�H�KaG�-�p�r��W��#�{��tq6�r���YG�Ʀ'VGUAi9�6V����(׏pqm����C�a����s�t�Q~���������x��$/͟�mPۗ^}��kG%�!3܌������Ѵ�\�E����:�u���hF�3��<����.�;���y�9�hF9q��f��n+j���5��>Q�1`b������G��_tڶ��K�7��;��P�=m$P��	�͍��acR6��	b�`'߿�����f��# 	;VbF�=~f��K$a0��R��!�),�g�*pMb9D�+���3�6N����K�U$#]���E���o["[kv��_�/n`_,b�:�ǈ�Ǚ��a��K8�:�յ"Ĭv��ލ�x�2!�B|��4��:�
4+942���1<*�V�T��x���:��tx/\��lt��m�T�
I+���\���v[#�X/��ť�m�;�X"j��sZ��TP��1�J4[�ٝ08�U�,�k�^]]O�Hm�'�p���a�g,� �B�xϱ�DX	�S��]��b�Ӳ�}S�U����Y�����~����=1ݾ}c�k�תd�h,�Z�4��H+��5&fL������7q�b������-ܺ��f�{<Ǳ0��Z������Õ�S�9h�G����(U�&-�_�a�!��A$��c82ق0�S2� �c>S�~O.RaH�n˟s}f�F���N���!���`��`�l��p�|N�#`~7�d��"���*j)X�3�˴�뜇mNv4�L�P��I���|��a�fC&�N��XC�O#�3��~t�-�l["#�T�
l�ۦBTxJ�N��b����Kڹ����3q��1Rŝ�^ߣ��6�j�\g��4�WCg�Eq�H��2�"z��c�@���1.���m씆H2<vjeڼ,�䰲8���,��$}l�}u�����1�_8��8�d���6ĻN1��-��@���t�WI���4FC���"..�2�(p]����]&�����[�x�q��<�rU�C�1������Ҩ�;F��m0��<O��c���Kv�J,C������f5鉠y����ɸ�b�n3M��hbm�T6Fw�u �&to������A�gy��F�RC@���X�oE��K$
�uu~��n�����U�YW�ۭ!R��څe,��Zi��Çx���I:Gi�2��b��)���2.��iC=g����(�����b���yֱ�)<Zl��G%؍v1��~���-����jd�I�p�*�8�� �A�	����~���&�.t�>/�K�&�/i:VH�k+���J�G���\��K�g���p1��j�s�K4�B'��=��>�	��@��O��$�6���e��_�Ͽ׮Ӯ�����RP2M�l��2v~=��
.�Y:KE�
�tfm�Ky��1y0�n!�{u��:��Ŝ8If���`#E�x.���P=�W�P��KZĳ/Ƕ�BX�h�͛��B�P0=�PL��ܲ��~��"���i�4�C TW�t�S]�q�1��%R�݈�4/k��P"�4�:��Y�㙔���h�=�F*�W�U2!"6L
g.�5'� q�F��P�el���������g���Q�*�-%e�~G4f�PQ:�z�����s܌��<_`��Bq3��&PZ������k��[���� L��|�7�|/�q��0b��	UG�I��ֱٰ������w�`4[�K(ñ<3�<?�V���ZrdX`�U�Ĭ�s��U���,���L!�z�d��󛮞O��ϊɩ�=�%�Ͽ��P�]<�� h&� c����L��ҫ�.�`L�I�a���/N;���q}��~�>DG�L��G��/�S&�"�kػM�+�N(�0��퍬��a��k����ǷP>\����i��0�` �a8�ٕַ`���k⫻{���l�?��s�����K��5kg]������j'���U��׺	�+)\c�⡞�+����ښ��2��|U��Ɲ����:13�n��Y�~u�%�8�:>�1���'�/eսՇέ^���\w�k�'l�EI�`�fdc�U�ә�?�
��ß�<�d���b����o�?�� Q}iؤ��+��P����T�P��d�+�c<�{����;��Y��^����Z�F�iއ[�X�C�x7��q��y�pu���=��u��+I:�Xu�3պ����fԂ6<%��fi/ڶ������K-'&��o3(a�q�7S612���5rg|������E���LL�P��5�"�Mtr%c����X�apa�㱟���z*h���ht���u"nvC{m���H�RV�R�Nr����:4�Ѵ�b�֓t&
�����Ȓ�i�E��L�oЕR�������hݤkz]�=���lI^�|�m��&x��������#c�&��3hI�u6���hR�����}��*�?,�n|���$i��1s�m:��������ŭ�2*]ǐ,Y\�����$i�M>\�-�:��3�:���d<a�`�[�t�<"�
C���T�Z�����{2e�l(d��+B�M��Ä�з���+��+�I�IA,!�nFM��8��!IFr�6c� B��������H�,�2�C��X�9˽;U����;6���>{a��
���˳�Op�<Z�O?����42��Ց亴��G�g9�Y*���D�{�c&�=�#ԱW���Ӟ�S�vzdb��̤,��z����Uln��P�&㋡��:��\v�ŋ�S$���)&t�Qݨ������`p���%�L�m�a�3���}0�����Ao��|#�������>>I��؇͹���G����%iN��8�6�hA_	�X��k��G<e�Dw�E?��;����]8��^� %�c���`��=�4��D�K/a�;���ڋ��oL#cs�����\7xv�8:n"�^�]Z�͛B3�XM�=v�Ato$ɠ�Y#F;2��$߃:���9��e*�uK�-1J�\`�����ՎQ��}�H �yK�Q�7Է� ��tc�����z��(�����!#cZ�B�^׍ndR�}t[I��"zN� r{2A`�l���T�ᐄ����3z7꤈�,�5�{x6ج�HӣT�I�/v��aS���:����<A�1�:w��3��gE����=j!�׭6*�?V ��d�K1�乩��m�Bq#�R�6�m΄�Y�B8�`s�%m�@�A̐Gb�6�#�׾��ي"���	�u{�R\*w9Pn��ǚLٹvdt~�t�#��:����o����}G~UPZ��~Qڮ���d��7�b��p�n��,AR,���88	��d@�U��*ڌ��OK=�<<����P:D�X��l&g�o��Q�.&���F2�����X!n�Z�|m�SB�9����!J�(U�ܷ<Ʊ������9̥���N��<A�p{G#&�B��d����(���J�J��l�-��)����U�b���"`~�!m\h����E�h����J{}cPW^�����O���ȥO�H��Gф}�F���n�f�M����n6.��C]�BA�$�Z�a�3��:DN0ү�ܛ�1:.px�0*�D��D<iD	=��<�j�n�J9J��Ǣ/VU.���o��C�����o䆷u�TA��E�ka���_:�����il�}��n�i���'�͐��
��_�'<�QWJI��,��|0g�S�q�<��뫛&OT�d��΍lsm���ϾvP\Ͽ.�(~0(��ez>���#	�m8m_�u��?��$�֥�w~����k	O�ԥ�߯�P��C���7��\ *B\
�с;�Ҡ=���ʁ�./c��,��E��	`�$:x��AG2��Q������4Vf�X�`�Xd@"�n�[q�D�T���g�H=c����4�>�xVMO��*}��`,���0��7��|.mDV��갺�Ic�����TZ�=_�O���_ſ?�ow�l�هC�[9',���XU]3;�{���a<r�ԑj�RV�g�E��J��<����Ȫ�iC2�P.�O1�,दk��_�	�#��&��3�?����g�t:#�Y]����oa��6�m�|�!a]���7_g�e��4l����EB����+�Eb��F��7tE%'v/8��h�ձ�IP�۪q�G6??]0[#��V�ɡ��iv�}?d$�_�ֳb�gH��I>�N���ß��{�ْ���i?>���:�Ez�g�S`*���Z�H ��{'Pq�����ʮAg�UY���%����`X��C�$]�_�r�O��x6��TQ\��o�o`r�ǀ�w�|�(����8���X\�����:���7��3��n���N*��}���B�y4�I����8���u����*��=:�>�:�y[[���;�C����j�x(r$͜�!�QT����̜�XGNL�;ַw���/�`�TƘgE�d2m�`2�U��.��Y����kɄ����f�5ǤqDcs��$�I�-*�U@���ղ�D0��PGp[I}�� ��z�]��5u̸YJ�Pm�,�|����A-EA/��d�a��_�:�"�R�X~ICZs
b��3����cT|.��;C�|]���z'�w߻j�aYsO���wdI�?�G��kKX�]��o_���s�{���<��367j�gQ��y�ZkTAG�6XA�(�D0���%�i����l[B	O:eL�}��I��羄��$����Ijg��d;�a�/��J߯���?�9E^(h�oc-�}�YS���Y�^_����z>��+�Ԯ蓆fx�*_ݪ����u�^фV>��v5몫f��y��g�.VM�Y���O��t<���_�;)-�QRg+�����[�e�������bX�N�����,���v���m&�(m�2�w16����J�4�����\:���u�/�L�tl��S�m<�g�]�#Ǎ�6�ڍ�*V���Q�=b Z�6���v���x��e��bh���6�u�{�ڊ8��U�n}��u3��9��P/���ud��{iԩ��]��/M`�ƙ0rB;R��F'Dk����9�'�F�Ɠ�Q:���:�M�۴Q�ǌ�Ĩ@>����0lE��0��_>ŭa�d ��8���"�������������
��sLg��)q��e�ـqP�qG�L��KM�fS����5&Խ�i�g!�3��uVչ����`�+�<��:�1~:i11��ɑg�g*��9J7f���[���$F�ǝ&���6�W�}}c��ǐL���г���Φ���7~�0�n<���Ϲ1��d���p8���{��n��^O#@#�	�p�-�16�����Ʊ�����7���H��G��dT4F%�٪@2������N�Q.��B�XA��OH5As�t�uh?������	��n �a�\���Μ$$G����ƅR�m�F��J'������tz����靮b���><�'��>��P�3[b�ܑg�וJ�������Ĭ��x9��>Ɵ�x>;�2�:<�ڟh�Y��roDoB�7��S�^U<u-5�'�uq��Զ�Q�b���&�gĭ�b�]���1n�z�����7_�8�|���8E�G#����/���B}��L��c*���Yň(��T3A�=�U%��m�cftff�ljd�㱱��Rg�F6�^�Hy�j�b;İ� ��`��ǳΠ۝��u�ʲU��ω��恔p��n.l�� ]��D��+�X�&M"���ܫ?�ү�<�Ԟ�W9L���"\ ��4���Z�2���H���Mբ������8��̅3��w�h0@�z��������6�x���U�:7����>xs�k�}y�~�h�(�=�Y(5�(?,���t��SAai�Id~�y�j�*��/�X�F�+��#7�N��"�ӓ��Ul�p���t��3����HO;�������QE(*r�r[�l%.��{�N�f<��*8!^�����ѷ�8-��L������|ǣ&Ϥ��6��	l�����}�i��qH&�@��u��V���wV��K�b����֝{4u!}�ҳ���$�����7W�؏/o~���66iX��A��E���<��4ڵ>�6^
�y��L�;5���{[��@�k�۞��C �&Ѡ�#NN��]g��W��\�)74v]�ɼ���K���9,2=Ry��Î�p�`�a���9qhr�<C�n�2N��d���_%�Ϫb�h4�D��z=1��ü��L�\�U�Xp�^[w/f���}��Щ��t����;�u��{��bغ����zc	�+��GwQ���h�(=@�.)�(����Lkq��%��n=����Th�=�J<vAI$��u-�6�bg.R�Ȑ�n2�K!J�6�Ol�ਊR��E�6�4��gK�«`P�Z#�+j�ȟr'�e�N]� �q�'�����!N��ժ�ß��efg0;�`0͐k*������)�g$#�jL��K��$5�II4�>��v5����Ф�}�dw��������%Ѭ�>:��)�O��i�34X[��<!Ұ�!�?޴�N�������Uc�=w������=��
fyt\��\ǿ��_�x���
.��Ǜ��0X���/7��a�g���v�
}u�ձ�#6iZ�JG��C��l�6��>v�5<=�2@:A�gO	���hX�&iK�v�C+��?�rJ����^��m�fTal(D� ����8$�uػ|�M��'�n�7�@��*,i<BE�I<u�D��V����#��K�l�XH����	�B�~-K�ࠄ?�iq� ���k�N|:��2��F1+��m�8��;�^D?��U���LgV氲��d�Cjf��[{X�}��s�����\``zW^�l$C���6���维�eĦ���Lʌt���n�IfB�
�]��}�0��cy�������I�ŻYF���d,�&��Y=��p��y��T�<7^��〯3|�'5��j6Ͷ5jM�s�[��x"��=�4�D�w@�ǠT��P$⤳~1��vN<�לK�@����5�y�3�������8n	��l0��1�p>sh��JTt��UJ5dÎ0�Ѯ����\z���,?3|�cx��_ę�<�Y��
֟�㤴�<�k��>??�q,d
��кH��Iϐ/,ئ���ۨ��p�!�l�I�I��=&4�z�L�%����1I�^����ݎ'<��&�ƧDpR����g���z]���0��i5;�����g�X0�$�����+Tϣ,�ퟠԞ�&J�Ί;A�����fw��*Wj<|��T\���g��q �s0���YH.D�k�ܺ���a�M�h/�8�2�W����QO��5�6�t��N�!+�-��bvy�f���b8�
d��f�31'Ԃ�B�z\�6�`xܷ�0M�L��
�ktB���.W��]�4��WM�!�Y�xnm&����A��y�� ��Z�������&�L����@�\�{T�މe7�7A�r$�?B���	����$�0��9-�e
���۪DLٷ�Ʀ�u.\̞�*6VQO�7E�S����zc:�-�)%E1梉�-Ũbz:��^;�nw�=zB'_7�LkE2;�D~ڒ>��9�N��p
� Cz7-��B�˰5�ߕ�Q���|@���.Ъ�hk��AY�F�c�I����l���i�7q4c=d����_�E�{Ty�b�S�����YRa��f�N��'���p�gc_c�ٻ����0;���,�Ua�|�P��-�G��xhFڈ�Q���e���c���%b8wq��4��Y&#I�<u�WG�d�	�	rub#(.�1��0/ܺD24�����D-	Ü��ٚ�h�u5�`Z�Aڤ��#�d1&-��椘Ct�ۻsr{G%�Ա{Ȅ>��A�"+!܉%�3>�O��'wN�<���&K>C:s�2��eX�S�&i�ȁ�:�`���F��|Fqn��Od�ɴԯ�4���-0aH�!�Ժh��(�s�:�R�9����hڰ�����QAc�1X����c�#|����>�������kQH����;�X�	�8{/���ڧC�`�fڢ�^ϒLuBb���r����B����ϣ���������H������D�8^��`w��$p�Y����N�.�{.Q��1X����}��#�GA�t�#�������c�6V��?ܓP0팂�:�x.����'��fz~��;��r[��Y:�E�l�-]V����^��F?��k�zL�4�6bp��2P��jc�d��tɊ�p.GGS�o��󾻇O~�v�\�"簻�a��[��M�ze
[۸}�3���_���m������ �`E���¡��)�ٌ�N8��BFU�!U�Si�g��ze���!6vw�A��a��g:}�"����y$]�3p�zv��ݚ���ˡF'P��bH����_��Y9nu+�%Ty�Ŏ���d�����&�Y��Y�[;�x���:O;{��*�ZC��� yg�����*��$�!��P�s�o�!$��|7�Ux��-���^�g_��s��*����L����#��hZLX��#��V �3B���/o�c�������7{��>�Ͻ��U��o(�
�B$HI�lj�$�j[V[�v�C;b�ab�O������~�qtt�L��v�m�%��H� A �j_�*�}���woV������2o��o=�9k�(j��>�o��:�A�+����Cl�l�pK����<��3�bw��uQ!i��٪�b/�;Q8r��T 	XÖཌྷ��"��oau++~B�W+��ܻ�$�g"+��r09�]V�r�ћ��ڷ�[����Hi��ױU�+9}`c��ruS�1�d�#��U׈��e[���E�f$����\�t����nro�"�}�N=}0C�V�D7I%��6�?��̈́�bW�Ó����e��~=�*0"�^m��64��S���C�kIM�G�n��.�|�H�5�:��ŴI��--����al>�����>B2#gaf'O."�� ���f��Ph Ec}vr;��vC��2���d��|X2	dA�P����V�%��t��[0�G��$��}r0	t\�%��2.��È�[���1$(p���[n!���"� { q[UjU������bÊ��H���3&k���LB8��ٺ���ї�#��9P�!�(�A�2^j8d��U���k23���Crg��ͻ��Bf~��b�3s]�`@�������u����h����%&��tJySl ����	ħ�MQ�ϝ���AnG4���ȃ���B�!6��}���b���R|aA��|TQ��o����;_5I`���"ɬl%m��zP>��sAE&ig�m�q�눅�M����1���m!Q�a� ����%S*hȾQZ"!��dD�2���NnA���)��=W��x{P|s�n�D�^�l}���`�3�/{��E�5}��hJ�$�D���Xr�����%��K����aC��$�L�'d�r���ǔ��kJ�C�n����p$��HT����Yq!><z���ց*D�?�%&�ϧ����ۊ��Eu����"˾��ae=[(պ�l5M
��������z���-ay?/Yv��qm�c�<2��K���aA�A� %w��$�n�dQL������S�0.�G��d���8��rb� *��R�k��p�E�ؕ@�r��ݺ����{��V�~������7�,F*��ѝg9?7���v����
���>Q����(.��K���lG�T;���S�k�G4�n)d���5��m�3�;a}Ξ�g�8tμ�74;�7���`K��lN�h9�{ٜ�Ӑ*��U�@;J���K��}�n�{�L���R���j;�:���
2���3c̙	.X�������#���p�k�fV��c�y��ȅ{���N|ggSY8S�V���g�QX�2m5�,�A��?|�'��}��2���66�ˣ�t�z[�۷��(�����\	"3�´�S��;=�7CeID;x���{�U�<�k N����u7��9�Ɵ��d�Ne�a8}�i���0[�����bs7�P�r��DH;n��	��3�t�G��~�&�������}�RY>�\�R	�Z�T��hP&&�e]�Tz�s{Z��׈��b��l�\�.���k�uPR<��>k%L�ŝ�"~��U��5	�L�b�Ӯ�~���3��#����*=y��b|�&�FqjiY����#h������݃���K�YS�w"3��K3�j��c����}���{�����6"��*�S�Mb��q1�qI���+�;!��� nJ�R�X�����8aI*ؐ���3Hy�Zې�(��Wh���������#a�	��M���lɞr���1!g�26ԡ�8��qF�t�&�A�>~n����G;�S衎 �]�%�����TR��2�Y��Êv���C
b���d")EN�i	P/���Y�(��Y<���I����W���ʮظ�س,F�rG%��#�%��x���g++ȗ$�	M`tdR4�3�W��L�8f��0W��jJ�O�{�x��9�*j-	i�������S��
���)SޡTm!hqF�:�bЊ�S{��!���S�b}b7��2v���Uk���116��Y����	nK�[��E��*6��%"�%�U��u{f�̚,~v�l�EFцmH�Zj�|##bk��	1���g��-�w$�z����6�w��$�a ���IS�LG'#�{߹��q#�\+ZH�)�D���Ȅ_֭���� Uq��073����zyL�Յ�C<~�X��^�]�)J3qZg�e�O-�ت��$jU��؂j9 kx��A^��!vvsr���|M"!��{��vI���I���?���A��6�H����X���s�u�_�QUl(YXs�Y��p�`��qmIbkbk{�ج5�Z<�؉H$h�����gK'R&��}G��ί�1&�A�Y^��-*N��b*�&"�$�m~{M�;_�4��J[\/���j\�`��&!n�AN��«O)?v��P�3��}MǱ+�_aǬZ�wS�{ӓϕ�ձ���B����!Z]�sl3��ޗQ�\6;J]G	]H
#gC��r��lZo�%��F��ݢ�n��܉��I�[Z�d0��DH�ŭ��O6]9�Wゕ��)d��4�~�u3����|��0N��(�/\v��~E��wQ��+qĨ�2�L�r.�0{�Q�܂���LH����>�}��W�u��O�XCXG���t��u���ld��e�/�|�V���0�.�Ж���=�v��K�Y��(U��T�%&���g�$��a����y.�a�bC$�� �[�RD��B�ul��aA%�)rgus�B�I�
r�sbW��c��͐�~I��Q-^���w������ iV��x	��u�v�J	���V��tb���h�a$�Q/�?9c��!�w9�w���N�\Ĥ�;�(٭�w%����"�ev���Fo�0DB8�]4S���|EI��r?��&�9��٪6	\�����<�y�r�&��M�$��:�a�"&ڒ Q=���S���<bmc�C��%�[k�GB���sp��)m�
����f�G9OH~
� Ƀ�r��J^S�X��&�VX!�~�ބ��(��Jۭ{��K��G�)X�����c�b�0��>�ď���1��R���n�T2��ĭgΜ������ĸ��~��/3���"!!e�Ɨ��z@�c�Hu�QՍ��h(U��f�k����ba�RF9W�j#����J��cd|X�9�l)	֍63�R����#���g&��2���]B8)���\�����a!c۝�A[�>qv�(a�0c�PH^'�xO+�E��%�8� [��\c��N��O�v�bXyT);��"��¯� ѝ���L	G�hWk��'�r>Βu��p�f�cX(�a!�?s8޽�f��q7p���L��
��6֒�h_�v������i1�1��-�y�Fm&)Qb�WKM	n"
HDRJf�Tͧ+�HQ|��������a$-��y��-	�p��	(�05#_�}	3��9��
=�g��>#Ϟ�3N��E�!�8����.R^��ֺ$�����s���}h�i�A"Ă��ձ�#t�k�m��M�v|-�I�q�(���Q�P����{d���;���4�e���NHB���ȶU���*�3b��:o{���:J����
�~�d���/��׮��I�+d��!��a���'3l4B]����8�O�eJF��P�0��W^y�G���-I ^����N#.�����%��Dn�g3Vc���*�Ϡ�:����A-�#؉��Z8ȖT�ݝê�˖�Ѿal��]I�.+��-�}�l�5�^�����Қ�$�.��D�mʣ%��n����$H�M%�ɌaD��ؤ�1�!�Cdit;���̶hżk���6�Q�$�D�)�C����� �Hu�@D�=�D�DN���g%��֤��)����4$W�Gm��;T�^��і`��_�&N/������r�s���Ù�	�ُ����>�W���wߵ��|x{���Pff��Q���+���ED�������WUD�a58ǬIK�l��Ŏ�qX,������C;Q�����ax��di�g�R�qك-9_�7�+�0��%q��v���!R�G4qge�!��1K��DQ���&���5�8��U���!��R:��i��ښ��zէ�/��I�щT�����@?���<+r#��)��>�%}m9�-�����fG�5��8�|�^</������uV��}�_|��d��󳻳�'>���38fQ�W��f��?|G읃�������
�
$
��YL��>I��RϞQێ�}�,�=~�7��d�z�;�g����]�8�\��,�0(�� �֞����Q3�,���XJv&\��+ûM(aQ⌘��h1I�	�džӪ���ɚ�Q�'�rM�S'ŜTϸբ>g�t<��v��#�x�tJB�o!v�8����pG����p������F'�c�R)G|P�BS??gz�}���R��%�,7Jx��		����d@_8�pJ��n`t:�p/��n��be��UL���o!��(�:����]�n����ZO�J��� 2�rN�{H��ou%�}���C	��nQ���$,%YϚ|G;�A���`R>۰���a��`�r����0wS7F�@�54�rP>ߠa����>(�/�,Y�h̯wPu )"����6ėd�7Q����l�Ef<�w�������߹�e�BP���	�K�E���*�"�r�I8T�9c���(�NG�P��K���J[ٽ�.���Í�w}�T�dv�cc����g���$�����;>6�ƈĲ$�����$�D���}�F�W��!�m%C2��A9��#�3s���$6�#cA�E0�.XT��;ْa�e��3I�n��o��$q�.|���̈́�����HkN� /W((�8���ب�vJ�p>��xGb��+�Q��0+_\��ة�؈�2_����nKB�[���@�b�丫�-I��f��;ԭiQ9�*JG�i�HϘiƾ�۴�"	=�(�55*	P��M���rK�����^l�>��� !����I�ό#'��@r����bO�@K�a@	�L�����<�r�lIr�h�KV�"�_��6�*6-1���N������0-��۳z����������4[�anC�q�Z2qኄr�9��q�J��r������M!7?���O$�ے�m(ܩ��zk��A�0`䌓��W�N�4�\�@ @� �� 91N��N����ss�wwG�ӡvo��(++d�"���b�Թ�F���U�P2�Ó�o=<��V��",jL�����ba).	�9nx��P�Xfv\�{�p2XQ�A�Tl5�!\��O��I�?6<��ey?j���k]�t��QY�0���r��t��B,��mM��iEţ���A'ׅ��U0�v��Ũ�:��?�tV���G�^>:%:ov"|X`����:���V�n!����c��\G�nYu�W��N5I�gg�j�P|���}����@q`>&���I�qnH�����*M�𶲴Q����]�d3Mc~!�g% 9���
�>��)n�nL�+f)e�ҹV��]�T���%9��
~V�[��7r<w��ye�"|C�I����#%��_���!ERl�gX��L���_��4v��2`)H�Fb�0�%B1&J/�R�;�l<�%��'ΜDJ��ō�b�=�%��>��8F�Lc�	�a匝�v�Ȃ�;����_����F�T�7�ѐ=Hl�$mg����˳��7*�N8�WЂ��|FVd�+h�����E|���b�ٮ9qL{�<æ8��æV�8��Y��:-�V��!5��ܮ�����*�\*�}(a{k�[�*��v���)����$���B��a�vO�0R7q���:G�w�K�������V�E.�8�ˊ��I�,	�XL;U$#a ��ޓ�� �R�K�N�Ӛ[}� ��Up�	xɠWR6ţg��g�:0��MI�h�9Gî��VM��a��Y�\N�����dX���ԪMuR�;A���������e�� �ti�4�c'�� +,���O���ܖd��7bi��Gu��C��6�gp�r�@�y��/-/ca"�t�Ν���H�p���n�����������Y�nV��	Ya�:�����~[��"���#����<v�����Ն���� �Ċ�!ama	�28ǢX\<%�Y ˟���'�Q�h"쒃��k`�7��ވD˰�v���ܐH�A[��N6P!C;�"Z�R]�v�����_������WI�T�Cd%��z��[GA��>�m�έ;r��j�+r����Ȋ�RHP�S|nkM��>�&/���'���>{�@%�'�)����t5I��Yb�9r߆G��"���$2I3?Em��<�~��O~%���EK����`�ó�.�#������۲���3�s�`d��u8` ����o�0��V�;�]�jMQ=d��s���L��V$�҂2Y��ՙ����7�u��Cv��CdM�&�����Ț&)��EzniDp*���JI2�����=�?�ni�J�%�4��Lf>�wG�ϑLπ���W_������F�M���?Cc4��%���Ȗ˸��7���8�è_�8e���B�f�=��fT�U5DI�������8gNf0*ku:G,.A`�B�ċ;2x3��X 7[�Ŷ�vx0^�sy/Y80A����]$�Օ�|�Q��QR���x8W�dL�2&���0>9��	[b�J;��I�\�O�RG�d&��ɠ��2CMl4�;�����,&�dЯ��������ؒ�9{F��B�/�V��᳓�,.�d$2�#��!e�܏M.���Ν�ۤf]8��&����0����%a�L��Z�;�[Z���e9nЭ���e
-�f#�̗��b�R}�&t%����ZsP�U����C*���2Z�=�u�$�g��+�d{	�q�c��_�w6+�bǵ$����g眶-���������pk/�Q�oI`C�/�mk�>���J��P_�r�0ƥ��$B[�vD�LU�M�)%I(�#,}�㍓W�aa�~���5H)����c��`���
�5�H�5�H�x�����+B�����v��8){X�W019����r?ɡ&��Ď�Z&y�sOV_��F�-�s���!)������1��R󫾹�:w�q	�̙��3(K���}��g~�7\�q1˽n���")�fƔ\ٽH��ζtfpt8��},�nonb%����$�#�ٖ����Tݍ��,ah�Ƽ���o-H 0��/�X}�!�&n�Fs����
�I:�0�����,<V�0fj����z�]Ë�m��v�X���ko]E�sU��*������
$�����0FPK�s�����~\�~J�"ʅ�$)���#C:������ʆO����J�Xj���������qq�8������'1��b9 �ZUEJ9'�dq~aQ�L��E����zv_�
����$�^��=
ݵ�j�g��_(L���n��Ǔ��x����8&S
�ᬆT)I��3w�t�2�m<��t���NG/��܌�Q<y���CI�>{����|n
�~w	ɠ����)���"J��b»�>�a4���]�P�[��a���&jr�Y��D$4$�sZΒ\0$$ڊ�>!� ���(����\ x��7&aP�Dƴ~�T�iJ$�̙����bI	r��fB#Ir!�)I拕���wv�#!A�Ic���X��+c�����
�5Ly��FO6��Y)�
i� 5�	 �A���ᢪ5�p͔`��-��T%�=c0�g¸�Ɂ����Ũ�J]�H�pF���[ʞ�������Lg��?�O?@2Ex:��@�����:k�hP�ƭ
4��X��6�F�������|&�'����a^��'�iR�����#��9K��q��<#�u&@1�ƥ�Ro�^'^Y��@���88�"2x������eD�P<i�����2S�����Gnw۫k�'�����A� ��=��*ѹ&�#���W��Ћ;L�Xi��S�[�b4������19���gh6�3�Y0k!Kh�P<("dI (뒌���wŁ"sj?��?��Oo�}�i������ڛ�X�n��8@]ݎܫťY\�xsS�����n��\�����?�ӵ,�U[�g�fC�xP)�johgY�!�E	�T׮��̤�������꣕m�~gFF��*:Ԫ�X�]3��	��q�KPB�%o���zC)El���.�Hz� ��B�ӈ$���JJx���N�Y�U����1��L<]yH2X����(<��f��l��~��Î|�
��s�8�Ǯ��~~z[ϟ��?�R�5�sM;�b��T_O�H�G�%��`h8)�������2���+��+lj~ig^Y��s��ݻ(U�&-L���~o�u^�Ňѱ�?|���n=�������r� An��scE��nj�3;� ����/�Gn{É�vKb<ynZ�!ӹ#�!�b����ݠ��8.���ﱂ�t�`��E��F��;������əi%h A�h\l:)������9bA�0d�{���ؚ4�#)��R�` K���H(�g+��9M9nb�z���i���=Y�`R�adߓш�S�wO�h;�<Z%�w�$}���,�b�*��Q�Ν�@�DX�Z�#	I&N�o	k=�\a��-��(���Kbf&�"�N�6��<~���u�nJ0>2d(��N$g��^��Z�M'���� 3$�P�pL���HD�BYg����L|��T�ݍ��b�1o��;;�+s��J��E��3b��dT�q�[�ԙ����<�Y0[�1L���#hSv%>���Ң�hf�F{P��3��f�(�qb-�t��b2c%�Đ��w�(�p��ߓ�����m�&q��VI �T;��vjH`E4K����NSi\��5�uHD㘚J��ZY��u��$@��~��M��9l�n� 8G���m��ʨO&I&����O�9eו5`C��mzZlDA�c{���qS�t|C���vǘ���Zn�����I��sz��>Z���a���zG-��LV9Ʈ.���rF��0D2�M�? ��������Q��?�5�Y���쌲��Ux�'O��K���1�,��>w?���y>�d���T_�p?oj�L�|�-�c#+�9���O@�a�-�p;[9I�����Hfo|�ĝ5r~�Q@�� l 4���:�F�1��E�6ϱj��V��Z�v�t��(�g���G��"��(���>Ŋr�x2d���^�]+�����Ϊ���f��B��k}���Q�'"jUS�emV�"��������Q�l��v�v1�R��6�#��b��Ԯ��uG$V͕�0X|Fj�O�7���3���7:�奮Q$d O�ȥ_U�~�B���S8wuIq��rE�>z�R	?~��PzeBG�]YF<IJ�6����t��$]n�gN�PVZ�^n��kaBn�O���dffCb��x�}�";S!�!��L7�FX���8bu���Q�0�q�YH��!a:�CI�>+`:�p+��,=�<�9�[�+n���	q�q�p�4$���=���ț���}	S<x0˵�V�Y�j��(���brI���1�PmF�w*�\/cH��\�����@���;ōn�?��8�	@��1�<�(n`j��R~{[�@���~��	��K�%Inhǎ"���#3�䒨��B�s�Mbx8��:xB�ؙK�S����ܩ��Y�������v�����?�Z��]V*�ݮa��'�ڑ���k��\PUv���*5��{8�?� v$3�����&��������^�5�7�ap�.�T�I�d\�<	j����5UG�DD���I@m8e���B�����PγRс������t
|�X �b�ł�e�l;bLzEqTb�`b����vr~<ZWb���q�.
%���[:s��������++�q9[�wM��?���y�C���)�*[�(\��R[�V���cfd��ۧ��I��yX=��wL�C���Yv	{���bN�,6�֔�wayQ�թ*�`pf詂�������x���� &~Y�(�"݂�fр$�ԦOLKP,�8(����ް�)�'�\9�_�g���]��M\�4��}�[�,���J���Q�O~�+��YK�>Ν��?��s���w?&�g;��ID4<uB������3�hJY�)B�sI���)sj�­��X]{��7��e�+/�쏪�N�2���Q�k�J&~~���^���HХ��j��~X��J�"A�2Wz��fԝ/�� OܻF�m �J�׻���^-+<��v����䄅�vϕ&5	U1JM�YH2 v� v(���M�_=�|���i�ZX���� 8"�L[�C<x�ᡠܻ}�	3J��y��D�9�����Ք����ģ�g��m�#bO��o��O�<o�ɋ,~���`{K��Ɓ��F3:�D��>!�d����eRו�R	�k�nl�W�๬e�X����!6 ��?|xW�QpؗZ��rɊ��� ����kB�r2>�q�5j�ܢ���S�V�M#5�N�����SՎ�m�H�٥UVѠ�ݐ�UG5�Q&��{�H�g
�j/5A�(�� V���b�m�hJ�b;K�i,$�R�Y!W�$?+���p�����_X�a���$�%�M�^Rف��"Cx�t]¥�q����/�Y;b�v��]=�DZM��������ZU{e�}z��6ʒt6�,�R&��eF;xZ���[*�CF����.^���!>�uSmR��Sv�Hb;y�y�!ʝ�dЌ8[^8ef�t���7cR`�cl�+�{�X�������ܫ��94̔��n��D�'�)�����VJ!'A{Q�ް�C-����=���==�"7�̓��<sډ��Z�ѭ�0)I���0�ḉ�%�Ŏ��<}R��FVۣ�!e�,�-���'x1ũ�9LLN�,[�� 7o����ٵ(Y�����ў�'hTj'5�\T�d۟H���ȹ����7����HXϤ2���^��%��əN"������h7��2j�&8+�Uikb���BF]).�G� ��?�0��w�-���J #q�&��>Ц��3�\��@sܽ�/g�3�q��G=_�3�SvX�yɠ�(<�c�M�O�#�f���3�#��ir"��,��뇆Q�E�@_���iQ�ЗP�c�(ڭ.J��$�	\}�"v�
����:'g�d4D���q��	L���]lcvr\e`�P:�.1��I$�Ii[;l��M]\��aq~H�����J��Y�p��<Za�jP�^�+w����Πe�=��q�B�"�?��^΅�ۃ�3���hp�>9=�#���LQfaaA}�g�=߱���9$c!#�ㅣ�����xh�m�L+��Z������\Scd�z:���Aj:I¯�]N�r��/��G�% LɅh����I�q��e��E�Ga��dxq1�~I�Ȃ�H�Ͳ&_-��6��*���[����p4���N��lZ^?�*��#�U�7_{�\e_ُ�d���G(�w� �iP/��p�/��X�����_o6���������Z:8j�o�R�VF�ShL)��D��$�R���zQV�K�g������ɠcR[~[D_�J�|	�?~�4�������j<�S=jY����%\;��L��j�Ή��1:5���$��*Z�����0�9���9qz��4gqP�ș��N���ϲ� Hgv� %e�uۊ" ����0_9��|��M�򛈑Q���0�D@�% �`bz��V8�VҺ�VH� ��g��ͤ1 4�$����;�W�m����:i�0�MM*[X.����}���Nβ<�o��ɺhE�r+����x�Rs��5$��� ܺ~_a1��ʻ�$8 ̒�B��3)��@�T�J������i%=-13��yY�.d%���X��ŕK'����2
�ɋ��~���-���@�)AN�U�	�iH�LZ�		P������%��I ��Y1�$�-���J�&�&!i��ʳ�'W����G�%�P�;�#P�c?J�T꒨P3.�+TZ5 *��'�,��2(�d�Kb綶�0wjх�� R��I��}�,���d��/gI�\l	�J�@�"^u�]\��Đ8��B	[�B3�����K�=CrxF�i3Ө�?��������	�\Z����|���O���S<c�vyY�K���[x�졲�qm�f&{���\���j}�ɛ��ڣ����8n҇��}\�Yĉ�����G���F���#
����&n��\ֹ�A�Og|���|ltݽ����������A0E��[e��˃1�1ƾv�ఋOr�g�R0������rF�ye-�)�]
=J偨X��9	0�������5���wyĺy������ƥ3�0=Ҏ]׽΄�mf��w��]	�,E܄122�[�?��O>�k�N���I�(6z���Vv���λ���ާ���$�y��]}�39L�����e^��I���>�u�-���
���N��2�]���FݧI�>y$ID�N�Y	���h�����sU=ӭ1d">k�=$#�Ä��L�c��sC�Z�TL׎A�c�)��y�E��&�c顴*�[F� �3�L�� wԂ�&g�6wUW����g�#���D_%?��>�z�� ^?g�d��Pѡp�Z�9I��=ǋ�}9�roBShh��O~�!�OMc�ļ�!��!�
����ױ^{K#�?&�R7��Ov����$�w�ӑ`��$�q�a�!9ӕ�~~R�ATKe�|:$��K�@��\�k�W�1c�rEl�twY��M�ayz�n�T���Ү��:��,�.�gr:3�����rǋ˴�d
�ڲ��Ax%1��(�Li2HR6�A�w�E����O��5jXk����L.�_�Ȟ�Ύ9�Μ��W^�p"%�Ql�����ƧFp�l��6^�S�j\���1�v�V?���5�ر��,�hEl8$	E��dq��F�R�L!ʎd���}<��a�ڀ��R����8�(6�1�MM zbJ���&�}=;��$=I�JL�kH\[Vb'��ľ�P鄐s������R�-V:J�]�Y�uM<��2�����S��%�#ƈ���#�X[�)jjllTbVӱt���k��WfG�E^6u���jK	)&1uY�I���U�O����������L�u��#��o�y}%Y��}y��!�5��ds3H��Siyg��?y�j�p��z��ILL���a/�=I�
Ū����EX�d8���ct�Hfg��ZޑN�Hr(��[Α+A ���f~\Iǜ�`��H���l�w�],ؑ¦��YFF�L��ݿ5c:n��\ԙc7��.���Y����)/^nhÍȷd̐��C��]#M�ئ��&鰟���(qĽ

 �K�D�Q9Β�q�����&��^�{�KQRv�s�N"�p$�?��4;+���,ŐI�Zc7*�w~�,-�1&�E��Wv��7��&���S�l�G��i�X�4�[v$Y8���N�|�����&$A0���~�%m��\����0e���ѵ�d˻L����ǝ�A��pŲ\y���*�.��	�c��{��
iI�Τo$�Q�HV7�/�1�T�GǑL���Ǘ;_N
���MdA�V5�ԟ��,��!8�	#�J)�3_��s�G��rV�/����[X� ��5�=�P�?j!>���^���/4qe5�K�rqB�ӏ�l�p�%������d@Ӊ!��fK��18��JH��e�Y����1�Mq��u|��Y	l	�����+��$a����MU��,���+������?L�~�G�BO�N��	�M�B�&{�u��m��K�,�c�bXrr�+4�q`�J���rܮ�{�-��c�0���K�֛�����3���j����IcZ5v)�@Z�~/"kQ=F+�B�n���\:;��^�'t>���t�$�H�̹�J���|�k�19�ƺ8���uݻ�\�rC�j	L`*�$7 EqT�;�3g�ؐe�ז�9�
cb<�������M�"gj�~=��)��6�pj�<�cg0߅���-�@����3�4i��M��e�ݎ�4�S�o��{KHg��LLMK VD�ZA�T��*j����v��dЊخpkwǌ�:TV�;=e��_+�s����^���}��pk�,S�rs�x��a�������p���������LzN��$��rw�:�tN�GN(�s��=���6.J�B�`�/������"��&�{�S��niwm�j�:ɰ��쬬=�~��?�?X^�Bf��onbco����bɡY���2jdG(!�����s�0���88Nw�f:��M"��Vᱦ
nw�I�ǐ��Βb��#Bp���읜�N�h���\��垄]ةA��c� �R��ۅ��l##B��dOG������O���*>�`U�S�!�\���4N�A�{�~���C�]��H�ޝ���k�^�X*���M
�6<���i��T���v�n�����W��7�*�OX\s'f$�q��Y��l�WU�ʯ��&Zu&4��L�B��_���`�s\<��r�@����CqX��܉��G�$�8
e�?��-7����Z�f"��:���QH��s�IԴ�Gr
ϻ�Va�,������IHl]ky���T�� <����֦�:��P���{��P�#�����R�d�6"�=S|6�W�W�"g�󒜌Ex���8����5m)�����O�H=�X�,|���L�O�v0�n�箕꒤6�3�%9L$D�C�0������I��wbr8��W^�u����w���ċ�{8��%��"��۶Κ���)v���0���>�Ԉ�S3�FX�ɞ�S(WKZ���̩[��7�i�-±��S�5���� �?N�����lW��2�8\|k���@����9�7L:���kj����������c�,��i�X����V�BK��1������]~ܕ������I���PH~��Ο�s���1�ԫDW�\ƹsiY�!�K|J�*%FΞ;��d�?z��JA�UO||3��{�P�}(bdxL�l~�g������''�m^|�*z�LGcb�r���;̊i�cooE�v$��N�"���g���#�bm�;nb�5�{]y��bhG��ŵnC��Η�����&�G̮��y���Ub��H�9b�YrE���͜� �-�5-Sb2�p���2��>�//��|#b�9�^�7宋ϖX~|�z�q���GQ⠔��fK������p���%ψ)����a	/���	��nF�;�����AW5}.���Ĉ�5���0��
@⏙��e
Җve�5-~� {�����~	�Y>���{>�U��T� whFX`�3�T��2R<�����K/F4�Yޜ`�q�u��{F͍=y:=�ү�~�����\�u���zh����0;����j��|-��+� �r��D����1:�e9	������I2x��]�;9�sO˃���_0��~�=�Rl.�������%I�x�����/�=�'϶�����s-�gl��5v:f�/M�k�h�m��#���
BäE��m�υ��:�{��Ԡ��<m�	���B��l�BD��Yic�EHu�H��s	i)L@K��������UQ��0F�gqN���ٮ�2�/C�u��/�q����
��1�99�3�Q��a��%�eRZy��ӧ��H�˶��R����W�W.-bjrs�����)����>T�ש�Et�ѵ�Cqڻ�\�U�nu��-�y�Vӧ�H�-�,�{�me��h�F���ݤ�W^�,��F˖s8��{���~����r�=L�W;q*���¡��?<����
�paM@of��*��SŎ,ש�UK�V}5RG���U]����|���]zk��wT�.7�%����N��d�-��R���ǈ�J]��,�J*����%b�4;���?�_�݇8-�̙����������7��S�5����ˤ����j��MqV�h�*ַu���4k�b��3�ԓ@�]R�F#)q�{�B8�}��~�ݟJI�Ǹ$�� n�]��$CZ�6����Է��-U�S?ܽ���jFx;��;���n�0Zr&Le�伆<C~�;�m��gH��(��(!P,�0��n�:Qv.ĎXQ�@���T��a�!�!y�1	�߼vU������x�dUa~uI�rW���Ν)���o��]��gYt�V��pu_����^S�p����v�k�^���4��������kMfF��o����~������މ��y\�����Y<|��]	|�>2e:�&c �"��D�?�F�O,J�|���ݸ!Ɉ��ڛ(Ԛ�y���MBu�:����)��&�{���~y�p�5}��f��"\qkj���<�/�����	�Ǧ��Og�͈�d:r���Sˌv��&��QAO�3lО'�Y��=�����{Wfu�ꪜ�rK�݄�/����m��'���$ǩ��OH_cr����a|�[�g�ȽO��?���o�~'�v�����*��y��3K�zm�v�n�Axt˧ϊ�������L+㦸:��~�*.�r�?�P|��;�=\C���Z蠯u�-%ey����$��L�����WZ���v�u��Gm�
/�
�c����Q�ǫ�yDǳi^-�1��|}��� �O��1QCLc������׹D%fS���fJ0�A�`�PQ�4�|�yV3tԐ���X�7N[�8�l vI�8/�ڕ�t!!~����5<�)�X����pbb�$18{�,�xu	[�9d�%�ML"���{_�=,O�kE�/Ք-9-~�{߿
��[ؒ�t/�S�����&��bcID36=�W^�����M���wĮ��U�F"m��c�)QQ�̖)��W��<@�(�V������V��',o����@�n#B�>�A��̯i��.����5��F�()��+��3V�v��^�EP����U�O�������yE��u�u� ����1ܢ��=�rN���	�����x�d7?| __��j��HL�h���2Ο�:ff���g�k�n8b?�^���G�G
��!I�x�Sj��>\�ƅ�t�~����H��_�w�����w/��a+/7͹�,H�%IfBw����kwu�j��<��b�}�F%�9'g�,�uX��{��U魞s�A�j:�ޟ�/w�̿�|����>��{�w;��w0�QԄv{EI؎��3�F�ɹbB����Uǂ��]�����p����8_���Q䐘��TɎ��z}u�b]�&zr&�Fr߆17��&9a�D�LNL!��Ⱦ��Z�$�D����r��r-�T�m�$~�Ja4=����p��a��X��[��UٳPP�]�E5�����_����{y�jO���
hHr*.�s��2-�Q�u{jP������G`�A8�
�����5ƥ��O��cГuuι�;Z�N��Zb����5ngЧ��B�`�� ;I��pvno���������d$�� �Q8O^��_��P�sY�J�P*����Y��O������6�R죕5���J��P��$r����d�A�M�L�S�1��~���n^��pX�)t����`koO�}PE�_{MYU�g(��u��9W�g��ې�����Gmځ�\茾o^�_/��|���0�SGIxv9�D�$�{0��5Z�����L��cc�H M,4N�HGG�cS����7���\j^e�bh�$E<XB�^6����D_9C�!|��eY��:h[������Hj����TO�\�v�(��[�?G�c�N_:!Ap�0��x��Ǔb��HL:��&e�$YFϊ\;LH�>]��U��y��I��u�-�(����!WW�IRjU�k��n�f�}w��\9��i ?�%��0@$���[��(1)���D'F@�ݥn�j���w�*5^�d�;g��m�ZdUt`�Z:�b� �#|��+8�xJMU�}	2�}˒�-�
`c#'	�gXC�}eW�k[��E&�b��`$"�zK�
j��V��������h�`,��Kq��L�����lgK�>�=������`�����ל�)����~��q,.Nk�'�H8%wr��BrF��#��
��n��� v�[���+/�Ao5x�RSJ�xJI@���褵ܡzjDv�Ys+ت�����&�0��jD	S��q_e%,��SiO�aڪ��Y�̎��䬍nn�_\Gfv��0�5	8O����ׯ�����i��q�����������z}r�����x�,����%9�{�}��y����_���r�G���{�cu�~��w�$����O�A�>˅!��t~f�|����}�%�^.�?�?��?DAlzE������o���5	"Z�|�f�)k��b y�߱�M��������|$|h��'�^�����5�}.�T+�>G!<f�H�ϙٺ$��_��I����g4IF_����{�P}Bě���E���Zo"�~����p������C����/+�UI��u�G++�o��ə��?5tdG%�Y>;�����$1�OMau�n<Az�_���3�^����.����Z�������j�%�C�
�w���ޟ��~���lǐvp$��D:{!��y�!�8!�ֵW�����d���"($��w.���Sk-M�����{U��P��vu��s���u��7�{z���P�zMf�v�L2��W�X_���t��"�7ezu#{��~�t����,���&�"��]���	#�"{��BO25�o*�4+�RKI�pfiH���?�/v��Gdx�X��]��E���"N�Nb���WB�paY�a�<��ƍ_K��c���%���">����ݻȜ�ą��x.	������k��9O?���e�quI��(r��N��K�3�݀)��D;!���Y\:�Ƈ��"«�^U�U�{��.��m�6���Q�MXP�)��++�Ayas�v�'�q�g=W��96��w��Z �}.=�A��m��V�@��oy�m��k1tF�2ݏ�q{Wr��V4&e�B.
��y���q��5��7��e|�Y*���!B��
{�y��\�QL�ELG02��z}I�'�τ�i�on���&F�Kb�~_�]V�<�B*ul��*S�1ćr�x���I�;P������Z����S���^�#ٿTr^��Z|vLr�#M0(%�Í��W5�	+�rT���충��G��d�U�m��ў�[�]B�5%��ĒV��b����7�f�z̥�ʷ�D�?��j)��-��ͳW�א��0?�������P7Z�l�l�kd5�Wߺ���i�lʞ�_���W�bB����o�^� �V Ο@|;�m��X�_~�2�WW��"/���;,ʟ�q�Ĕ|͋�U����r,<���̿���<�����8^<}*����Ą��mY-Sf���{=���7CcI���yh(_t�A�q�c����!\�j-z�)��h��oƙ�d~Q�T,ڊ�qw��Br�Q��
�`Y{�iqq�W^�E�HࣛO��H���G���A�ё$N�ڵ �߸�����6jU���ř����'Ů|�t*�3��|1��eep?W���"=:�sS��'��	���/�r��t�^+\��2�G\�`8��k��h���0=��r����q��Ls����*�&�S��CvR����N�.�Z��Y����oi�Q�4�R��gVhy�	7�c�l+�Jݫ�@�:��u�Y�Ue_�T˻.���������b`��n<؀yΘ��ɹ1\�X����vM����!ع�q��I��]l��V��)�f�0-A����vs�J�14��w��;x�� �����È�"HM��;�Խ�b���t2�7߼�pb?��=4%���A�kg�U}�� ���ғ��[�`k#������ay}�_���a�&.����V�]="�#%0Ɖb�����_��FN/�wv�T�Tx�of�8{��S�2���p��@�J���c��g7��)��*9��A�s+u��lC�=�A�PD7$Q��}���W�o��և�
��Ձ�2;�>,����$!�W�^D�W!Wșʗ���}�]\9;)k���>���9\~�<>��w�=A��p ���
R� �Yl�p��+��$�Fp��>x������"�eH~Ygw�M�bd"��Aj,�X"���@�Pǩg��QX�J�����BzC:{��#��ckF�҈���.�	��Hͭ��e�(�@�ԃ�% �}5���_��Zz�X��?'�!��a5������s�bN�����zY^ט��ggIrBi[lјⓒj�#v.�bi��'G$hG(!�(��TB�����}���(�$�MRWoH�ǒ�S'�w=!��G<���H�
-�)3#�d"�����8��WA�Jǈ�*<[� 		tf�1��~qjCr�.�a�IE�W�R�P�/~�K����P�W<Q�w,5���%G,q;��cI��z�a�d���k�b��	�\7��	R�kf	=��mH���A�1:��`�JM	��$���� �1��2�<L����$�tJ���Ir١�g;�( B~�ʞ�HJ�А�V�UTn��(� �LzB��U�Fby���q$��.�n��"\H�B"�z���XF�.+I@��Gz�/���52�5U�lDl0��:���)5#,t���֪�[!�=�P|:�sB��6^�tV�E��_�S�_;�3�����v=1p�۳h�B�m�K��^�$&&1�Z�{�u�G�I|�͆��˙eǦ��Ѐ�R븣&ݳͺȽ����>�Nd���C���Δ	z�-��eBŹ-"��e;�j��<6H��dk�����	���It/6��JO�cO�_�I4�[�A!�'ϴ�V�����>�����8���K�����)��0�!��DFl�����m��x��_u���p��_��#~M�B�~�ֈ����Q��NS�o&��\���ڮ$�|�����B�O�\�O�����n4�X���.C�J�:G�n�(㸚n�a���7U�[  ��IDATO>MK�|Y��4s��c�!��G����2�O���12j�XG�}���,���c���h�K4��șr���	��g$�[^^D�-uĮ�[e,�L���Y[J��Q�D1d�S#�)��S��٫���bz"��Ks�g?Ɋ��H	�����7�V)��Ü��\�8�kY������?"�l�|D�}FcU�~T����t��g$���'+H��J��ĵ%g-��c�y�%���u����� @�:GQ�A�����I�MS�"��#D(+�AV(9�&�fܦ��(�U��L#iǣ��rC��2��&i5�����v@�[�$���0:V�����G5Lϝ�XU��;��m�by	s���8�-�6D��l[���cmf��q���r�fF�^+L�#�j|,��/7o�BO���9�2�槧TkΖ�5�"�ɓzڽd��lj"�+�Nj<5=9&�!5ԣJ�E���{���j_$�s�mC��x���<З#��
�v����#���cː�y��j�M����`P�9���9�z����_;OjT%pR����U1X�a~n�'�x�pCRU�Y<��hT����@���k������ݚ��c��o��
�31dw����;�V�G1{boO����^�Uq:'fp���p�Jp�lt��%p��<��*���D�H�oļ��bP���9�>/ZS+��İS)ܾ}W�����P�8��V�/dO�kk[�e���P����zY�B�J�n������\&3K_��~\��&������q[��tɈ�3m���Z����&��2°��e�'�adU�F���Ce��Ƞd�r�����RS���~�PƽO�� ���a��k� ����-Ir0�Ӌ���fE	JŜ{�&g,ܿ����ޗ��#h#�N�k�.I�)||�<��]Q���>��Rw�A��w��\�0��wװ-ɍ¯d�4�,B��Sl4�b*�|��$/�$n��s���8uR.YH�[���d���]x���&1�5�>����oF_����)3.��H8�~���^�%4��G�\xhǭ��80Af�D�I���DPa=Zc�-}��bY��|��wɅ,w�א(��$�m�^D|�M��q�ӟ��R陳 �\G�GOq�������^��ߏ�p5��A�x��$�v�ӟ�B�WH1�hW�|_��9�\�DU�uJ����4����˟���Ů�y��-|�ݷ��7.bu������A�(@a�H8�4�J�,g�I�w��uLL�~�tro����R��� +Ȅ�L2���yi���t|��4}��t;�0T�
+e��1��L*���
6�IÀ�o*:j�=fP�z�Cbk�1g��dD�=T�L�VI�c�"=�-X����Π��(C�_�<|�YI��v۸py��c%XY+(�D>�+NV��}'N���eۇ���'�H� ��	��;�"����$��z�ko��/`e�����j���!^e
_�ַя���~�lK���;�x[�[W���'����	4�A�$��Ut���w�����#�m��o?�҅7d��ӛ*M���a���p<!g�%���Uf�n�	���5�n���%�(t����S�kp�N�B������VZjO9�Q�D�A�	9�H� R�3 c�M���'��m^V�5Z�|�W�e�%�\o�gy<@xG$���=�4�fZK^KO�z��_ �J��5Z����5M�E�� �
U@y��\�S���,rfTd�D��y�g"vD��Q�b7���Z	��<M��Sҧ��?�#=�ȯ�>��,e2�Z������_�u�@A��5y~���Ž�Cy�r]��/�\m�y��Cj�����WW�ww�޽���!�ѻ������w�L��o>�������O���/����pġѫM�U�Vc�h̘��@��ꝸ�`O��3z���L���~���Z��צr���Ġ��^c���X��X�����̌�3���	�7�J���=�A�߀��E�t��;�٘g �O;� ��U�A^�@��_p8<S�ϓO��L�0�G"#�J�e����|�L����˜���N�����٪���ץ�`K�tfj��)��@.^�(o~��l�~��\K�m��{�&6d��yY�x��=�5
����`� �#B�SO�}��+39��66�Ʌ��'zV����g08ZMC�2����+g�`��г{��������do^���ѵ����Pw=~9�L�g��g!GnWm���n2P���B�ux*`�j�� Z�Zz�T�HF� {�W�Զ5erԱ� $�X���c ���\O�*4P���IE���%���.?�����Յܾ��A�	�w���<�d[<ɵ�u	�F����bϯ����W_{Z��}���.�����W�b��o�(r�P�~S^}�!�~r�Bc�?sY�~��]�=��)r�aT�9/��tP�D!�+�O����ܥ6����m�;T�d��k�yI�Kl�c#��|��G�J<Q�m�W��8t�6cwNgF���٥8�x�@V��b6a� ���2�ѠwR<�N�-;}f�<j��I5�^��z=�"���kV5��A�m���N�M�R��b�v�B]�	fa+�� }؃�gFVZYB}��<O1N��yL{��B)�z��gɮ1�K�f��l6[�<K�����3*�Z"9�H#$��-_g�ln�KS�H����\Y�؂���Nd��Qf��Ә"W�=�`���O. D�j�#�B�pY�&o���o<Ӄ�������
_��2;�	����"�7(�vM����}ljd��u^B��ٺW���g����m��C�t��<qqI��zS~��?RԢ����ߗ�z=�����\Vú�`[�YC�Vj�ᇟ�g��F��(f�\ٿ�l�?��Mf;�2�,�A�b�y�CX�_=�'/����%Ous����� �� ��eO{z�fRQc],U%�|��R�s��@Э%(E�kL?QL��^i�0�7B�"�2��w��r��pJ@��|]���N��/���e��g-�.F��	�r�����f�����JV��e���w�e�� �Q�}̂�̽�T�B�^({�r�\M�4D0�iЦ?q�O?�\n~�@Ν;+�uV�����Oh0ؒ�m�����IA�/W�\��d!������
�oj@w^�J��$\6��rh�(��*����i��y��M�u�#g�J�:���N�6e������
��k�;>7��Ạ����X\����q�����&�(O���SD�"�,*��ب(�#NL�PR���l��v��I�)` 2���p�` %w�}�ۉ��
�Q����d�(���#)����@��AGa
���4km�mlt������U9Ҡ�܅��W ���-�6[�ƛg����7�W�����3��A�D��̅˺����9��Thp:G�b�������ՋQFJL��<P�tnsY˺tIY���Wn����p.?�'O�ٛ������T�[K�:r��9	f�N2����e���2�I� �%��Tj�H6W�����Ie�Ջđ�<ZJc/�,"����*fp�=��r��"��Ի����Hʠ��	S�R�m�j�CpU,�}L����{�7䥗�e�BS��Ϥ�y�^�������,���\~��'���c-�?{�]�W�/�������W��հ������H~����qq��'��w��޽#o�qI���������d�Ξ����y��?���L�;%������� �T�;�m	o<�����[��>���%��K����m)T�8�Շ2���"��R�JqQ�'�~���`�]��/�	��{
�Gdp�dWVZ+�T���{ �hJ�\Hu�����w�b��Uأ��#�Z�gdE��`<`���\aL�s�1�u]
�cON'����L�������#i?�x���J��5��6�_�Ò�臏��߼-��/_}}W��^~�9֗_|<�k���XE�@��_}�������^���_�+�<!/�tV��ȕϾ����j�!_޼/�����W�r��W���i���(*��>H��Ooj y��U?��ٴy����k�z��EA��P��߽CV�ꜱ�;����W�ǯe�~7�J�:������sBp�ĝXI��
P�ħ�,g��z�؋���t{�Q �
-"sV1��^%��c�{m�W	n�o3;W6V���=��Z���M�!�>�7FM�8���,bOe����ښ�>����Z%��/}z떔���߽ ON����|,E=׏�ٔ�'����U��_>��֪���]��kw��ڷ���Ŗ����}������ O�ܒ[��rg�[&�}y}W^}�����k�_�����w�-�>�*�o���;T�.�]c�>���K��8d������|��'e�������r��P^z�y��v$_~������z]�H��)�OC������Y0G����&�(�Z��G��K�z.�g�����k(�d>u4o��(�V[&���G��ZЀgF ���5)��=��J�=(��^U����L�O�e�lE.�è}�rWF�c�\۔i�$�]ȭ[��9�5+�w0��ƿ�ů`�P�j{����������hjP���֝]j ���P�ѐ��Y��3y�W�e,���,�\�B���"��9��
��MƉ|u�H���Q)��������ޝP����C������[_ �?�n虚��FO��:�9�T�NЋ�T<P0�
վB)t<�����0	��6��$�FM�ެHke]�
J%���XW�)]�`9赡��Za�#V3נ�����4(��P^|zM���s��ۗO?�2*���%=3/cI��+r�!��،�p,z�^y�9�~�ϤW��P�yQ
M_n܄�̐񝭮<������7��=����%y�)���>����b�)˔���E�&��-�Q��5��v[m���yxԕ�rП��qW��O��hF���X�%�|�K�
��)�hYK�H"ق��lq�G�U����V�*�'�Hq#f���MY][#��c�x��/G�r�vD'�8eF�ǘ�$�f���8E�ެ���?Ϣ�LO�ZV 5#�C��E��]Y� Jg�&��[�:8�T����������U9�@-ٸ��e�\F�f��a,|�(�+m�Sy��o((^����g��;�*��Һt��z�c6yB� �}�0+;k�e���υ��4�(�rݨ���Oě�fMl��;���Y^�4����S*ahȘ�6N$!�����6�kJWJ��0�-��2�pt� ���	W!���/�1ۓ�����
B[�֫���Y=лC)�5x��\l��KU9�,%�9+���@���%����a~����?��?�/�ؖ{�����^�^|Rvv#R�p�j�AkJ1ZLE3f Q���]���Z]���Wd<s6�K�� �J��1KR�����I�&����q�3�����<y�8Q�J�x2fP��h6d�@=f�Y�ۄ2P�5f���<����'�Q���Lgv��\�Q*i >{0���Lp�������y��o��������h�a:Р�y��g�1Ŝ�V�5u{N�'�;'}]G�N�RI�kП�{�'T�(~���t�����~_64h���O�dU���^����z"}$���Nu�K�e�G��
^AAs]A4���y��%��?�c�?�ͻ;������K� �F �9%�,p
\�%�9��f��*��'�7�]B�7�����`5E%�ޖ���7 2�����r1�����ZKAk�,�/T�9q�cL��������5F?RZυ0)4��U�ңW�������}�uw�4H���+�vn�~��%GrK#�RS�{S��,���� C��U���?�I�ξ�窂�����ѕ���ջ��O�N�l(ڒ{�(@3S;X�%t�-����u�2� ���s$��;���'/��_ܑ#��UJA���&�"d�XR����������G�`������0����"�]���K�Y��>�{6`r@�	�ع�$A�\	�T��-"�W�u��7�gE?b�tC:��ƒ�v��F_}��| ��7j�� ��_�=��_G
.�dB� �B]���gW����=�S:�z}Y��@K������W�z��k�M�;�����
j{���Ғ@���p"��욞���ˍ�3H����p0��f� ���C����h=_�|�p,�ݹ��9[?���Mn�)'�.���y�T4���c����=�,S�������?^�W���z�泹yC�(����I,�����J������(�.k���`t�19'L�A1\��稚z� v���ex�>8�K�־D�|=0���@io��$�iC>�l$�tK��X�δM�@�ϗw%�^�3Q��ae$�r�Tv:2�u�ԗx?�rG��\�z�}��BM���\��a�:����*���@}kH�����0�Ʌ��}����������1��H���}�����~Q����| H���%��M��@���RJ��F�*��`x��=B��x}W�0�f�N
��.�W�)|VP��0"v�#�vZs��2�Pꗬ�Ģ#� ������?�������@~*_�渕x�A�h.]�Iʧ_�x4��x���E������X}�����Zj����փ�����M�c���a�v�u�@>��Q,/�_Md�
k2`S���_0��lP�l���[����&R.���AE�q�hB���w�>g�$,����^Ǚ�X���53��H�
�9���}$)N\ ���ќj͕r�6E��$�{&bŒ��Ȯb����͊�M�D��b�������U�@ЂA���ϋ��`t:I���e����(�t�ܒ��oKs{!���������YYjW�b��u��LB?9����,WecsE�P������Ri�>t��֞��=���}=o���V��XV�sW|�G�[_ue{���So�X ��7�7*���jJg�ʯs(��v�>�2���\zƲ?�
jS8�؍˱�/��#5.�@�#�?��`�R(ڋ��5F/N-)@@�Z��#B�KR�ݵP�����Ľ�`S�,DdR���._�C�g#��xe�[��A&��n��α��}fpq(�4x��W��2�"wl��U��F�{�3y��K�������r��|~���娓����?8�P%�7/3B���W�E��ߖo�tV��p��cC Y8� "`�0�+mRc�͕Cy��u��|��u�~�ޝ�t�c߈�#Vd�̨�.�6��Wڳ\6^,�Hs%��2뜥�$1TGP��k�H0�&M�j�t�(I4�cPx�$|C+�� R %�f�4�Y��jX����y.�pY<�š����<�ܳ�zm]~����A$���~Y^���L��緥7M9�o�g�潻r�³���UA߁��'?׵ր��o�"��7u]՘)h���MY�s�ƛ��_������G�G�^.�OvWA�^u�&�O�+(|��uWȀey�{,�n࢕h���OyRulW>ߕ�z������gs�,L��[��)����t�p�a�)+u��F���=�4c� ���eLL�}G@ ��5��mMj���4-�4�Y�}8�"���iG������Y��Sp(`�����Ѽ��Cy������l~},?�ǫ�j�2�ʛ�<%�g/I��/޻��j�������ݕ[����=#��s���T ���!�<ߔO>��<��ʪ���=��޸$/���ܾ G{���/5Ry��cNFL@�����a���P��.d����_ߐ��1�����>�j�rN�o�eG_�Pj1�+��o����w�E�2��>潅�g�?if
���}M��CCd��l.2��݊�:�|��#�5�¶�4�M9�t�P3���Mf�^"3�1�H��(%����m�"a�^HdOG}�ygO�w�<���4"��� _��K̕,+Xj/���"��{�Qʻ��&{_�d߸}��z��]���#V�V\Ҁb�������rY��nw��m��_��$ с%�R�u`�es,Hb��\@P�S 똗��<��A,�GpA55��obYLn(�H���1����f�'-��c��g�%����W��e���T�u�w{jw�r��`�x�{�� �F���5��i�S��:�@{Z�<f�B�RIˎ�] � P����:�E�J�(4 �'j��r�Αl�`�+Q��g���w�7�#�&��&ŊF�	ں�S�k�h�+�s���u�g��l���{�@q�I�wt��Z
��ϲ�=b�^cC*p�:��:5��ꮰ��m�ҩ��/��f�¶��|,��&�|�����N�gၩSf��9)J.�N�췞�٠��zE�[5�Ly�=b�8z����D�<c�P���.4�����>Z��9��I{QT;T�j�p� @hY�D���eJ�*%&4���n�;���Cy�;�����שl�d履�Z� ��v���Ӆ���9�]��ϓ�>FM����z��z7��[Ep��?�s���c�~V�u"�#R��\ �a\��GT�En4�4��N��3Xp��[nT�3``\k�e� ��6�HN�yNH�=<��#G$�r�B����?@�}M8�3b.O�%L�G�&��8���>�4YLL�̴@��b��.� D�o�9q�P鉭��c�v�GЏ!z7��58�+�PֻW��`,�PoD�[NZ:�-�az�'��
�u��b��l����0W[�,�:cyȁE��\�Ԩ�����K������m��gHO] e��]�!�٩��`1֌���!䩣i�[���G�ѼS��mJ�	+t�уˮk9 =5�p��`�`kG��T��/�=DR��K�3�3b�d-��p_<�k8<����+��G�����D$?����j��y�D|�A[xo�@�z��S0R��ML?w����EAJq~��$�'�j|r�f<U��58T�;���,!��{����aW�o��
<��~`�t���g���|�'��l��}�Xj�9��̦�<��?�}/6�<��Sq�LN�׳���2����T��	��w��w��衽���k�\�q����أ��3m��7Ƃ`��x6ƭ�XT��������P ⡿��Ã����@{|C�7.���5Y�<�Q��T�s�&h����
lz���;�H>�쾼��S
6_�k_�h�h4���$���+�?���y��#���w�����Z�7X��IP������`*�T�Ц�h�B^h������ �\�i����;�����lmwh�z z�9g��HLf�\��+y���(�V�7V�5�,�g4�%��g�A�1)���M,w�<~l,�"��fN�R��g	�0��������U���	r*�%���g��$G
�n�ۖg��ب��B넙T�0O��k�z������^��8��/��2�o�vN�sd%���<���}�{_�3aG�C��G��k9<\H�}������:�@��v�*�5Aef/��3R��q	�Ԛ�~vOu ͹�#Y];#?��Wj�SR�T,Y�9�|�����3W ͼ\�����۠mp��.=�8*�G�UU6�'�{���/��3�(QD�� �%�z3��xf���,�fʍ. ��H��o+�B��T��hP���z��X^�����W��^�F!L�����|��U��o�E_Z]�����ӯ���j@E�Te�` 3u0���K}�����������2V��
�,ukU��=��υ*��mр�j[�dĪn��F��ϝ��ڑ.{�����T8�		P�����[N��E��`�t�<��9
�9_�hs>���1.��3P�6K���&�9��:�9V:2�`���:�Cw�lkI׵��U��5�@���������QXQ�Lƒ4�?�
3�����p�Aƕ�B:��\`�qY������Z&E)U���/ת6�]_�ނ}�Y��AE*`��D�|�����Z(��mY�-��HZ�Yb��*�L�Z�a��C�:�|�U<]g�TJ�+�RS�\_Lj�A�++�N\&33��y�k��J����G?�n�q�hX����HД�Z��l@��&�婌GS�cd ���������|#��
H�0B�͵�,��ka�G!3�31UCa&��0Z��1pF�-Z�0�,ֽҢ�~p�y�����0��O8{��I$��ctT~ө�v����y���ύ䕞��R������P��AJ�\$x����K����*=��g��PZ}�k�����<��@�����U��ٵ�������ߗR�9��� m��H+k1Q����K�w~`��O4�*C�Z���u=�U�U�g	{��bu�Ƌ��3�X�L�X�D�k��%�b��DbL?+Qհ�g�KR����ykg���1��L�:V���$T'�֗x?&������+r�$�B��Fvf8��Mm%pRH�]���<��/���da��M�NQ�>�+�0Z	�QY�b��}8�Hࠪ���WX���*�`T�A,0�c�d��� �?�8bU6�����a����%�N|)�Kd*��: +�R)��5 ���#(4pZ�f��Aq��]�C�锸�ȡ�3�Ogb�we[�)�Z�n��Ҥ�"��QT��7=J�<�)�RW�|0���Bf31����s�n�����=����ǐ\�!5������� �\~I�}ߨ�3�<J[b�||.�qj�L�G\Ul���F�1	f�y룶qV<H]Q"��7��y@�g����"A��&�����O�$�j�^�j%�[����&�����\-�*��>��ݳ)��@m4�:�E(��"����h��蒙�L���y[f�.�ńF{]y��L�r��w����~�BCd��X����Z<�3�=cRjO�Sҹ�C�P��$�+�>����k��ĝ�.����Zһ�@P�<�g�ViЧ� ��$!�=}Ll�g��I���V�R��j��M�2=��a>u�-|��e���;�r�Ԁ��~���0����4 ��PlVۊ�	}z�����.{�������
��� �G�/d
I�)��Bz��ܺ�͌Z��$-	�й.�Q�@���#~ܕk
���Hn��%��X����9�}�P�u�����Ԩ���	��Gc��?\��J�VW����"6��/�zYRϲ�(ۃ�U�U�`�^h�1����߫��Дn�#��wyIB �0&�(�[�-`p�0��8���d'`&�7v���,r��bD�E�jcY��o瀆���3���jQ,X��`���*2���m�<�i�)N��N�y.Kk��L��S���x1�w?�*W�j��X��`L�Y�`�/�RX���=+�@�!{*Џ�yd[#���u}梼��mRBf�,���DYU�`.���/�ֹ>�����kC/��*��[f&�`Ѓ��5
�
�p����!Д�<c/��3����@�Q_ˊG�+��(�j� �,�5b�
Ȑ��;)m ��.<�FP��@���<�!�BW��Ng4PŒ:%4�<�+�G#Vk���	x�;����}q���T,.�Jq}��5�z��Á|��Wr����2A:(�0^_ݸ#G�e�2��Y*�~p_hi0��{�ȹs����RW �����Z�򚂥�p�|q}��C�����@��L�AAp�*}`Nw�����/�S��Ai��� 2��xKk�<�'�!���V[]�M͹��)�:6`Jʉ�p�����4V�����)��|��yf]Km
�`��t<c�T �=	�<�����5Ѐ����e����c&�t�Je]�2 d��;D��+UL�Dl^+�]A�#gT!,PfE���)��������������c��S���(�=*�f��O���� �[P+Ef=�UX�uJ�Ȅ<�����;�}��b�ot��ͤ���ZVa4x��ZL�!Cj)zΘ��rZW��e���2'$��?����{Gx*��*)+%��@b$�Ψg��ђ��)�[&ja}�u[1�B6]�<�nu}���41�S$=�~t01��9�srr�u�/���Lda�䂒.  �mA9� ��t�;��r[O:^o4�q}ؓ��7�]�#�}
LP�6뾈���"�$����0#�C�ugL�2�wyyC��e��L����)�֯�>��xd�H��^�(N�w7��*av�������^! bP� ��ϱ�����������@p82��Y`�_� ��S&A�f c{@�l�%?q�	��t�D���(A�AX���g@��##�0&����9�éA˪6��id�+ f�@ ���P���1b����
�Ɉ�Rd���
�j/P����`2:J�.�(�T�~$@��b�,f����M�VA��Z����X�aNk��+L>+BY���󇙸��Y�{��p�+�)���c<�H�TIˆ�DA�V�A'����)FB�?g��/nHpQ�)�Ĳ��!X��Qg�)��L ��Z ž.��-�	Iq.�g�+�������[
vO�������H$!D[��h�Mc­l� ��a��+oO9�c����i�¯)�{����ڏy��cE���-�}ЮW�E��6��0md���
��&+rS���,�_G�P��XGX�<K��9Խ�81�2�Q&6�
u*����'��L���eN��>Z�L�.�<��ʴ]I<gۙ��*Ɵ*�ƝB@&��Ղ�fhL/B���,��L��dl��*m;���ъ��֖B�i	f,y��1�	ŰBY�����9�y��5 J7o1OZ��ʼω[��I~�@$B�ض>HTyb4nܕTL8S��H[U�새d��*�%���ǜ�Pa2��#T��?�f��V�c�Zt���PM�S�۝ɵ��euuU�_S�h����
H�~�@z��>pE�bU?��8;�&��޺�˞�=5�+rpܥ�JM�
k@R.#뽐~w$�)���h�KsqB�[(�A�hȍ`!Q_�{(+KKj���VS�]�����a�̺#˞���\����O���0Iz��rn�o��Y4�K�� �"N�Ke"�����}�p(p~ �VŔ��@!���g��..Hf=P�Ɛr(�3{��1g���K �����,-�ā�c�]8<쫁��V�P�L�2��
UH{R1��w�Dz�T�L�����w��,��	��y� �����^^a�$�\�R�g�I6<N-�QqU�h�z����T�-B�E� U�(�ۜ9��i��މ��EcN�4sT8qP�pT�!G6-�m`2�� �N�R-1{����`�p�*�0�f��(	��-M,[O.e�|M<��PY>��]ߚ���@f
6�o��. ��Lա�@}͙�����0�-�U}s�8�$M<��U�w�<3����Af�Jú7�z�����r��vP`�w������F/��6
.��>;zA3}��hJ�ª�y���5T���9��h�������.w�Y���sC�Ĥ�����	.A�[��M5��p8Vc������AF
|^�����f�5��ƝEB	w y4�{�3T2��Ǫ*��� 
{�@�X~$P@E֑���)�ֳʑ���[d���zD����VP�R�K���z�y y'�
�*mQ�O�}�&
�DW�f�m��ʉ�fq�c�8R%2���� �%�x��W�E�Y�Ӂ�^�oV��<������6+̜M�Nq�8W�q��Su�#tu�{�쬮o0)�:��%����X�P��������`�ؗ)2�Sݏ9�o��(�qD�Ì6����	t�PA�"�BA���/�D%{�%�b2�n�c�
3�j�͇N�_�u����F*#���y��{��*Ϟ�w��$3%'l��d��cWo�*��)�)d���OJ/�G��G���ʨ�����>R]d XOc���6,��W=[�����i���Ʉ��B$�R����H �s���5�����=@M�o�� �Dq��A�eɂ	��ĝ)DT�]L�ע�@ �����y6�yhhK�C�㢐���"��jPG�#�a���R	��vT��M�SVq|��aY}�'��&��"+/��=Py��JH(O�
z�AaN���J�=D� I�V�ϭ��@�`>p��^��Y��Ȝ)+Y��1Z�I7��O5PG�g�5$ę��x��5s�i0�:$Ͱ��j���;9��(/p��������ၤ�ޕ~�ϻ�1+�f�[�e�
9�.��5�GɃ=�>5�Rp����Ԙ���5)��4h�X��k5*b!���ʧ�D�Y��3����ofɛ��Jk�9-�*R�?�q�S뵴�,=���n��1��h���[�QY��6g�@0aP�1��\p�?X��Y�����ϳ�k(�a,T��!q�b$�R�4⪟�A�~l�Ÿ�f�ѓ�V+T�L�"��Il.��S�G����^�`���b�ki"R�5�k�HHख़!}VRa�K��d9[���Р�&0a �1�+���A�*v�0]5.�`3W����i�f#�~2C�~9��j6|좏J��ayf��}��"��4r�����%�z���NiW�N����I�5j�8	�<�t�����5_����XB�bw��?�Pa��6V쓁*��km���(a�z���a������n@��J������@6�\o���Q��^�k�3�M��KZ��Y�Q�z��+�%�ؠ��&e[x�Bf��d�K$���?a:gp���2j��#f�,KV
�J� Gۨ4��;C�@�C�g�A�3{>�fD@�R
�yҀг��.V&2��R��#�aH����8z��R��糬??!�6��ܨ-|�G��=GA��3�4��q�JV��׫��f� �&ݪ���7��%���0Zz-X
Ob���dd�X�K��
JP)) �n:�KUǲ���D��CV7�4�A�������	��t�Xr!�LN��S�=)��#�	1�öеei��� lwo���t��h4G���>��e��iL����-0�6�{�1�1М��-�s����j�gIԗP
ui��GY��yG�*fS��)�wh�fE'��C���Y3�^!~��X��=)0��X!Őf��r�VЉ�y�S�xs�tEI~S��)�A��k�}&Z�":f�g�
���orN/�/{D-K���HT�N�:���{:�?�V�)�F[��$�u9�@�4W0�9�Z73��'��/��L8�D��i ��),���N`*�ʝ^f�:2�������x�uE<�L�D)���B��; Qt� �$��AϨZX� d��W���B��˄���ڣ��Y�Ä���K�0����E-�P�y�������11Z����,q":�'=J��O�C&��׊�4�ܿK�����<���1��� $!������G%Pk٧���-ǚ�
���D�����n d����H�n.qh7x|�q�A�����j�Ŧ������-�� C�Qm�@@��[_A�UJ�A�GUT�(8�O��="I?�=+0������Y")�k���h0��0#ݰ�A�hn�' eh23�n�N�h⪻>�*+\b�+�������ĸ%3UVg(ݸ��h_�?�y��+�v��ԉ����_��%�[��7�b,���"��\S��e�r	��!U)�npVa��$0��&P���>���w�lH(8{5��Nd{P��Q�QAD �P�a�f�o���i����D���S�(bU@pf�@@%*�]*]��k22���Rj=B��Q�����"���G�J��o������UA <�]R��x8aOs�Ƃp}3k�`�lߒ����XR�3C��z�򹩒Wݹ�'�E��(��[1Ӳ��8P��=K|�
 ��bD��dJ����f��ժ�GJ�`�`?ث�gg6�����Bo!�BbabIM،�8ɵ2��n��G��,W�&����~�Z�Mt�f�
ŭ�o`b���y2�;YOK����O�D�.���N���֒�~N��#��`QEϬo2������)���WwDB�>����@�����p8�Z�v"�^?1�b��0����`'�5�k'�����g�VL�R�_mU��2�z~1N�#�|��)�3�O�g�P�\�,��Dz�J`�E	�'8��ÁÍȗkMr67<��#'s
�Ў�����:05�0KlP;\J�����v/�xa�Ϛ6�'��� �'L�h��{3AL(G� @��+X�s���p�7�����En$��ɳO٦�2��ف.Y�Z�g/(�Cv!
�}.r�%���^��|`���`��R�d�FB>���ֲ�ĩ��y���ߞ�p�0��>4ܺ�sf�6&�GAx���$�	�l94���B���9��5t�Y���R�ߘ�".x��RpVb��*)�BA���-+�d�� 4^6T3z|�Ě�xf& Cz�`�H�<y㴳�|/8�,��!+3�&
������Ն�C� ��E,�x��#�����>+�� 6�)/+���A�T!����-��-���N�����J���a��bNx��]5ʅ�G���t��[Hi �N�s�8�> �� �Z)���ɌʤX���,�ϗ�Y��%+Ve�UIX)��x�x6��P<рt���QUǢ>�������&nq�\��9�,�Ѭ����3�ܠk��n^d��ʒ��6�f�T
d��и����B����aH�%VH�!�̜gY�1+�FϦc�Q�p�A��y@_�@w6��<
G{T<�cKt�YO��t5s��
)�w ��T��Tq��7����Æ��u���K�Z�Y��RL	�Y�1J6Fk����b�J$
8�0����	3gu�p6u��sS!k���$VP��t�B��'��]�ۥ����[��E*נ����F���� `�>�X��5 ��k0���J^^^15����0I]s��hb�H��#B@�`�,Q	� F�L��Xب#+"#� |���@��Ͻh�w D8S-eui�ʟ:�l�6s��t�g<��'^T-�X4��&66AA<X�pHp`��$�!�$#�Io*D��#�ԒcwN�:�7�	�=�<*�C���!���bRI��luq]*��~�������Y�@3uI;d�'L4�B]�=7��1gƖ�VU 5�.N����O?�j�We��k�\y�U>0,hHh��j,S�q���F�V�\��~�Ijb&��§ ��XT��c����;�ېm�R�8�<�%�y' Ǽ۶Ǹ�FWď��@�?�
����w�ِ싫���(cQ���υ���	��CEВ���&9�?!7�w��|������T_��b�:@�Ɵv�%�2f�R�z��8����h��5 ���٧�֋ϓ�9��Q0f@����/X=���ǵ�B՛"J�����/�ц����#�
� ���X�j�L�� rqV�H䠏AR�a��9g��R"��KW�t����H�C>�)�G�����}Ȩ�p�N�G8C�[��'`��p�
�� i^5rZ�^��g7s=K��|7otN�}���SϒU�:����w�CKRЧ��F��b��8t=ӿ����jK�;=Y�Ғ��G�����QK�я����j੸� F�m62V��ʥ�|�J�sI�,�t�D��¯w�Z�Q%�%��T1{}[��3�Ùx��Lm���BG�c3MN*���9��?�`���X�	�P�ˀ���%�����(���ˋ�������9�R-�мsMP�'�P�1�<3胁o���،�K� ��L�W����5�ٯŁhtm�K�<�&aV)� �<��+0Qh�������zń{]F��"^p-3 Y�?E�9L
B4b6P��(fE�@��>�w��0���Ő��_���o$���o�`�s�g�?q���'�T"�����6�;O��U�I�N5�u��"ā����3p���\��;\�ʠ���i�'�|�"�ąg8ה�<�����u�� ͌fb�`��dϓz��@e�+���R&� �rͨ���$��9\�,$/= x6ÂC��f`���퐍ay36�"T����)h�����SШ�9(���b0t ��K�Ԉ5��X�4.#��6��<z�y%��M=���gV0��c�8	��*�:Y��ۄ�9�-�UƼ���Pbd�砿�����޼i��Y��d����3N!7
��U��%Þ�� <�j\`C�c�x���>{>K
իj���Z�͹]x��l@���6T8"#4��^��#}�"�J5	!����@��ZQ�T�%��%�(�G���P�ń7�C�)�oUN\t��d>/h� N!�d���v9V 3R0�P�0�	r�]^8g9K-�dYU�~'�`sY�>[�uoz�����@|�t��t-
����IU��٩��v0��ᘯ��H�I��,�`��6��h$�@��N��L�FE0�v!�X�k��R.�?��!�+�a�h��)/���l-QXb<2��{D��)��&�:�ڇ,w�މe�<S��+Oy���_j����֏�3(r���� ���,:��x8�5��]���M����6��_���uC7K�hM�����M�!6�4�R�R<Q�
�w&�\���e[�g&�~��M���#w���2x@u�T���k p2��9x"��T:���-�FZ��-(����hїY�+RS۲��)�+���h��l�߳"��Ǵ;>�G:���H��xf���J
��&E5�}��ڷӝ���Epr �Q ����@K���l:Jq��A��zh�|޷ةG����sV�vEg߰^Ȃ�x}$�b�"���5���Ԋ)���TD�.�{O�t��,�Y�(;Q�+:�K޻�ģs�I�H}�^�!��g��"�+}���=��@M�kp����vS���#�ju�6�9�&O��*��D��iW
�ؙ5){k���"`�c�#�%%'8���4������`��0H�d��~zD*N���}�b^ջ�U3�3�� �Ư���S�ſ�I� ς5��q�]���t�+�}�U�y#��J�,r���@�� 4��Q6 ��F��MΦS�{�Ѡmfժd��T}�4���prN刌����uL��ʾ��}#~\]^�����n$�E�6��+K{P���tu$R&�-Őg���α\j���C�����k�RiVegg�	����މ��>א��M��=V7���U�t:R����=9�ز�P�23��$X:$�g��p���8��_Py���<2��[�|�qL�s�� ��bVd�9�3���# ���l/-1a5�ظ�gn��)����*z�`���~���d�߉�ПyFiGk��qρ��x�Tjq�W0oX^|(��uCѷ�`u!�lO̩ؓR"�B/$	��
!.���
���%��N��,)U�gk��*��]�H�� �(�(7��˜E
*��f:�sPz{��wTn=����~_j���Ҙ��ha��x��Zb뙃�A0��c1q�Ő\k~�+�{0����!�O`�L�� 	 
6Nnø7��.��4�Qf��1S��:c���ŀX�$Vu���Br(u���{���̞R��H:PtTW1ܕY�݂�FDq��D��]��n���z��-9��-C Wt���ٓ��d_Dz�_��;��w��:zdbv��B}&�1z��=e��x�������:��W����T�����c�gmJ2�X�����V��c8fl���Py��mǹf���KFP��3X�K�K2Nû@���b��9Q��L�O�j�1�Ĉ/$
I���A� �Br�Z-�7H�SL2u��DH-�`���LlPL��O��a2מ�`f.��Xb!��[R���>�$қ���-!Ʋ&�V��_.��B�Zi�,2�I�����e��n6�Q���z k�8+H@F
ʌ�B�^���l|gQcd��^f�.c���u�A1t���Q���^0�p�Q�#�I-�F|P���ďLV�2�h����1�� �h"F��E_�f�"hLf�Yv��!����F��/�͚у3��(=uM�bǞ�������C� 8m�l�1�1(ۀep��1��ˢ����.�IPІy\�Ɍ
�IT�%�����
�yG���!މQ���;�Ra5d��^Pv�=������<����4��q�s?��0
�C����x���	��sV�p#�;'.�N@�1vi��p�l׿�	U�t� pJ�~�\� CQ���CD'48�p�8\n�����թ�(�=޽G�c_��J��X��D��`hY|�i�\��HΜY�g��D���E_AW4��R�Z{��/P'5^YC*H�@������:�t��^��^�T�k�:�&@���V�.�I��0�I e�Y����,"����L�M��d�Wł{���7$��6�v.sd�!�2P`��)*]<��	R*$`oJd,茑��R$�����*Ðǖ��{�\��T_[�jR���rꪊy&͜�+�w�̇j�"�#����ͬ_!�2pꆼ�9\]ҀX����C���:���h@�,<.+5���l�,�c��ɥK�H5ܺuC.��QC���l_���L�=R��{�9�ܹ�@��H�j��G�-6z0
"< �)D�e�kK)��gG����U�A�� ��"�Vl��ow���z���RB�,��z:tM"�T��AB��	���6�e&�TB�9s8��T8C$4 ���d�����{�<Kms^�v �@��/S��^b�kf�C�v$�J.ɞ ȥj#2<�SJ3��E��{�0ybb`A��QO�Ų{������]m����V㳩������b����a��_����u�|k&�ƫ�q��!{�g2Q��G��9x�}����M��V�� �,���[f��rYЦ����7$e	��c�L��E�#�`�/�E�>1���;g�.�
��5�7 Eb?��5����ܨQ� ��Zϒ�Z F�G�C�<Ui�a�*���jWZ
�ㅵ�$��S$�\a��&�E�������x���P�v�:����j�p_������,��5ew�6�ﳗ�4P8��C�eisI��?��!��t��X� 뉧���.�����{���;|x��N�ɑ􏠎l��i7��m6����U)�MĐ�$�Jd��.�؄YHO�y���f���=�H�Ѵ~>�T�էc�/T�7Ϟ����oB5�Vf������K�2с(
l��a� `݋
�|E�@�KW��)΄S)�O�`T[�w߀!��_t1�Gv�c�����¾�{Eiem���5$a3�ɐ�"�R�NU�Й3Mŕ��ڐ��\W�:���zE:���J�ZݳÝ�l���`w$;7z��}Oz�����Oz�Zk�Ϛ&S98�O�,�MGzFu]�Y�)�+%BK��	:}<1[�٨- |�Kԏ0_�s�d�3H�Y�ք	�T} 1��P�EO"�l���z��S�H�5�go|TUٲ�>w$m @BLd<p
�<1�/�/!�d1����ʖ�QŸ�>��b0b�=èb���삏��w�l��XLt�`��&��
�r9`f�b�
�ML�}�H YKJ�xu(��<����u���(K�cHP������b����Q��݂UU�GAj�	l�g-�!�e��Y]h�J��Z�U��1�yϞ�j+a�@��<�w�*��Q<��d$sÏzv'� ��資��L������Nd��?����@N��8��
GY{�@<+�Ⱥ�� ����'h��[�X�D�1���/!kķ1@�Y)�/��DK�a$iQOd*-��(��$&TdzEPp��(�K�X���`r�oI�T�̤��7�6�-K�X$ux �������9#Ðe��irîir;��Q�@]	[-R�P����~�(�;C�M"�^Gǖ�B���r9�]�#(��A�g6P��	�ϙX���Fut�U�4A���� �<�}#�NXe��NӲ�t�(B�� ��&]K�OA+��ŜN"V����˖������}Q�ϲ�<r�#V}-d炔u�7ז�]oJY5ΐb��1�^a�|�ʀ��"�z�Ќ}>.����h���3qP�3.�1�ಡ���S5
T���yj�_PTg���nPf��n��P��ȍd��0�2p��Wp�])�u��5`�� jjb3q�5�7�.��\���`d�P� �
����V�"A��(�����\��xV�0���f��ǵEE��^A���h��g�L����:�M`�6��Ɩ͵Af�������e1̤�M����Ȕ�
	� Tb���jS�B*��Cݏ�u����7�@M��cv��ƶwxD`Au�i�{�p�YI��Zf��W�ɣL݊�U��o��\2����'Ӟя�d���rf�àQq,���5���`}g̻,��5[��΃����f��i�&f� ��R��Jl�d�qw�4u��!�/q�4�↖t���S�$�캟Dg�ه&2��Pt����x�2:���6�fIYfAC�J&u5���y	�1m�ҹ��yfC�}�\�xN~������������@A��2ֳ;	�6ڞ�k������!y1ѯ�����)C�?�T�}p��&�.
$e@���!����ʲ�7�����-�O��ޖ���
vٓ�0��@n���2햁� ��C�G8��*G6��z�%2T������;��=���gs�s��5mfTBR��V�-���,���w�� g�� ����
'��	��z��P�T��8ؑ'�yB�
�#]�'�b"��n���?�O�\�����������]��X����t�>��I�#�Q�bg�Q[�}�+@�+��!^�䨐NgLP��>��}Q�	�X�)�&P��#劮��T��o�gdk��vF����P��6w�R4��p4�����~��ڎ�"��:Tt-E?�%��[���&:C�Ό{��3�H�K���}�8��G����"[���Zz����?�D��Ç�r�,���&�^~��r㫯����O�Lm��ͯ�J�{�Y9�ߖ���˗�ͷ^��?��᛿��������޷��W_��\��y����z^.\<�q6o���+/˿�W�F~��O乗^% ��7�JY�iemM���BY>�N�0�q��r�$۷�H�%o����y��tP��3,�%�%�~3�Z�Z��ܖo�����x��ا�v��^�n�Gj�˗(�stܑ���~����=JS����-Y[]5u`�V�g�#�_�"[[L�T��������#P�\ Ȣ2����<yf���a �J,뛛��=���֖'�}Zn޽-�G����<v�1��zݎ�:�P�Ƌ.�z�9:f�q^��ܹ3��T���-ǝcy���#�|~K��]��~������2"'.5escU.}�r�¦�5*l�9E�|���?���\��RM�b5�I�m3��'���nO��3]�tA�z��O�|�	����ت�-�-|}��%y�w��ڋd�!���+Fb���ch��Q�6������}���z�1ff}}����r��]�wpL&'V����	˭E�z��\-�~�w���b䊍�0&,�2�������C컬{R�����5�������xT �����T�]���7����������?#-��_} so�管�r$�;�K�&ҥ�C��E�B�s[��3��|�\�|Q��->c�ZbK���!1��5΂<T���>���_D�b��,<���Q����P.o�$o��2YH �Wf�j�`��^���j��'����S����<���C�I�sc�ȸbw��6�C�i�b�#�%����ef0�nl����'.���3�e��� �����1%��
 lp]�-�Fd��V���!��B�IW׫r���'��"��JXS�^hQ�Ƙ���d���%��z��dy 0�r2X�}$B�]�0�P	)���F��*	�A(Π/8a�x�o����Z���"u�}R?Ш]���@�j��Y�F=V�p !z�����Zd���gEf�tJe ?�<�z��
�*�ϰ9�"fЯ��C:<��3�n����C!(�Ǧz�l�&�HC�+��r������I��j�YЌ�Q���n���07�jg���đn��#5P����f1s`N&u���Jfa�� 2J#�{fj�w�$���}A@Q�0�%�����87e�̚\:�$W?}O���F^~�;�v��we����!�k��
eR	��hF�M��+3Y�4�@�ݣ┽�����2A�~�#zf������zQ��7��QI}�G*��e���{�z����陜����>u�+�0c�UP���#���j�� eTҠ�7��9b�XZU�s�gT�h��@ еJ�d� �g&�P���n���x���������1\���],=>��-)��ՙ%z�P!/V�llC��H��e�J�@�2<ڒ����^	� |0P W��R�<�s��`6"H�ԱV5���(�Y(�!3�sk=�� {������ZM�#/o^%zU�V�'r� �h�U&
Y�)�2��{5�<O��D�`�N�d����C`�Ze�υ�aPOP�� H��A���at��+*eD�O�¡vD��� I�(4�Vg+�§�3�ߏ�7ӏ8gx���f��-� �!���P8�لc2v��ɽ;���rMB}�w ^�xV�Ё^өye��*�Ѷ|����/d����7�{>�ձܺ���s�4��*��5�����*�x&�)6�z�EHH�]�0��`�OBYV�����PgT�#�OM�E^}/�y���Fjg�m�}#)T3���\� ��Π����kP�t*��co���1�2/��oVJ|S=k 8�{�%�t�1�Ԩ�G���� �s�B�_އ��M�r�jS���� ���&Ӎ9�f���Zh�6�����T�}�U��府?�"w�Gr����9�&_��K�疼��[�G?�=y��'9��^О���*����;�
���(�q��-V#V����i�6�t?��l59�g���֖|y���>��"����.��/�
e.�FA�n$;��>�������a6�74�9���,g�=xp��$EP���@jumES������Y�X��}�ϝ?��J�]����e눊�`�d.A�9?�O��|�5��o�Wy�[o�O]�/�>����֫\������$o��ܾwWF�<y��6�����lnn��/^�Y��w���FEz�9��'�EA�4�w�ۓ��_��_��sY������g�����?�p�����&<��Yk���2�G�o޹J�[7~��lK����U���O�w��~����vwq ��9Yk�dǟP�*��z���f.--��Yu@П�XB�:H���FQή�}0�!��ޡ���㝎�����إ����=�C��rv�)�B�l�zy�
?��2&�D�gOƇ_1�C�!)M����A�_I,s�d\��tT�eR����JIz�� T��#=�J���̖e>ؑޡ�Ͳb7u+�^O������������ᶾ�\�v�y+�,˷���\��۲ЯM��ș%œ���kIO��RM�R)��̧���./�p��gˍ����^���H��u��+j��dVG_���k%��~\�o8���>�}e�RXƇ��\@oy2!S����/,t]�*f��aK�mAe�icfR�g���
�����oo#�k {F�5^}R/��@R���ƙUVwF��z�e|p�&b�-T)���#$ض��Mmf�Fj�j�We�Y���!�i]����כ5Y�^�a��s���<�������h4@�!��@$Ȑ������"�������a3B��R�i@(+(f6h4z��+盙7��g�^k�s�`*\�Y�ý������Zh>̆Ju]h�w���Dz�jh����&�~� ʳ�\溴��T�b�-f�o������\���2<�T�xqC�t��Ο�k��翨��\c�cƥ�lW�dU�y�@OGGR��ׄ�m��nn��;��*4(5i��P<�nE��c���i���q$�´xAU���ɱ)�O*պ��Hm��t���뷷X|x����y��H�f��i`�����l�=+��@���jEv��2�nˡ�R��͌��d�쑑?Ev�����G�l�<]̞�+�D�xC�`��#(��;$ӧC��D�I$ϕ@�4�9��:H�����yX�rEyp�����y��<;=�jG_C�Y���@���d�ʐ	� �_Cg���!>�|?��F�Pl$�(���*�f���)0�ޙ��A{��F!H'��<bZ�`c�y*��`��zA�/��{�뒌�X`QP}]�x�!��!����@v@5Y	�N��b�bRL$�Dy'g�qQe����9`�e�����iƠKBE�F�PR���p�|NxET�"б�3�$�^V�1��%X�f�e�c�4���M�Aw`NM��d%��ꔮ�)P��X��@���!ޓ�&9�Ԡ^V���;��1�>#��� ̈OY!'�2p��$�Q��W����F����.���?#��{���Ư˯}�-���3&>����RM�mh�8���Թ���̌��Ls�
��U��cY���x���uM`��4�������'�X�<E�����Ҡ��;����t�1Й��ȍ�טl?��� cB��ji"}T����?�Pd��pt)A��@p�
����9*�HpN�������	g]���0�0�$"�8t�X��q���@V]����ܸ��鵟�y����q��\u1��뽪������e�S��ؗ{w?��&ɚ�^�>��&��y�W�_��&�o}�u���r29����	���7�������n�@߳���p5Գ6%�V�C��A��:�Z��Bqb¾�f;��px��+�?{������.���a=�|��*�w&���(f��_..�5��+kLȏՁ �AE�փ�X+QJ%��
t�V��b�j���
�rHb!���d4e���:�w�~[>��}������3�9��umx�	�X��?��nU�����TGM�7@F�iqF���\���B���V4�?���֪����4���m�������Oߑ��~&���M04`8.���xE���I ��'$,Iк�<5b�";@���(&L�a��P5���E�D�76��q�\k�K�\7�.]��Vh�z�3�Q�>gr98�lx��&�(:/�T�Nm)����]T���,$��i���\�q����V�G��}h�%�+ZnKج5���i�BTo;�>�R@�{�F�"�Ȃ���F� ~NVeM]ג��TJU��At����6`�C��F,����k&6�x��oʿ��?����,>x$_���)'z�-�P�2�NZ]ΕO����D�gE����.d9�:��B���کx2��d_�_�3�O>�E�&&;��&�-	�ԙ4*!��ᮨ�������T��`����U��� g���.'��)ˑ~�V: �8h0�o���V��WO��L��&;��~�s��Ϙ�����]�>��ь'�=�
+e?�\��V(�|Ni���3����t_kȦ��R��O���P�?�'�'R��Lg���lt��}$�j݇���}�ȿ?z����@��}Ύ���3��sNƇ�L5A��n˗߼&߼�*o�ɞ|�#}��'�`J���?�@���?U����{��?����d��L���#��`C9��ԌG�k�������B��R�@2 ��c�m�%s��<=��\c��O����p�273�Ձ����gg�9|r�U9�Ʌ�?̾EɈDA}φ�C��g"�NOz�h_W[�$:gIf��(6K��!@�M6w�<��tO�d(=~�I�ӻj�^���)��C�����vN4ٹ��N�v�5x
���H�\fjs'Gr��@�*�<����lx"��^�m���sy�Ɩ���~E�O>��AY��^�-=}�������r�g�B��T1�q��39�$���a�~I�i-���&+�v_�����T�@�{:�̅^/
�,����/�ĕs�:�M|q��WU�׹��L����g����]jG�t&��J��N5#qWW��jw��W0��uE6�a�s_M��ꥹ�+	�09+SPrW���c�F�u�	)�S!N.�$�C^�C��������TR$xj��Zԓ��bJJUK6������FH!]�Sؠ���&Y0��a�略O�U��*K��ѯ~���7��]���YQ��"v���k���d��W�U�g��$�J�߀s�(Uu�nV�\'42l�g6�Z�2a�莎/���7����j��UM �K=���k������:�;y/)�I�$��zB6g�
�4��j�W5a�XmH[c��Oԏ�=�K}&��/���f?����K���> �aS��4����p��fCc�9����1�K���)M�����PR��50~Q-��٫���xΙ��.�I�e���yE�rR�I꺇>������\)zRԄݚ�/gu���@$*��	[��Va0]�����W�찔1��`uJf�3�l�n�>���׾.�wV�{��!����_~�&1��e��+���0�0p�k��*��&���N�L�H�,9]�O�y[.b�Q <��`�B��ڀ< �����H��\��ؔ�C�dzx��0���?���[z�+�!�Co�B�)$��	���,*~%��㠓hD�'�X1.Q��X޸�:b$|A7s� ���L��oK����Ѝ�F��Fd[�FmE�S�/M�@�]�>ب�H/e�	S���Ʋ�uk�����H�G-�����"]�x�I�Xj��?e�73K����rH�G��M����H�����D>S�}xg�!vP4l�W���T��Y���u�5���hZ����x�K#�
��D^�z.k-K�¤��n̴���πb�k���tk��M�,�&�V ��0�O@)���|�:ą:��Ԙ�H �K��Q�Eu5����NΪ/Z�7vz��R'�.�)�&LA�?�ddK�v#WQ/��smkzM��\����f3�;����=�X�j��5X�i0�����}���S�sN�.�����e��K2>|$��6�ۼ:bb��B~X}�3���w&��t�N֌���Ya�?	�Y~��K:x,��u�QW�g���S��+��(�Y�G�X�A ��[Y���^���K�׹��h�n\�Y'��_7o�kpQ!�lu��m° ]X]mjҼ�#�{��hV�����R=՟D�%|�]�̈�ΰU8���@沮����ֆn�C�Є�$�DKu�lt}�h ��Fc��?Ҡ4ы��B�c�����:hu����@����uʍ�7d[�����ܟ��)�M�;�,5&uϪ}���⹯��3�jo��Fv1a���J���<}�`_���Ti@�$�7�7��L��ӳ����R�;a�Ä�?��vû+2���P�a�EC�S� �v�9�v931<'nW�ݖA��������:���:T���X��%�,}k��P�y�j08V{�����ir3����&&c$����L��U��&�$I�ak 0k�g3D@*�+�7�oj����7���pW��ڶ��rS~����o�X~�����@i�Q� ~��>��������<������tu������)eRb!�짺��GG���7��X�Y���<Cc�s�:�?����Aђ�~��_�b�N}ch�%5���=}�I�T���9��g��ߐ|�E�����vu}�:�0_6RS6�frr�1�t ;r:8f�'WR�$����I��ٙ:?�3�������H?U��':�9|����n}M�����t�2���WdmcMmrW���L��P̛hП/b� =&<Y���Ư�����K�׺�ݿ�w���]z[,f��6{k��uM���.Ԟ�ܼ!�4y|��G�jⲵ����9I��%@ �*<:�M �]�׭��������wA����ʷ�IZ��QpH:�3p�\Nx������_�[���Ȁ��4���7=�����1��6�� !E̱��l���u�o�z������hb���o�ş�û�ڸIF�?�mU�j2I&������&o~�M���*�t`?�|) �8��@R���4l޵�.�I��Nc�"����	̨3���T^z�%�L�(��R��[_xS��/�G�C#�~�%����N�`LA���+��e���_���hwCMAl��H���*
"��&����w�������=�\�K&��I��@������S��h��/|��X���^���u��t��=�{�o�\�D�G4����Zx�R�%me\��&8���yM`'�ua��)�����:�ا�Z�W��MMc٭�U�+�tO����^����i�SdȯR��R��Lm! �뛄�'t���Sx�,$�D4��"��O0��~�{���Ϻ|�~S���`Ou/OA�1n�`����3��o��
�	G����-�z�����e{wK��exy�n'�`��	��SD=�̴e��m�����&��O�{�C�]�׀���1��v�(��F�B PdZm��󏓡ڜ��#j,b6y�"�������ki.�]]��뻲������!�hE�wB2�xn��+��h0~qf�9=��a��\6-��H�Tb�������<9Nd���>6%'9�W�����L�d)M~��@d���s�PXd����������#3�^N��0��{��lC"��GLz����f��FPE]�NK��z*w��6�0O��9h�8:�t���>���a��<n` ��ڬ�ڀ�����\{,{��Ǝ4�<⍥ĚB�W�&�'�ɑ�:����e�����]�m��k�V)��<�E08Q\�v�x�kib��� �8�s4�I���d
x*3���93ؤ��#��dfՔ[]�ݡ����#sTYV�|�8'1�DR-�\e�6R�B��J���S&�j�/f�`�pB����P�N��)c%(�f�mF��˷��_i�9�j�C����n��Aa�����\��Y5�� %|Ψ�B\�54hE�6#���ʖ�9|��~�z�F���J�3w���� �����s�{��D.8��9�� �NG`�G�b���N4H��T��5H�j28���-�`@C:�S5�`�B%�ځ` ��j��%�떪���!��תֽm�l��ӡ�=���	n\ہ:/�.u5Hq*Ps��pr�:�H��l��ՙc��_�NF���M����5ܿ/��X^�=��7�ݷ���3uX�{�Ͻ.o��M��|�Dj�3]Cu`��B�G���r�z��͚�N`>"m��x�b�1ˆAq�ߓɐ���j�]��2����z�I
6��;���Muz�d'�T�z�cBH/��ӠM�� ��1W#|���n�hkK��>;M�_痘k�����[��:�+��j�� q�I��!�bɠb�5#jʊ�[o�f����kܬ���/kb��=����q�AHfv����}i����K�4�3�=��_�-�5�L4��]�έdC��[�n��N���ޞ|���u���$7yP�&�)�l�7�L��DTj;�5S$j�Q��*�da�t]��DU&@��>x�@����������[dS�����I�����`��p��η��\�d�x������V�ZSG,��<�N��O�<~�(��L�����Ӂ����w)��>BPY�� �P��JmH��]d��կ��ۿ�
�i.�ɂ�D�r2�}7��`2�AU���P��}=Q�@�g����WWz�^�qS�`�D'�-�<ړ_��W�������C��{C�ƺ<�?�RG�����qTq�4�8H����=��oF4+���-d�3�t������oG�����_P[�6~37͟O��5*��sZS[�59x2�޵�[��7�Ν;|]$<Лԟ�\J��y�H���@�bh���̃�����~M�6M8&��gz]?�?�5;��_�{4�Fg���Q�2Kƚ��{D(.�����/I�oL}�!��(�{�s,"�\ �^W�	��ڂ��uØ��h��k`���:�g�hྡ����XX����N�?�c��u]ۉ�/���ɗ��e�~������i�ٖ�����Suy�8{�����&I_����ĺ�t}�T��&
U�3j��+m��L��B�
eI~������k����zK��&Q�&��Q�-d�Zʙ��	���ٹ [���̦�� 
@��ì"Hn`����$=���|<��X�x��aq(��W�DR��>��Ox)uQ�2Ŵ���I�I�~��
z͘�B� (�'�c<���i������?ԟ�i��n79ڳ��Չ����C��U}���LG�ob�@���~�3���*Xn���ԄzEm?�H��{�֕��3y��>K�c��.������{�ȃO����.����>��n����@����>Χ��W^�͸p���9>ٗ�n��B����lI���O��
�R���?�w~�=��g�����9�����(��k��s
��"�*��́)!��ș��
�\J��&��QO�`���t|;�<��,�86�ާ���O����`9�~�d �h�q	X���ui�Ծ�B̓�3���=��c��ĢuC~���8��z&=�����"F���Y����=�ߜR/�4&ؽ����9����9�F`�cHE��a1�5�dҍ�V�vCߣ�v�ѳg#��^�&[��R�X1*����Ƭ��Z��i��q���ΰj�=��bR= L�drM��>3�kM�q�Άg,P�͗���8V����_��:f�u�N.�߿�s�я���!���SР�����qoܹ�ڞ"��,�k�+"�_�,p����\Lt/鳈�=S��*��I����V�Y�M�06Wc�5Vhh���{TÀ35�P(s�Ktv����UѲM���Ā�s�j�*�QAN��,�@۷ݬ��ku�?���S�ssWZ&�����1}�2�$t�y6BO���q��I�k5�#�ji>���(��L~�ߣ@�^w��s��Ey�)iSf�d��fR�`��F��`<K�^>�MM1_� ��'�*�:�u�GÄ
�t���U���75Ѐ�~,s�f|/F��rӣ)�E�T�8�db�kk�խk`���fEǾATH� ޘ�$��ĀC��r4�ĮɎ:3�=M~�<<he#�S!*I;��;���xs[���NG�T�n*���m�A���tրW�G��U&;&D4b%y4ք�[a琂�1K.�N�A�`nl��P�cy���k�j������X��-�gU3H㍽9�5Ⱦ���d�L  ��5��t%���B5��n���fMnj���0�xo>�Ժ� �7���}��-���3�9W�,L ��$��Pgo���X��u��&/]ߑ۷n�i��� ��uo!qB��iҌ�'5 �Z�9���7�PC������N<+�=�OF�ǒk��������)���72��n����!`�B���bȢ���&���8����qV@	 Q���������]��r�3ߨ�h�0���]\��F�����e'��6��Zut��A��:��iv[eY[_��)�.�#Ώ%i�ؖ���U�]�Xu4Y?==���		�s}|�C�8�x�l��f�Ɯ��$LIX����$]߶���������6���<��nʵ���&���SV��^Iɘ����k����7��=r��l��rO�i�z���B��]Afsz:����ߗ�w굔���o�_���u}��N�ɮ��S;p��KO+fP)#�s`R�	{���1��Z�d�`Pj�>�IaNv��uij���#��򦞇�>��@���p�0�9=�ԫ�P<;<�D�__G�/<{@���ݏ5�[5*y��fSbGڗg�鯭�4It�1/�M�K�dfˀ'�fVhLmb���w���2��`p�����ͻ|m$�G�������l>`;��P��-X��m AŅ�F����vZ.dV;:8��Ǿ��������?����/�g���3���T�����5�;п���_�����l���ЏIh��}����r��8*� UA!׹�6����9�c�����yUn�t[�[G�έ0�$�����@���L�>������G�5��7��������9���,�^+k}�퓓����[����P���?;?c��~�� ف�9$i`���}T��-0B1���\�7�����ѿ"�D�1B��)'q|vL����m�!�ս��X%��\��t���چ��� L�2��l��Z���,���������74����do�APEc��&���-i�لNm������?E��It��BR�Yb���QPB甾:W;:bp�{��qW_�Ν��7��ٓ�d�F��t���dqW&/\�����Ϳc"XDϐT�v�X� ��{���,dE.(A�Kt�P\E!���5�B̦!�?�Fc�$��W`s�b��.)�]-�S���>�=����yL{���9�����\�o��[�E�b"�%��{�������MH���V��Pqt�C@7��4~��o����i����y�k���5����uY�\����|��O���R������9�_6���$/@��C@(bb򓟼#shoB�U�������ϼ�li���ʘH�� �]�Wnߒ����-<�=�X���],�쎳�lI.�nf'q��w�a��d��&��D$�:�EƠ�Dm�5&���S:W������$��d�B�X�\�:�����:o>�$Z#���v��mʝ�ޔ����sM؏�0��}�����St�:j�PL-k,|�qf	��Gj�{O�'8�(WI�n�"��HU��d0�SMΨ��Co96B:�@�@^��7�L%�"R�,��4z��
�@��yqw[������VW�ۺ�{C��GOP�Mc�^�V�_͑`d�kz?���d���L�Y�Ĉ�� � � `��
�ˤ��͓�����5�]��a~9��|���MGF�	Z� �QU�:V�̓���H���m�~M�d��C��A�$���_5b.�ĴUW;��m����Y�!c,��KF��o�0�6JdN���(ew���.a�|&�5�BB-C�&#&���F� {�+<c{L��Q书���D1I
=�aI��`_�7���:;<`C�� {���y� ���&
	���	B�q[� N�� !Dv�ﭫS==��?��LM�꺹�5�74���B��a�mr�!.���b�ݕ�.�\&�DF�+�*c���K=x&����F�1u!��i�Jz�&�v��+`7���GGP�e�
�IH
-=T��N	��/��lF��dG����&��c� �ld���y��OO�dM�����H�AH\bt��j��1d�[;j���o�;�˟~�	WU��e�ءB����TyvV׍�>!�f�(�МZ�����F�F5r��]VKK��D5�Q���G�0. ֽr�N�3�r~p �xb60MT� GH�y�q�ƮLu}�=zL����x���U�����p��;��<���!���P� n���!^�m9|�H���w[4
��T0��
�h�Az ��60�"�ż��K5�XT���bo����ɐ�@$�
���[}�N9�A}�/��� � �M#���O���L>��C���?��XdK�,T/O��V�@�}q�{�ڒnoU~�ܧq 2��\-���Z���uk҈n2����}!(< �����]H�S���)��E1M)̸�,T4��t.K������h[:�֖>��R�#A�����Г�� �	'��Lvxm�k�+���"��ͽ"��%���P}tl����/e_���N�i����=0ܰ[��j�V�w�V�3����7�\p�ȫH�p#��h5
�����$���L��?f��!���p.z�����+Rku)����K�^��P�'��r�D��|K�(�Q:���&�g���c��|���kr��.�I�(38l��&3�ۊ����9� ���_���=���h�a��K�|�ɠs��� �O&��
:��$��^�Z�p���1�{g��hJ6+��qet����w���]���%p��I�P	��uʓ�#�+��-0&��Z�0��\��cT�ʀr�E�o��Ƨ����x��K�u������~�ѓ{��{<=ܓ��icF�H���w���7_�w��}�DA���S�z��X�;��*�~G���b���H���q$�O�<��i�J�%M"Z��!@7
�	�	�6:��[����"@�B9�<fq9�����V;|oh�!��t����p��3�% �@v��	�!<+���4�-%�v���X��P}ywkM���P�-�����A*�h�y���P!��lv�疐%%�8���C��'����.��g�^P:)ԆG������2���=��Yl��G�8۸����ә$�\��`$|x_�UG^{�5��;,��T�)�;qn7����_�*��i��������%
R%�	��H�P�@y2��Q�ι'$��L�00!t�k���D/��A���AƇ�2�7X�4
��iV�}�4d��{MZ��[꘏�K��ty	���f&�뇼J��0	���=
�I!M���y��0�%��	G�����s�$r� ;�AyL�Mf��q����u������/H1��5.�W��]��J�gesc�,���Խ�N!�?&����o0�L�SC���e���EC��������ܱA�@�Ԩ�.4Mh��A��%��Hbq��0�����ff��ٖ�oIkmM����j2������bB>J��� �4t���	��E����
�Bao��L�s��}+�Y����(��F�J
�+�Z��`���+yTN������x�ޖ2��j�8G�$Y��(ȔNX}蝫��8��}�!0V�z��s��"b^�ڐv�#1F70+]����ε�lƮ�3��������,��$(&'�Cq�A]��4�>l��qn��н�1c�N�hIg}]�v7��� �(�T�=2�%�dx	�:�J����3�4�?���$� ���MN�r�`0F8��[ّ2v}���/�gAe�� 
&��7#6aL�?��(z7X3��Ʊd��Vy!}@�R�`����7����%�"�b��~�ߔ|w��O 1@���-�ըj�u�Fp=,$�a]�����.2V�ˮф�!��f!�I0��K@��)�M��X�&)�j����&�䃟��*ҩ�[xu�UA}��4����0s�5aRTm���F�����#$�u����gKcop�ԩԅ���%N�@����������D
g�����.��MkA�H��R�kU*� �a�A��
�A1���3�(�p�������Dj������)V��@P��$�r�Ti0�KId�m5頰�9Y���������?a7n��Jc��A(��^~�%
ݢ�C�#�1�_��	������G��ك�\&��R��	a�1w%�P�D;����@���!�� ���*F�oq1MMM�И�:`�b��B������H�18�d���ዼZ����6zR���oӐ,@���R�)�@zN��a�0�,>DVq]5 ��?cq�/�4�D��N��wֈe������c>vJ�	H
'�Xt�j�|�Ş�XaP��Ua@�Q���lln�[�.,:��9t2QEI �%	�����"�d�sT�Rv�I��9!���@����Y�;}yAݬ	����Hi������S�]��vάKM����$i�3x�T��ph�$zeә%:1�ԛ��N G�i"8��8�<cR�IHJ�a�&�W9۪&�ph�����9a�A7�cVN174A���a�����
k�FR�:�9�~��Lc6��Z���Me_q8{����V�aɯ�j�\�_z�����>Fd<CA*��n8fSN��|��Y��¿16 ;��0^،#�C�F�.�
+�{Q�J���"���H�����ZR��m�I~S�����	*� -
�j�L]Xg�9tuR/lF0��HC�h�˹������ �p3�55xу r�B�(�O��KQ�p9�_�l ����Z��_���I��@��.�~�d�拷 a.]!@DuK�QP�EC��r�$��y���/E�h�1���FDc3��1'A�~�<˦֔��=�s�ycbB��跰�9��"��d�Bm��k:��Z���V�6 �=}���;�E�-!N�A�3f�'���db�B;�7Jl\8��;�)���jY1id@��̟�o\�ؠ`��Z�����P䃝E5s��st|&w��'a�k��Wk�;�GX�'�&܀a5ۜ�m ܖ28[�#�~]B�"���:�+�#��`�Y���ݟǐ���	u��%�\��dL�(�^,@�Rt1�O�F�7��1֚c �1�����M�m���/C�����}�
.�$sc��g;g8���[G �6D4�{T���⩡�F�ז����.����z�,�
I-��HBӀ&̬��8l�g �A�dY��EL��Ԯ�\o���%���Y��ՌqCƅ��2w;��9g��G��FhB�+��0~f��0-_�0�NMO}뵗oK}uE.�|��Uc؆�`����J����&�c�*��&�-�Q�	a��lFB��z��=�AN29v傆%�A�� b��u��(�����$�T����#kl��0��'{�d&ߕ����	�id��8S��+���@�88�&%�
�+}^�z�ʳ�D��L��x��"�}>�:�� ����	��XHǌ��NA��&H�R+�s��o=�P�)��5���ԿWd�8���gL�3V�����5��iWC�Af�歙.;:��  �k��3�[����i�U ~�"Wш��d�ش*���$&��1���17;�Kĵ��ÿ���	f�����?��*>p�3g�ˋ��U� 0rFL.�&m�� >�O�zJ)�x�0�Z�sA�Ve�끨������<a5[�<�ɝ%P\S,`�6wB� K̊!q;�J�ǯq�$7���4���b���fvf�B@\Xq3�A��7�H����C��&a���?e����A�H��6d�̌�����Z���C@G��.�݅�\N1���LH=`����tt`��8��?��H�Z4���qN��˪1[a�Aj�ڑfF�F�{�f�.`�0�f3Md���d�͊~Jo��"A?\�y�cۈ���Zj�I�������_믰��3Q���#���k���M8 ֜ݖ"��R�Y2�B\/��8�^�`�F���q���Zp U�Y���٩R�Fq����ĐYP:�ud�m<�Ē�<Hlm�q}�2��1��hVI6�i'��_��D�'�ud) �s�L���g0H$i) a�*u-9$I��q��J���c�Q�r�a^h�Q%a�P̢p�I!�&u ,��f Й �����<@��3�"F�5`�ݽFg��F0���0m'zY�!��w2�CEr��쇢�`(���FJ���)*}q�JlH�BN�J�2���8��0`�(��d�=��WC�I'ġQҳ�{���q.��46���d<2&�up�@J�F[�řKD�sh���e�ܒW�,21JM�M�:tv��X��R��A2��e���}�5���$���\#�;�����^Nym�VG��M���Č�&�����,��<�9l.�>cN�EN��ٚ�.R^$� ͖�v���گdms��ث�9f�ІO��0 �Fz�jg0v �)�AX%q�?��W1�D�GFn?l$"�+I���e�� 0�H�FEMh���}mxkF�ùvO���x��kHo�R`O}x���hߺu�]�X}57ؑ�yĵD�K�3}�`��,��~@p�y�X����q�t�$%��%޵�kd�q��X�fI�x�v��w{H�F��[P��X��gBg4�s��`"��u�t/�<[�xgQ�M��U~��Fk�k�$�^4g�F�ɒ�RH����d ~y�,*�z�ۣ(?�,^x�7�/�E�1���҉d��`�.�eK�#�1�F@�s����܋�0w�b�׈�2{@�%1i�%�P�:�H���
��uә{\G�#.��{��W)rӍD�}HcJtMn��Y�m��U�́$
���w�r�CE"�N�k��-$r�iD���>�m�f����s����5R1~���Q.�.�x�'�|v�?���1����>�K�ϼ���J>�%A�ja�K,�8!޴D�;�qf�!;��,�F�A��d��ϧLާ�!m�5f�<��ϐ W�n�͗^&����BFj0M�G�Ω҇"���5`�9�b;�5���=Fz�c��gp~��q#���#�A�E?�:@�����k�)vi�e'�� yq�E���F�?���0��&�Mr� z0*5�䣻�e��+/��04��)X���d"��LB��B/"!&F̊8-'�b̸�3���7�4ER�;m�u{�n�Eqt���۲�ׂ��T,�o��=�#@�y��%3�/秄:��yd�y�l2���$C����PxVa�aWi�
���\��o������Ha�{}	��;�~𖫗%LM(;
���o��C�IX�v&lT�Q,5E�\��K(�>)�8�Pϐ�V�(�F�MK[q��� ����=��t�!H\!ك /�N���I�j�^����Kf�CB
����f(+Y�4�xh)�X9�l�H�э"�O���az@�TW��xZb�iS���m$U7�0�D0No	�pT 6&U��aLB���֫|&�\h�,�YBzwTl�%-U����Ò\�#�R��̓�B��0���X9�8s��%:'<t�o8aPȀ��� d��M4[ܰs�6xv���₁	�	���U�ܖ�2'c�3Ne��9��$� a�H�0��~?���53� ˠ�L���\8ό���1'�=P)D"0�FB����1��<AEW!p&�9��ܻRN[e��i0����s�jPEd@���<0��ἅ��Sǒz���<�1�,BFPMb0��z���R�J�w���d_"12�&P��뙆#�`"��D���u�Co`Lap`����d�%֘��(4�)2��� t-87�D�r�
�vv����{��e��H�����G�?q��Yn�Ē�t����,l jU2U��'I�U��A0I�-
��J�:ْI���c�
��KbP�frM4A�d�d��.��YmѤ������d0�R���3! k��m��7�IEBX8����0��kP���3���~&�wv�C���|�`W��ģ�K^3:p��3���p�!Y~�}L�~œ��9$~���>����I)�$����
p��]A�1�l��`�:��qn����	���Gq�{p�'2x"��U��C�\��1�w;�Se"k�Y�3���M6����C7I� �ւ�?���e�M��gQ�?���p�9@߇��~�:uE/Ǻ�Fܒ�XtQ����/��gK�	�Ps�4Q�<��L�EW�Vbٝ�:���U�1[v�ř��]B\�΍e��K��6�<�
��!�M%���*�1��C��$o�����
)��A+�9�h3!�{��8�)�Y	�?%���\4���t�M����(�D�ۅ�y��;1�����}�0����ߖ;�;��8���29�X"�1Z4�U(4�����E�H��Y8��M��H8�p-�΋�M�S�`���8�b����>V����a���eF,��q�k��lJ����{Qg��p��:���Z�/3�� ���׃�gf�
��Z�2�s8�u�*�'�\��o�S��pa.�����e�MvZC2�#���r��#��*r��^��<��Ԣx\D���[A��?|!�IO�x��QϘ�[�����"��`��L�,�3g�ק{���&/������L�����N/G`�Ib����'E�q+��n��ʊ�1��?H��!oS�q5ē�0���nȽREQ	I���<��@�GaT�R�w�zRf��~�4D�;~N����KH�Ry$`�����v)W|6G�C�?:m��l�"n�X/p8$��A(�FN�ys�÷ ���d�$�Z������6�u�	��<��o���f{�פ���1b��~S�+֣q�=o��(d�K_$$�2A���c�V�y���K��A/Lbu��λ?r�zRV*3;�Øm쀱'�?[<Q����K�gn�W
<�,ʗ�W�
�X�F��|	 ] �̈́�g�����wJ����B
Y�.+�J�u� ��B�$��g����ipM��gPR��}�p~7���c�q�:uh�
�-�%�Q~��D<���HY�O(�-���b���>rO����Ĭ�~T-r;'�b���A}����:/��T��q�I�,#uR�衶��8L�I0Z�4�a(�L��K��(��85�䢮�Q0#x�8�]Lݜ`����Yg�ʊd���lb�a3 �	��U#����	=�_�sD��p����Y���Z%5a��o�$��q�	A��	�`����O�Z�^��I"��Ab��Go3S�O��8A'���tҰ�\��0�A,���Ԫ:���ZP	�oV�l0T���3R|/`vET�񻜫���1�����}!�G������~�a�Q��Y�3���9�=EW��:ЋC���d �X[[[�SS�hʁuS��Xّ`�/u{`(�I?�-$��
�Z��y2������$OP��!ܑ1��Ybb�`sE�
���K��	��ȖCDն�/1�Y� ��<��4�ߵ��x�4Ya�s�U���"��lh�R�5A0�uR������œ�&η����+l����"�LP������h�N�|��G,�ߚ$
@���P��"j� +��Q�ݫ��f��[8�$�8��Aj�Zh�Ng���6X�>-�ɭK�DC�ɞ�ϋ3��}Hܞ1Lw���7���:a�!F�u���YJqa���%^<�"C���X��?��F�L� ,��g1��n��Y!�e�g���Ofu��_M�� � �* ��7߿�9Z�/��".ܫ�Ug(�5�WP��:�dʆ�&s���܉�+�Y�(,���9q�H�Ec�v��x���f��}���h��@�b�	#O�p��<��4t�:=V�g�؂h��J�mg����h)�3���@nٵx搛�A
1�<����R��0-|��~"d���{Q��
�3���ӨF�8�냃}��%׮k���p}���DHn��Ι21psU���s��^XA�;	{e�xɉHR2oۺ�,x��ˋ�r��,R�=�n}NX�����?C�qDG�y%�q�-��zo�~�2��d6�z�+��Dy�[+>n�º�%ں�FcL��d8;����7ȟ�/7�:d�-�٠��D�F��,e�hN�u	�ƌ�>�g�d1��rhdDޙ	L��	�q����}2�����i��L�3~P���:PH��E"r.�$�z����!�7_����������e���?���\Ɨ��ؗ1>�g������S�M��ԾqKVvoh<X���sH`�HDR��l�εP�(��(0{H	��%Zf�Hc�L2G����LJ�2+���;�k��:���k�ɉ��D����%>
Ek�u� Y��0�0b�b$�)	�R#�J�A�q�M�;��D3��Z3�6�?@�+��l���l: F�YB?1���֙�dzX�0��>V㴝k7d{�:���V6~l�B��͡wbs&��h�/�������#9�J��P����'K?^��T�_��-{o+U�;X$��`�94c��s1����y�8$��BѾ��(c ����F�K��D���,8+��"��Qq؋�ߍ�7g��C`�Z�P�.��c��:D�ي"E�����]�~gW�����n��7`��A�䊭]mK�ܫ)f�,�@�ǋ�o�>�J��\��2:7�S��o0��C�!<�M���/:8���Ol��B�d�*D
-|,���N����$R��'3^��0.�̪yj$��� a6ɚ>h�!IĽ�[RA[�ݺbx=$�L(��f?:S���Y��Y��e�;�@.7Ja����%N{F7�N�ABY�LzQ�C'l��@���o���yW��e�C��N���>Qçr�#���64Lخ�>&H>s�*������J
O�',�$��(���Lx}n\����9�����[ToX ����1��x���m���rHے�ԓ���A8�H�%ɖ>"( s�1I�,f����mP8;8��c��T�!r�)s�{l�?V-7\Qm������	8fB#&��f�I�R����	�I��G��`��sF��*4$��H*
�?�; �&��<b`��>#�ǲ(gI��"��%1	�Q`U@~�;(�8bG0%�ϊ%ecѝL���g���^�����h���y�W.��g�w{@�S�"2��2;�c�`�ͷ�ELah|�].(:��;���*�D�HM�J�I�@�� ��3��%�S��IS��z��y^8~�#��,a1��B���$l�)���S����1CY�V�g;�-!3*�*�+ʫ5͗��绣Kx``���߄��sK�ǀ�}{��W����l�s��)���/���s:�=�K�Ĭ.6�Hi� �'�3
2�ͪr< �n
,1� ��@B�����#�Jyp�D�@鳙�Nܣ�VU���$���NM3��?�dP�_D[@���e븋�=�m��xĬ����Xƙ?��
m���rճc��`CHQ�������?�����(�PH�1��D;�Z�M�(m��yQ�΋�'�1AD�;�g�@$4�h�z�m�C<��	A�/_��1{(���Kh�W$�$��sE�� .e�Qέ` ��C��ו��M=[�Rk�H����	�M�l��^�q@��E7�AV �l�$p�]���+5���Q�x����}'*2/h��4�y�j�ڭN���4����R���ȁ��Ҩ�n1�o�ށ˽#e4!�`�	aN&��(|�|��f��V��A=������ڑ�oK�ד�ڪ3ȋLf�꯴z2��0Y��	�$7�Фb2C	N"��l�Ȧ&��N__g.����/����am�ɲ�zk{�k��S+�J{�D���uf1����s��3��՟�7W��sy�[��Ďqh9�p�򪑈P�ׄ�V�t��R�,|4�I)��r��đy�%���O�\�E1��X�k� �.��0���h���fM�+�����80G�ad,`H��Qh.��/��JKT�Ԍ9۝�]�~M�S�C �(���A?��Ż�}Z&s�w
��OQx�z	;����~'��Π�̛}%��X��AK�/�n��e���`3`PO�C �5f*��?�
U�9������x��&�`�lI���?t!�Ad��˨�3&66�j�:]���=v�J�-��/ ]��A�:-��<�O��W���H��a��@Յ�^z��=�&,.��93&S�cWT:��E�xoT���nU�4���>f���/�=iw\8�#�0�9�V��#JBK�����IE��b$��� ��lfX�Z|\@x���JuT1h���Ov�H'O��U��$DoA�tYq�b5p���H6g��r�a�Q%B� g�gI���B�$�϶"*� �H��#��I��,%��� ������j\Q�t�iaf�d�[,�X[�_i���͎&Vm5dM:���{��gd��+bݏ�9gZ��4��ۀq�H��A-ll�x�VMw�^ͧ��k���c�����|���0Ʉ�������\��͐{���n�K�Mv`���1�IQ1��]��xPdL������9]�񘠱ǎ���������aQ�3XƁ{��e`3)�Ef#�Tq�"�oHuu�ZO@�\���-��I�@��� �|�]O1��;��;|/�"C:^�Y'q��0<���0f����̢#foЁG2�L1w=R���#MgD&@R����פ?v�8�r���6[xP\���mʖ�g��F��YP3A��"+B$�"����Z1a�w���_�a�bŃ�<]��	Y�����r���f�\/50O4 �O.�0Q�ᔊW��͈�����~6
(�ʉ;�*��]����C	���Y(O�#�I������,�T6��R��9��Nէ�j�߆��]K&��s$���f>�l.��tI���%KB��`FF��|��7�P�>��`ݍxĺL��J���Gv�s���k/���H8�bb�nS:��[�F��?�h8�'�ROdZ(��~ ���&�[}O����	d��d$kN�`͘·��"i���<��c�O���(�����	vlI�\j�F'�$�Cqre�ϵ�:���RvE��r�-��n��H�X$�R&-H�ᇐd�'�Q�Q3�lcQ��ݮ�\[�If��?dERe��$�`��f�,L��*wV��{]z;74�I�֤���?$�9wv��S����Ĝ��G`�d��E�z��j��x��*sG��E�=t��M���EƖʎ@P[W���"�����&�8_�K@�0z�H�n����L.u]�z�5��6��2��$�!0G1�f<`����om���ߠ���p(�x�s�{ A��=uÔ~9H�BC1����Y�KU����[R�ܐ��m���LƧC�A3����|ċ�1�$����ɂ*V�Ɉv�"(��'�X���g��1���'	���XQ�6Yډ̓Q ��v9�q?�H̸���S2���Or��9����$�2��d���������8�G-֔���f�/k��Ի�c��� ��`����sŕMBE42�3�ڹ.7n�@�p��!���$P9�~�V��$a,��������E-�����zQ0�|��!���p�X��dg+08If�:3`�0.[fK}�9�� ɋ̾Rwbɀ���;E�M�R��=
��K��l6Kx�~�:eiZ�PY�&��sn�ݼ�,��RǱ���	�L�<�n��~ޒ��b%yQ������*���G��+6!��y���$V1A�;	�:���'����/9�� |�s��:eYh��S�(aާ� ��ˀ��If������o,����|�K�m�*b&,K��	_�,N�*k�&^��������id32_2Xf�JH|��.1�Cv+�تoА<��ӿ�5����l2x�%Ol����~���6�� m?�v{`���A��PMt����Є���c��$DG���7A2�P*7�XJ� �a�W�d��Y�P�Zw�ed Dg"���g��T�w�
�:E�san<�H[���?�{�Ч+ a����H��(�NS�:�.�J݂��1��N��t0VZ�pЍ�������]�@@���S�z���Z2X�BKDW଼���g7��߹�n�pBtiS�iJ
pxҞ0���G�Ȣ��'h֍$�HZT�\�Eb��(L 
55i��(� �hR5�Tft����\��(��1���B8��]�4M�1��rDW<H�L!���%6�0�NjnY�2��e2Q�Qp����E����R�����@ K�TAg��dK��.�Ӧdrfd�H�#R�;ez���qF��{�8�$��W\a�E�n;:)��E �X� h �@�S1-��U��w��(t@�{�z�'�vW:k}>��M.��l�	a] ��~ �G�Q��c�Y�����٪ 5�?)KЩs2�8c����������,Y� =tۄ��,���ᲙBhS��~��ud�;;>�������N|�Q�����j1[����_̪P�l��S�-v1_C���1��=�O��om	��f�嗓!� #)ދ���V����L"F4VW���D"��cx|$�{O%>�A�#Bw�.S������X��pqVp��;����;���i�5������0˜�Ņ�x�M�s���M 2�D=&��nx]<��gO��s3uo/ȼ���3	H��Y��!$%�А(ZR�9�����h�-��]^@�>���xk����;X��Pױ��{b��R�H���پ&e���[\w�O~rO�)�B&��c���勤 ��;����R$������E���^���QXyQ�y�I�\2��wa#�
J�]��=�bm�s�L3��� @�kC����A޴��i���7�y�hB|���D�a�;��о�bJjs��Y��䍀�
���\C�H�oޖ>t7a����^��8��&�c_�Lp���8{��20��Ӯ���d��lݼ%�VK��:�g��*�k�u+>DE�MB #�n>{nq4m\��LZ��ɄS��<�+R��0q|�_���Dh@�@�����9!S��b^z�x���)��N-g�L��]�۟�J��/��md�`��I�O�'R��,F�&9�\H"�(T*٘������O�f,g���g<��D+��n޾#�[;�z&����c��L��ϬcN{T
͂y���]W1M��{�k~f��p��]����"�}��t�p�}-�&�rvȃ_x�Vv5�k_��j�3]X���ζhO0/��a����4vE��CHD2s2!+nȯ#0��8�>/Z��:���rqޑ����&�g��\�``������,I���������fI���-{!�)���m�+8˨��}�fW][��AhU+t.@C��Z%��eë����_���zIQ�&3<8NZa3Q�u-��JƤA,I��,��Ŭ�?_��Ɗ�x5�mD8+3>b:mӄݸ07&W��轀%o�	aW���-C�e%ܞk�U��DM]��w9�4u&�N��`PdY��볙�X侞�������Š$��;5�y�����Ψ&���t�z�1�<��wzB�Qg��1*�����BPv+S�^f�0t��9Μ8��`^�ق��A�KK��U����JˢO[̝H	��n!X.y0�Q6}�'Gr9<���^��8O�ܑ d6���F/MC�^O��(f��<d%Nʶ�DNX$���b��(X���R#Ȁ��u�9q�h� I��S�]'�e@�ַ�Y�J�н �}q&�VŘs�6��� ma�faseAj(>��L�(�R�#���[�m.#29��d6�ڌ�����L+f�X x���'�y	g>L�V!�չm��&��������uHy��W�_�iC׎�z���	$�x�qb���Y(S'�(|B�s')JX �3#�d}./F�Ԓ�ƥ~�OP�$���dVM���za=5��`U�;�����	he�gj�䱤�c+
U��\d�,���{�8�{����8t���Јj !R���Mv��u��)�#�L#$��l�1��n�Y&���K�t"٨x��]T��#�PS�`�sG�Q}�Jd�`ҙ���#�
��!��l���>G��I��lA�N�i���
K�	�%L�D��5�"�~�,jO��mim����4;v9���r��X&G��,�|@�>�X�wb�12��Y�b)��fxq�����k��v�}aꌪ,���̊/��5c�4h����2,I��C��`��t��"@�Ue�6d'bprH��g>��[C&�0DQ�\&Q��X쓲����HT�Z��'��ucL�lz�ibg1��1
s'?c��{�/3y-�3�㥡��GcC^E�]М��FMV_�-��*Icz�f����<y���rX"��u��XP��|G?J���ݐ�x6%5Bv�qfXT�LN$a��l9f��E�(t�CA�D�K"�f �6�A�s�W�
6/�ē��bPt����/i3x6L.#Ki!M�z~9�if��2�c��9d6˪jk��!������ )ki�#2:O�w���p����G���` ָ@q\����*��8���k��N/���-Y��f���ez2�\���_�h�'cV���ꍺ�ԉ^o��#��ר�����\�4y^1
�)�铢�������_3%J����ӕ%� :z&��A B�<��w��P�kiR�1�i*��Eg�dZ�F*	�q 
�,C�E<c��2�8c�{��s7G'�;����D���t\�K�p1�&�Q��$���#=߃�Qz�8�W
��e=�� C��1H�E6p���	�i�y��*���e�����A�gK�G3�U�~��9P�'h�H�!���a�rǬ^e������ܿ^�R�r��{���x�����r�sK�my�,v��XB�Z����L&�.��s�h���0�m6�RH��r 8��.� j��rl��%_��=����=;<��s�ù� �z8�U��W-q��rJ����dԬk\�]2����2�!\(0��%b���ܙ���c����E[0ݺΛ�톳&�2��8Pp�87��"|`<xR�?������&�CTEQ�F�Ѳ$D�e7��1/Jd^�,֬l���z&�1����N�a*`�K�;����	�q��ό��U���՘#��`>�.Q�#��&�5V�|�X��_P�o��",D��b(9�IH`�m��Rop[��{]��Abb������O�"O^���؇����kG�m<�G9��<�Y���x��s���	�����;��h,�Om�;q��X�-��/���0��� M|>�G��.L����{W�Y���&���3�[�p5C�O(oD�H�
b�"QEj�d@���2?��R�v�܂D�J<7�`.7IRr�}���?��Y6fC�KɜP_��;��
�E��9�[�4D���ap��aK�a]�0Jx��ɔ~�����[$�d<��G�P4<�
(oP�,2��;�/��M�����Ë�`��c�`��`=�e$�(�9/�[B��No�s֐�:]]��T:M=gv����4�I�D�vf6]���UJsgqd$C� X�\��i1-\��3��\��?,L�����eή9YFD���>� �T1���W��P��O>��dL�腮'u� ���b����gĦ��<�+
��a2�??=�� �_��,�j+�����/
K`gpO�HΙ38���J}mC����� ����X���B��
`��f��ﬣ%"a��˺[은 �#��֙��)�m��H���N���ZM�1�u�$�@+��ܠ�;Y1�60}����y�E��E�}�6���ɲ�����g��`SF�vG�Y�1�dI�`8s��1?/܎��uE'S^S����(��.f#nQ,�F�q����HF�V��uM:k;R뮐�wr>�Ç����LVA�� >e�hd�d�y��ND���Y{� ���<�;�zW����ޠ�h4�;03p�MhEJ�
)�I+�>IO������8+R��"�\��1�C `��о�|�2׻s6����jP�}���4�]uﹿ��/��/�g�*�Z\U7f����h<���"f����A�7�(��s�6�7���|w�-٫J�T��z|�2�ј�6�{��1��jҤ�ٶ���wQ�u��� �[|&��Ǥ<[uH=옂(?;Y ڋ�s�vX���x�����<�p&���V���.3vL(��+6�T?��N:;��� ���4���Q.i|A�jks�nU^�'vܷ�#���U3��1!��nE�ohxX�NS�-�Q�)�j���� Z��k�s�I���_��o�7X����T���t-I�^�Piʡ�G2'\b?����������-Ck�TI'˳�����^u�C�m�g�+gTE�����1��C�W��5i���D,��ED}Q$��]��>���a�L&U��c�S8p�&��\��F����t,�s�����+�hk�����0!.��{6��2sh~N��x�#�؅I���HK��q�&���:�w������=U����_�����)_��e��{�`!V�N���~�	"C�������3��5WM��`tϩ�![<kP��ª���8~1������x��̚EF�⋞����ݗ���D4��E������0�t��jC?M��-����`�3����wlT*�q���?�Mi�w�߷*L�$�H��Ϥ�o�fz�� ��|%��`�Z�*x�JE��4�4ĭ�oeZ�e�Dh����E0�jU��L
MO�q���8���-Z$<����F9�Q��^����@C`R�ːD�l�#{T_A���R#�Pv��l���Ϣ��R�)�sNKp5 �tH���ʐ3�ݪWQ�.������O�M�>4eXm
���X"A�=&�ܯxy�ݲf�����ѩ��k Q�V8-]Z[V"�(���n)��� ��\/�%O:0c��ن5R;��|�3x̚&U������6o[�1-U�Q�:!��DY|��\ߠ�$���#�|�Ё¾�s�	cP��5f��9;a���$r�H�`�[�Զ6�)��ݮ��ҕ����Vx��D ������:C�����*�Q����n��h�N�K����v��Pq��?ݗ�70�K���ىEc	�fI�G���+�l1�ؗ:ך�-�Ոޒw�w$�1Z�`1���f���S�TǢ��mX9e�9O�ӡ��0M�pDK2i���{7{LK��+c���uu�X@fl��1��Y�֖WV�\Y�" ����yT�$�Z
�|t]�j��s3���FL����gٽuw�Wq��p3�(��%01�	��l"�/����@�o���ٗ�b끶�<�>����7�O3��f��W�LFin��w-Gݥ/�se�t��7�����F��}�{��z�TM����F����(0hR��ܭ�ETח�Y�0 K�9q�%���lJ�s��z�L%�%<O����'V8��7:��t�f�*!����U/p6\?��O�����{h���"��vi6��I&#���m����>'ϯ����5&����}_{������}��p��%MM�#�9r*�����D{����L�����s;Q_�&�	2Xm*apv��y䊣J}������M�_7���?���a�d���1�<��k�*-q��<jeS~u,��j��Q����i�Y�������H$x�}a_s��)D����؟]|��"�����Nˬ7m�2mI�ݠ}']�b#O@E�^ҘV�_����|�y��I,F[aj�=GO4M��˞��Yed`�󌏍a W���,��� V\���~�����Vm+�7ϣF)��?���Fij���b�*�bϻ�:�TgU��J�I�9��HSV��(�Fg%���ظ+�D�4�6�FMLd�nw�U����W�Z0IsX�Ġ<�ʘ	��a$V��%�#6�
��vϜ��\�lM����I2n�v�(e�1T����^ew�@�S��܁���Gڦd�ӞJ�fT��e5�g��D����5�Ѩ�x�x��.�iX�֪�&��ꌭ�j+���d���&r�<���ymߡ}���Y6��г䨼���VVqI?�Ρ��K��.�kx,P��l.x���c�􉶁�I)�֦�I6-:8�G��(��̗���eD�������	��B�`9}�3�j�9#/�7t&�FHD �@y��g�c�_�}��]e$�G�-���]g��wыQ�����T�������F:���f"4�a=Mx��Q�\�,��%��3y��1#4���֗�UǥI�{�:�-�|6����Lq]^�����B��<R5��C��O���E`�bKWBԓ������ͣ�nN���L]JZ�U"i<"N�R��{�~�g�H��ދ?�+����?=�W�V�^7�.겆�b��&ͷ�zs�ä=��}��U,I�"�P�S��{*������6���+<��jE0�/����b��Ѭ��(�K���J_��'\ ���9�9���YW��@�F�Q�FO�8��"�D��։րXp�����E}B=S�k��n�ف�[ѿ�NQ�F�1Ҫj�ҥ�tt��@.���;�M�~r��G��g'L����$���4��W�=�Fbp����ęp�{�ZA�\V�듢����*�.�0P�K����n��X?q�A��;O3���Gҷ�x�Cp������U��avɮ��]h������f����/��a�UN	l=q
�)�Xe�մ�/�J�x�9�X��bes�B����~��§�����#Z�2�A����̪ _7���+�-��~���ku���VC�F������<r.�[�q�&�[��l#�'u�ۡ)��4hl����&�QX#n��T����E�2��R�_M<��HX���� �49{�}�A�X�?3��w-S�`�����w��'���R܍���%�zZ��q=WN���E���藟��aҐ���qI����V����y�S:{ք�t=�jTeuG1����p<�F!�\�,��'0&w+?R�;����:��
\�@�ٰT:�z��(��2�=W5�����L��z-a>_�x:�ei���Pή�l�K�ѻX��f��~:=�*j�|;D���^#쯳��p��y�0��b`��P{gj/��Nݷ��ҙ���i�f)���9�W���y����D���d3yT�=GڛF�Bzp��E�b�m�6��@�-=>���}(N�!78&g#�ͥܺtղ ��fk�9F��vC^��ҍ"Ј.4!���L��7��z�����I�{�sz6�Ni��	��%C,��y�qm}ё,�|r����pU���u{���)�'$�7z����іg�1C0eQ�+���|�Aa�\ZUF�NCG~�Ķ���\�I�9�j�Xa�JG���τ��	��Y�r�R
$lFό�����DgW�F[ �4QBivc���#%����,o`wm]�C��s�ʂti��uv�u�m5���r^^U@j���Fy[^+�Lֳ�:)�W�!���ق؜��IV�Ic��Y�'�/�B.�X��4J�ىQ>�
�u�<XOۙr�&���˷�Y�EF�I�Q�j�]���������懊�0�P!�R�蓀�l�[e��k �ڮ��|!g�Yl����A�7��Z];�6�%]��SM� y��U��6��T��б����M���T������]�}�{��{',�ɂ���V�r�}�/�v�Tܢ��x;Ƃ�`BZ;��d���$�`�	��� *,�}M�91��DT>��z���̾�
��C��
q�|zT��̡uu�I�kh�GM�{�Ҿ�����|�����ϡ;~���/��]5���@ⱴ���W�}l��{΀;�M4���a����Y�lC*�O����F��z~���~q$��)j�g�� 5��joN�n�*�jIm�%�Fi�\�(M:��c!b&��Ž��6�vjA#�hݢ*��a��p��	��G�.jv��0t�ϩ$:�E0�{����R�)�ϞYnJ�k�^�2�fi�4Sw.Qh�����d7Nբ��� �aw�v�W����~�F�,ԵW���N!)�V*_D�˲'9@Q���^�"@Д��5��u�L~د(+�ƍ��Dcz���sK/R�r	��g�FE���qT���I���s˦�$�ܞ�'P ��3����5l��88+�۳�F�P{崿���g��
�&�B�OBEZ�5��$ؠ�z�C����ͬ2�V��{�3�g�(�ZU�ΤK���85��ЈU��VQY_G]��\25xI�O�[-�M�D�����ē�N��X��v�xŦ( T��vIf�c�.�������(�x{I�h�}|�E`w�C�y9_������Nf]��[���E*�[1��m럕ge�	�e��
�Dttɤ��k�Ib��Vo*��m4tҡ�Ʃ�+�t	��*�QOz���V,�L�aht\�(�R_+cgmY���U��YX��z�h����Z��Xl�����D�(h�C��'�O�L��%���T���m�p�j�r�۳�^4�xχƜ�Z�\�����B�<����AM��J�$��2���^���g91�wV\�Q����:i��⮒��̪s�T�ʂg�1/�|�g�Ie����������A�c��Vu3�n�aU��*��L�z(��aВ��k��7��ƣ���%oT� �Y��=�hj2!T�(����>�QW��'t��}'vC:r_=�ym�O��N�1�Ĩ�|gK)�J9�8w���1cX%�d�������ӣ���t�dN}�V`yZ��Z)���&O�G�ݲ�6�5�~����^G�6�3�~��y�7^֤�C�֌�aځD��x���>���Cij��ܫ.�;�X�y�woku^�em�EO+������{�:�O��<7��̆���<�R+��,�ݦ��U@���Nv��o.A����;�1U����-G>;j���OB#��{�]��)���)��N�V���
"R��J⼣ͺi	4k�0���l6��y��է�~Z@JlaV��$P��ԖXM�[H�l#��&+�Q��&��H��Um�@���C��pF���[GjpCӓ�������f����:�V����,1F����,e"ϓ����I3&�vT	��}�뻻h�zo�LH��XKS�m���3�L�>�dOp9�X���մ|F&7H��Q��%�cE߁@c� }
�g�+���^��*�S ��*뵅��<��d�d�XmU�Po7��f.(�s��
�wn��O�CՄ|��0��K�@��a�_������O/i�8)k�܂��R	��zo��[�~��2>㘝�-��[DB�����Ͻ���ss��� ����Ͳ���;��צh_�`�T�h�[D=�������E~�U1#�z�g����W->a1�wI}M�S���򺚈���@{v�908����g�e`�11
����αEt�h�I�D���Z����V���|��?�Y7J��t(��ir�7����FU!˦G���$t��=����"U���Y�.Rm��J�{`�2���xY�6��_R��G���q��P��Z˚�U�'f+,���|� 2�w�����!3*�]¸�Ѝ�����_e}W����R��X!����������*���0SD�TT�]ÿR�87���u]��{
�4�lo�w6����/��U�Y\�ͮ�����}
4��6	Ъ�%B7�ՍJ�Q��@ʢ��f)ZRkU���*��j�X�;he;u^߽g�4�Y6���w�R�f0�:�*�����#���d�}��L��ytu\�*�{�nA-,���b�i�g ^O������YW��ڧ�0����Z�U�� �����l�`��w��Q��]F��m8v�WS�� ���B썳��q1qrl�������Uo�������O������wڼ.�{�)OjE���n�U�MV�W ���)�F}-Q���W`���:Z�c����Qzݒn���g��˩���䙴�ٯ.���9O�14C����e��mV��"��@��+�1�b�4�R��i�KgTBVrt�6ՠTM\�����ެr�����V1�\��j��=�^�_1��V(�P>Sfl��QdG�J0B9�Jy;�khll��;7H�g�=��B�G�{֘qq�OM>���t/��{�����M]g�g�لM�[ܵs�Y����	q����wo�(��%�۳A�aU�]R6�#@�6��h��6��V�Bd��C=�lj ׯ���Y���H9������/׳��{@?�f�Z�L�ˆ��ʀ�I��F؄���O3�|��I_��G���q�OO�08��Ny�6�˫r����^�3Q��6T�=�}3מ��=�6���+��X�o#��ֲN�����2�����˳�D��ց�=�2`Hz.�nPT���U1���Aw��y���ޑ�拿>r�2r�W�QՁ�!
���#�W�Ă���������$uf��N��4	���3?0<��#��ss}u	�3T��,����P�g|j�oߖ�sM����r^�w�Rj[I=�	�ő)��89#�}�������
6�uZ�kr�L������X����P�C����Z����@;2]����9����.	(i�%�I�@�qʋۘ,	�=��0R�]��"jً��4s�.V������:��w��D!�����SO>�3"Wi��)y?�N(�~�J��e�?z~��&�d-�Y�c˲��r�=�0:��>�ƪئz]����~�P�������uL�̠,�����:�f`TnV�d�DrN�.
c��O
�������A�#Z��������`I*C7�0[B^���6�c%�%�����"R�!�c4�2u�Tʨ�=�5K�L��ح��Y�d��}��M���z����]B�űʤ�G��s�(jq��ۢƈf�c�����Z) ����T����{w�2��4N�O�:���~v�S\>�v�5�$�����%ĆvP�Vq��	<z�$>:W��7.���i���[�=�8���S�V��mln��00fs�;fl��of��w�*�d��#8z���ΰ�j�֎�W�Wĸq��pi�\ީ���s���1m�01BS��v�(0�WT��8|F��3Y�u�{]���
�e�ڕ�F-������}�
�8p�]����#��?���-�2��VZ_?�z@�Q��s�Q����½_�w��_{@���=K.�T��j��fCk�w�U7A+���5�G��f6���4��S(��Bn�4�s��h|A���kf���|�����:�U�FcR"g�������4n#t�r<�7�JG�����s�>��	8�O�D?���t�S]��yz���TE}]�J�������TDT�>�.4EL��2��(�r�Ig�b�P]��S����Rӂ�j�^�Ϝ���s}�p{�(~7�gw��_��u;M�x^�Ҳߌ���P�B�ט@��U��b1=7���?i�O��ҹpA�wn�|i?������ҀA�`�f���e�̀��1��6�GB!�Q�+˾1�G��8�?]SL٫:EJ�nL�'�T$]C6i>�5�ku�3�"�}���v�ڤjul����Uڙפ�t�yJR�[��X�,&AE�f�t-&]Bƀ5^,V���(wv�QPQ_`Q�陈es�d/9�=�6�zr]��zA����#%fw'<*dvU5�ì�Ό2pZ�p��۩%V�cv�����/��{�Ú)rGz�:Z�i�,&��!�U5�����	�O�����y\�rMqhN��ᾞV'xOI���@0<��O�ט�c(J���%1����w�qn
�f�
��DM"�q�*��*b!���i��2�֚�Y�Aum��m���}�ix�4�@?��$�.��X�*U:�8
	�O&a2�6���}��&�{s���R�4F��Q�ȝ�y�:[D���U����=ve�Q;��˘��es��cx����%��s��pI�����;��s1�Kx�����JA[�8��% "���͛X\���#��hkd|S����_~M)�a7���k�2�$��5r����K����{-���`��	\7RQS�'W(��s�ЪpG7���)��벾@�M�	烜b3A����JS#4/v�)-��*f�.٢�@���Z���h��ȟ�
���j��s}Bp�7�`��M���.�tȾ������?�j�_}�Uܼye	(�?���z
G�Ř V|��K�����ZY�s$E���O�^���~��{X����w��U�;>Ɛ�>x
�>������A����;������3&���3G��br&(JS��Z@N�ݮlBu[��K�-��5�C�^g ]��ʨ�k�զ�E�Ih��X�0W���Ĕ)�Q�G[7=�[#s�dU@g�j,c�
�xM�-��/����(���0j�q1�1W����	�KB���Mr)سng~~���Ӳ�L>��~���p��q�����uI��#��#��DQ֟@���^�S��ĉ�ǰ,�s�:�668=��gp��Cr�C&m���x��w0  ?���ʧW�nk�ƞ�b�~=Ҩ�fƑ��ـ���L�78Bg��+���M�`��~���"�/�|C&��f�odL������WIۛ����\2ڃ�):f�U�\�������(�V �۲5��\Ә�9S��k�7�o$[�g����m�Ua��=����]a��<GZ�{WW�$7Ы�˥c� ��ˈIL�{���my�	s�������%��e�M����[����lZ�ɪ����3'�����bGb���/���Erh�>�����XZ��!j�&�y�<��}z�\X��Ʈ�M~���5��)���#�R��c�]��2"xoV�ľ����kQ�7b��E�
�̛B<4�i����NO�W[#G��x�����fC���-��	�w�%/=���opy%���sA�o��w�ȁ��u�Yq3���b�>���ʰ�h�+ߕ\l?pb������ϋ�`�֨:�/��� � ���Խ�Ц��%R8L�'����)��6Oc��C!5Q6x�XT��FimR�rټ.<�i����%��'��IIf3��� @G�𔺧��Ҳ^b��L��6ڜ�b� �b	RP��%�G�;Q~fLup�� �lH<��gF#���a��"�+)�ڮg^������RQ�����/I��?�@���ێ�=`ޕ��q-B���,	b8��O� kW.ц��V�Z����%�;%�PI.��rM��ʓf@�^��)*�6Ǡ\@JT����<��ɠ�Կ����&}�+W9랩>%<S��@�����fr�w�)M��Oi_'ߛ�u�rf$R�W6��@�z���K�l-UǺ���2Y�
�$3�X��L�����3U% �P��	>�}SB��y�\o�V	�ziBk��������nC�;:���{���J`vn��@�Ͳ*Rʜ3�8[��#r�2�翳�(�5�hxh�usV��q�g&091��
+++�֚Z�⨃\��5�$`�9^ZZR�lS�w��U��� �L�F�l��!���ĩ���Q��F���1.�%�P�G��d���&�O^�d�s�J7�YELF��^#�+�Ϥ��O��©ǖ �5�'xnYa�9�_X�	�hO0���@G�L\#���.�uv/t*��L���CV���O<���ܾ}Gi�H��Υ�8�6�K%�>}��η���a��}rW�$�I���&��S�>�U���5ܹ��?τ�HiǎÆE�լ�7��M\>���<�������αyZ�$8K
Lq�(�n>/�#@C�������<̴{�,Jr^��*�U~�=&�Q@�R9&J�l"�!�Ob�	0:�:(�Iʞ,K�q[�HowS+Z%!շ�0O��8a�P�)���H�ǋ"����;��8��K���%�H{Z֗���nk�� �f�(��In>v<�k��.Z�Q�zzNr���r�$��l��H𴽦t+U�L��}�ߏ��y ?�ַ��AO��D��}�̵����\��Ω"mS�_U�iu}�nE� !����G����S��H6K�"K�@�ףp'SPM?��S�9�,mqy�I���5,߹m67�gM�ej��}ߦj�V�_�A��C�4���� ].�b��e���̇��Q�[��\��V��Օu\��c	��䜈�������-��;�.)H�v�#�/IP�Ő�C&�)?���'�Ҹ%������ԛ�o�}[�DFL��>��O�������-5#6�k�����ʤ��{&R���ؤ&��*��ϊ�weFx��"vv|� ���@z@@;��SbmV���sIݽ`Ԁ`\�|�*�hjז���q*_[�FJ��n%<�-Bzry]�2j�WV��:��3��J H5�h��3�{"ӈ0�U�&J�F���S��;>�po��&���Xe*�|�$FŞ��>Ԫx��q���Ыo!��?q��MBe���n��O^��{o���[�O�w�q�I�Q�%q��<��n�����Ȑ��&�H�f`>&��3��r��VWX�9�������s�2E�O-˿/_���Z�5�?8�o&�$4�8��&tl��K�Q�M�)�"v�C�^$��9>��kG�3*���?TY�k�.*� �1{��F�j����^�� *����o��1��!]͡�����+bUv��yK��`�פ<�,Y�2I�~z7?:�QyF��0%�ߒo%=���+;U$� %���k���z[�iҬr��2�Ɔe�3�V�w�Ք;Ş���q���#WHJ�j����bK���ӟ��ӧ�����Ң��"�vk��OUЮ����,�/�4�V|�4E:n��=���B�/t��=�(�C��A?t�}ת����|�tv]�J����sĔjh32�A��Yg�Y��4V7���v]Eє�J]�>� HZ�炊��x��� ��'˟�,��bD��А�7́�� E?s��� �B��-S��B8:H�g�d�c�8��i1�����U�L���?pŁa�v+5��?0WÐ���Q�L��u�ÌH�>��������v`�\��)�^�������~����`|y:,V�`��X҂���	HS��*W���G����8p>�S�� ��Ksa�魯c}��9gM/�����l2t�,U�6���2�*��E�hOD[9��(��^6%$�T���H�n��^LW�둉���_6��+N��_��_��+W��~�������(J@ˁ���SX�\� ��H	��L9Nvy������F��߮�kzb������م9,,�<)A�{ｇ7^{M3���N�(�/��
�n$aa� �1ш�\����H��'dU�-��~���K��� �CucjVN��8V�|*������Ӭ���r�� =�N�Y֚�1����b7��CSUsMݾ�z/�1�����tF�T�_�p��l��'�Q�w�$�|zC�����`g�'10T�qhqq�s@�_�t��}��*Ǣ�]���s�>�=���9	^J�\Z�3T-	hI�48��g�`d��o��7��P+�rN�ݖ�4̩$-H�)d��NQ��6AS�4�wQ��2�H��8�|d\�̨�ɬ/IqrIuqϔlm��+�-��9�L��)�%���*�D����W�.�3����]�tR�SB*m��K�#w,�v�����0*��=�Pտsq�:�DYp�
��Duҽ9u���%AP���? 6�-���-��8�'|w��1����G�o}��!|�K_���$*���=��1��o%	@Xո��O$����9�LLd�����[o�=	���o�3�����e��z�9��B̵i�B"ft|	�SS�H
d�4#������+���i����Fg��,!)Al2��'m�	�āR����h!��ɤ����;���o)	tˍ]�$�eҮZ���rHI�{�a��"�@e]�]�zalTGv��	��d�ང�Wܥx#E�="�9x�X,Z)U�hW�)8T\���&F�0L�% {U�� �����y�N��k�^,���fE��:r죑O|������,�SlTI���)L
����Y�����yX��JQ>������I&+b{7��:���I�{��~\��c�\�����G�������F;AZdF>��1Vey���a�"_U�&�~y�p���Y_��(j�{�ϥ���*f��(%w~x0��ݚ&�fĆ�Z]��M/pB0<��u�{����eu�>����d�t#����ќs���6ַ�����αW��UƢ���eT�7TX̓�,�]H�z��W��-<}_[P���� FM�}��Y��\���aʞl�ZX߸+�G���v�4���똘��x�����+:�`ff���� -gϜT:�w�}��W��[�GCȖ�18�����LPĴ��z��t�&��k�9����:��Bm,HM�ZS>������j�3�Sb7`Q	�!�&A��$�ݨ�&{���/����%��Q(L�1�zj��X�(P�{��j�	��@u�;��Ϲ���%�;��ZՕ�x���7�]l.��K�  ��IDAT/a���^:�ٟ�O>����ؐx�!�-38�}e�r�=>��&�Z|���}���{���w��>�����+c��7^GM��W~�Wp��A,/�u-K����q����g>��E��R���7��O/akcG��"���������OI�.`E���ʵ��D��^�H���<�6{�cK�/c~?i�I�O���K�]k3�a\˙���F'05;����n]��8��,�~$18"�R��N}W���k:*1Sl�Iǣ���il��Ն�B^� ����C�(�' @����J������0̹�+��u��m����hI�\%�����TvKS�o�RA��#����6���f�Jz.{c������U��>*����c��%�2ı��S�\]ï���R���ϟ@ee����y}T�w��'0"�2;P��~��U�<.t��g����(á�M=��?{�#���d��J�%�b���o	C}O�E[�15�c�ţ�6Ҳb����&��t4$��x_Z=�a�ڣ�G�YC����K'��mqB�k-���+�GU����S��;��e��U��Auw��}.�����1����]��%���h��B�ۇ_|��x�o�����*��6XMjV1, ��Սu��]4cm��1�M�*����l2�]k�Q@25�t��r�X-dEfW��Դ����Y\���~�=��%�H�8j���uM��/��yp谚�:�;�h�%�Y����� 2��
�(��G�g�@�w`0�=GgS�M��7���
�q٫f���*�ո�6!�$�����{�R���� �����������k;��R]��o�*f&)���Z��ũq���&&%ggzh �ܹ���9�w7t-�g��I(+ns���+���&5o��f2����=/�$3E�I��p��A���".�lDYd��kV�Ѯ�ؕ���E1��b���uNRL.Wy};�+�(W�cK>f
����JH{˨¨�sUY�z+t�V�Z�{�W�=f��`o�,c���wȾ��č���/�T]gn(�����8 Rc�� �tA
�(���~h�����;&�)��,�0t}�1��Q����:ɹˋCb�Ϗ�CY��C���4J����W��bDYy�sf]����\��%�SK����%��x���qS�~D�)	��wB�hI���,N?���) �! �7�^+e�1.{�-wrG|���x>ciaC���X]���oY��c�N�J4*� ��zt�_˷��HK̏��e�ڜ��_���SɬP=,�s;J�p`<4*x6�Ԅ������<�&Ʊr���Ef^۵m�3�'t�!(�3�n��j/\�ǳ�%iBs��v"��(��ݺr�ͮf����τشx{�w���O_�5\���M|����bN�ANli��)�Rw��wU�nmy�";M�*.����kW�V<x �by>�:�x�Á����`��'���n"?XDabqq�#��Y�k�/*-�S�5?%w8)�"�`���*`������b��7��E�F"��wI�����82#Z���j�*�&e%� �c�gz|H����c#E��MsX�s�Պ��P�"&��Bj��A2��v�Z�a���ڵ � aD��[���dS&� +����|�cBÝd{-�-y�}�i�3�p����՚H-7�J�5��t�py	���1k��9LĊ?�J�;<1���O=�8���̼�����?���?��_�*6t��׵buW����Ɉ]�ݏ�)�25���ͮ�`��.��V3ܼT*]y��� v�L���0� ��٤�!�(��_�������8r�>���}�����cg��u���y:	믆��K*VE�H.kbՓ��I�k�����Q�Tu���jF��w�Z7Ƃ�fJ�����V\�vY
Q���&�׶�W�y�Y��d"/d=��]��.�Tu�*b�j7������/6���Y\_��Z��g��U����X�{<\*⁇DVl�������8��<t�槦���n� ؐϘFbd���~�k՝�L����+	hE�<����&t^QΏe����TJ)}LM��I���3�z�	,$��gp�����Q�l�^W5Ƥ��@�+�c�SԸ�)6��m��NS7j{	l�J�%+m)p��=[����m���+P�o�������֗u�ư���L�ٛk�OY� ��T�n���>�U39�>����(�$��\R��J@,=>Q�����wΉ����_x��:Ο�>v?��_ǵ��qW�ﭻ+�@�ę�1R(⇷o`��e�u�b���1L�/1<�Y��+��B��)�����t���X�U��*�E1��)�(�xG��'v;�}h�o���<w�n޹��W.b�x	�'����[XZ/��6E���?��B��^7�>�����=��T�P���nNl��Q�Xi�Qe�P�v:�*�t���'1Xak�rw��֥9o�[ǖ|Oj�(��� U����T�}/߽��|�Q�s v�� �@lt^�eA��f.���_9'���FYb����,Y|�����c��-�Z�;o��������,Ț|����q��`��Q��2��F���$d�@�R���sD�6�x��6��kop P�3}��=��{��HRn���Y�pl����1��o�M}Y�~�c�Ә	�x��s���7��e�b6xQQ�Q��:�x�aD��%��n2f�Jl`w���^�,o�����bxdX�2F�j16��F�1�cQ���$����hy�~�̫�j����&�'v��'J��Ϻ-	�n]�k7��oS��������W�:^�ld]��-q�u	\�7V��֖�:q�(V��� |(���>���	4����2�#![ދf�_�(@b3�,%����ת&@pG�A��s*������y���k��*
��|A�d��@��f��>�/4j��v�
AK{Ir��ViR��V�F$����Q!�5_p�]��5ן�p�Ѯ��k0��R.-nr�5��!� �7��w�TI�<�<NJ0���o�\��
�A���R�=��Q�Kc�`ՠT)P.`K�/���M�`jlL>SW�L�ؔ�jSQ6�S��M��O?t#�A�-�`��+/a�Rű�'���@iqT���7��eu�ڀ�-�ѐ�Z�iR�0Hƴw��ځg�˽�Uj{�H,�*sF��><�w]���'&I���qY=��$
9�W����V�) ����㸛p��9�Y�|��j?�4z�ۑ�_�eJ�;:���0ʷ�g�N�?�qb�4��5��:0�� ���O1��0��^����^_һ�h�%��A��g�GW�"� s�F�&qR֛��L'��/�K_�"�]���Eڈ��óO?�g>���Q��Mٓ��{�/b����[L��齸s�&���Kw%Je�@8�>���l�u����a2��3xA��F�rZ���EU::_E��-&}d��9Rt�d��s��e0<8���y4�e�6��dTɒ��
s���4Y=ק��҂�B)y.=u&�~+���-�P�I��w����rA���G)X���{�#�xE{�>�qR��kH��y�}���"��<���AU�do��Xa��š��U�&ke�6��Ʉ����Vvw��_�������O(���W����ݿ�^���H	�:��)��o�=���9�y�`k[)�B:�@�̓Rǻ�z���tUH'f�`q�]m�YN#Mp�Q�D�"�JCJ!-�/�e���vyI�����&kT	W>��O<�a	������(jb&'�r�����m�֪M�do��VӒ���)�2rpV���6T�%},'���Ν�g����ǧb�fi���C��e�M�-	2L�Y�#k���-�X��ގ�zcK �E�%�o83�sEqh 9���~� ��G�⣋w�3�q��}b'7����Oq��Y�~�q���y�Eo��&>���8�|�5T�݄��@X��1�k�ǧ&��?{V`ӆ��&���zM�>z�Zk"ZF}G�l��BU�6�V����&:��MU���P��Ӳ?E�[�������fg�1R/��
�tUD��V���VL[�l���̑�̞g:���r���92H�B,-�$�����7}��H_��3���P�}�r�&�d�m�'+���a��#j�j��v$�O�~z)l�/����GԖ��� �T�����խ��+����:~����,�����3�ॗ~�}�����M;�����p��]�'r�R9��}J3s�I\&(ey��"j��H��T�H=�#TS��o�$��B��s�T����b�H1���1�>���^&��?~�Ã��g��o}]�����7Y�<gX
X����Ds_��4���B�*!��^�Ԫ���{ׂ&�l.���(Z�c8~� �����
&3��s� �cė�����_`��ij\�V1��VSH(����%q������8�c}f�&��/>�[�Zr��^|���Cd�����8�����^A"��#��O��^����3�eOEL>��cGe�<M@�rM���M�f���t8Xh�)���e���[�����#ˏ�a�v��)�+��0�`ݔ�fK|v�R��}3��g03?�}���%v�埼�s�O#7���49cVln,�L���Eb����=�#����~B�4�Y�q�
�����"�GG�Cύ
����L���$���pXb�Cbg�������:�cE�B,^����p��	H��Y����Y��cH�g�p톾�P��3�P�<��'�2P����.�;;h	(����Bh>���ġ�3jǶvvqc�6���b��d�W1Y�mh����m��&CF֑N0:m4<���W~��u,t�4�=t�4�Hjr�(�|��V����u�}֫8��5㲧��F ��s����@�a�Gqj8NB�(������G�[H�>7>�_z����C���?Rg�jc�L�T�=-���f}?�-5qĮ.b<f�`}���:⬍�뚊��;7ocsm�Ȥ�:X�JS�M��&?V�g�����{�v�Of���F�ر�-����|�G{��~��}\�tY���%�e���ɑ����K@�K��ZY%ŤT*�o~�"�C���_�1����b �hʯ�NM�(��7f��xSYSbk�,f����P{��?�]KN��3N�V�գ���އ����X�����0�9 Nt����01�A�
��\�����si|��hsMx�������M�p3�c��t�zՕ�}�p,-/aV.�Aq�Iq�s�v׶�9�*��=�Ҁ�~���v�g7�g�������|89�:��0>2$�Q �'�#����>�ۋ+��^�LU�ػv����_�Uy��*m�_x�L���u|�K_ґ7n���
���q�=�A��&�pQAZޯ�Ĥ��N��T-�wL����>�E}o��v��b2n�����и&8��)FG��	L��^�\U��h���8���] �l2q+!̴�i	�`;�����{&T(F�A���W{6����Ϟ� �80��꤬�}Ǐh�amks�E��;�3\�5�s�!}�t	R%I'�@�G�t�P���Qn�T�ի����q�8q�>Gyg�CC�>-�1O>�?���E�����_�n--+�8�� ^z�e�������X\���ߓϟFR�=SBV!����?ϐ���^ii�Dvq�=�j�	4���>���,+r� Q��=<Ʉ����&@���Rs`n�C%ܹqW.]��7�əu	d�B,A����0
Vh��k�A�EU�e����� �h�M�Ë/]��� �=p��<sV��7?��ﾁZ{��H�
���Zy���>yn�G��*D�w6Uu5&{R� uh �����Q�>}
?x\�w���Ǐ^zY��(�p��E������/��?�<z����>� fŎR��[rF�DF����S��9p
��!14�䮊e��Qb���s�*�Wia�8�0NO�8mdt�Iwo�Dc�f��r�X@~0���aL����g���C�bOF��>^��Eir?f��)V����������߳�~�3N@�`�g�*���E�U�U]�u��_�3�Yz�_	������ɞ�b#�����5���^��sE��*wwG.y�����8���"�g�=y�Q��A�#{~��e<������[�8v��&G�n���O�/���*g�����O�����U���c��'e_B=z���x���ͻ�­2r���s;���B�	��1S�q��4�%Yz�h�h��fΙ-﹙f����V�KY_e'�Tay��+b�:8u�����Ç��:_��	�?����y}�I_d�w��@�l�g�IM�璦]�T��pj����wU�1RH%r�Y�T�6��:9O㬠<� ��ƨ��!Z�$\6��O^����>�d޸}�fÅ�<����#�|�6V$F��C�Z���5�]��Cy�}���k[`����Um��������ۿ3ss⻞�7�&J#��H� S�(�BqjՎ�s����u����2��
�=�7B@籆�6JJ E2��Ҙ�'&G�x����ߨ-k�ncD���}�i�K�P=<R�w~�U�<#gT��7Z�7�˪���e�k:�6������OfBe{[֣�TԺ�x��Hd8�C��n��4:}�ҲG����Erq�L%5᜖�K�p���n�vy�^�(:/�����9��ǈ�?�����W�V��/''�Ŕ���- ��=4��Ȗ��.��f168�����~ �>����ӿĚ�)i��b��1x���NA�����Bܬ۞��v�Tq;4���^Ǉ2�8�%�)&k6%@�ԡ̕R~��7���k�P���ի��{䱳r�� ��3rG�O���z@�Ob�-�-�o�{E�T
�GT�G���CL����^QJǔq&6c}U7�k�bVb��=� ���&V�??�)q�MV�����}�l�BB}ƅ��+��!טcD��W4p]�.&{��l�\o�:����|{M�~yS�w�XBI�2Y`[ee~e��S���X�V՛�v:��%?3���ɣH��"�c��me?�'׉W2!�X��)�퍬s������������� ,���N�)^����c�F�M�S��v0�J@��Pn�VT�ce:������@^)�l���Yq<q�����W�����-�%r=��I_{rt�p�h�ڧFU���"�\/���6om����l���r�?y?��ѯ	���Q(�(�uFIΌ�JV�hW�h��7�l�UG+�8q,_����8  �ef��8{�a�گ�:>������\�	ܕ���K'�&���_���2����=��׮�C=,�|�Ͽ�C_{,o��3��y	2�6�8�~�h��Q�\���R:T�>�s���NԀ����%O�=��6������#a�8�7��8�Y���]\��>��n�'j��K�J0��	�9mXn�9�(�)R�"����VS{VYyn��Ρ!�.�yBEn_<����T���� px{�.��X���Uy��8u� Nʟ�inv�����9|@����<��i=ά�0���=�J�9����w����j�����#緆/�k�O���^CymC��+�䓋x���8����S�!5:�L~��)������g�(��F�hF�S�������p�E��5��:U3�:����\F�7#�Ь %`d��4�}�����$����4=+�zI�޺����P*\�Q�� �sb3��-�+&�����q���΁���iqn��fid�H�|�ܫa<��Y����;e}/iv�d1�ŨnK��I�)g���1��1�i��>�9�\n��e/g��ottϿ�sx���Ul&�I��'������ȹ�����do������)��2(�H�d��cS�q$� &{:]G?�!���Z0�P�wr�ƾ�1�3���T�j`/+mh\!���`8�(�C�@I���'����		
��{��99���� $�iy�eQ����Y���Sdpʌ�V.a�m���/�E@A���� hdF�,�5��82\Ǐ��/aJ�?���,�YlK���l/	�*�62�ٞ��P��7�h�R�*�,����&&&p����E]����0�x�	|r���jrf߿�8�^~�<�՟��&�'�}��_�KU\l�������T��;��hLbpjV nB�	A�p֌_1�	����=eJU9u.^`}�T�#%2Ƥ���|�Eq'�`�SX�vw�ܔ��d-+�:v_|�I�L�cP��W�=����Y�*�$`}�9M�mnm	ؽ*���)�sI/�w�B^I�1�a��&�=)`F��f�*�xa�bZmy�"ڞ�*��+g09+~���v���s�.������D��8[b���b�P�wE�ʶZ��#?�����?U�|D�k^l���z[GJ�$T�^S�)���Ժ ��fdH�M�{�`L�翪b'o��FgJ�5�F�a��ٓFYS�O�*7T�5J��8!=�j��ZwU`C��T�U��
��3⫟���X����?��/�����X�^ō��J�?���16���V\�J��/�<���y��jo��6�,�b���BG&�v�=��թH�4I��CClOW�҄\���w1�A^�GC��=OE������s(��,�*-g�cW2)srW�e�.���E�e�([D♒��C��'1ɦ ���ӁE�<�dU19�����2(��Y��)�g��=��)<t ���o����տ������^E�8,�7���	�bYV�9h�I�u��̋ԍf�E��jCe�AH*F5�?~?��1L�ع��w���7��$>�">]>C��0��@/ ��Ul���@�`�_����������}W/_ 9����ĳ��$��=�˯H�ǞH�o��=r�SA��W�,>��-��=v3@=p�K7Q]^E�%1$��؞S�=�sa��?�@|q( v_��sx���W^�ͫ7T�sL���XM�ɢn
���sXZ�����8�oFA���E���t�=��x O=��Vn��/�
W>8�����c�14=����*�j""4z<�LдC��A~{8�}u�l\�VM��kϺآ��8~`���r�"�q�e�+w�N��7�jR�����[���ߐ3ǭO/�������wt?�z�}\�H�]�~&6�)��m��j�-P:O�bq�k�յe쬬�;5��42��d���v��9�-���>B^>���w�^Gv@� �j����n;���ҵ6��LF��^t67����˗J춴ov\�1�ϧ�^�}j��^��	�7+��{��lHF�_yu�Ϳ�s8����/��}'���4U}�|�U$�/���Sy6��F���t�{�>������+b���R���ٶ�#��B�¤S�8
���@6
j���f#��:<��6�J=�9�����l@�R��L>��2Q�\��?�4�(�������>x��T�S����8�.�>�lj���1:7��B�� �l��f�;&��-��˳�?�pg?{���X���d����F7���I	o�n��hI�ܲ���I�BzWA6^��|�}�x�k�iv��*�na�<ַ�4XkJ�|��E\�|I{~�U��>>s�-�����5��\A��t=�.�	̴*�8��YUW5�T,�?GE��9�{HgH ��0VL!6?.�i�W/im\��y�\O?�8���/(���_���qb�a��Jj�ǲ>���f��:l�� Z����:q	����MJ�k�T�ih����i�ZB�f	�U�޺�ph �JO�-���rV�~���5�R\�#����ܮ	|��ʙ�bCr:�E9s��yֶvt�Y�6ױ[�ĥ����3ψ1�����ڳ���0 g�ǯ�M	���#(��k�k��q� ��hFx{�w5
��sQ�%�Z����=�곇t�X��'�A��i_Ed�}���:n^�"�y��=��/㙧���1���>�o�p��i�~�����J�Z� ��J�N �96C����,R9�@��I�ZG�B)�Ͱ��Ex�%�y��Y����.��i��TV�}���J�����V�HU%`i���&�}u�,�����ʇ�>,Ap��e�+E�ҕ�(2:�wjj��*�C�&�"0	���A��i���yee+wV�ؘ�����;p������$������^�ػ�P�oY�f�^�aj$��~���V�4��S����3�������}>{�~��;������UU�{C���_���px������i��_ô��o���}�go���`���7E���/m�M�hoQ�g"m� ��.��${��J΁��<v/�Rx��Q��W%�����aV��m�mk���U��DS<�.�����0�����ydJCx��S�+K��,�B[���wT�=�����)m���J�ݖ{P�3rcq?y�-	>8~�0VV״B������$%ٯv��Ǔ��Psv�U������H�Q�g���R����ĩC��[�]�8����"��R>��������6^�Kx�38����/O��U�����G��DB�`\�����gr�Kc:{�!��ݢ�rJ�R�Sq&�Ǌ� y*�5([.���oP����e	Vn,.�ݏ.���Wq�͟�}��d�0��dS�~V ]<��\��mT��_zR���ſŹO��ҧWUF���E���?t��@����6���C�k���*8��|���J�������{r���������/��/���.�H�\B3L���>-X$tlX9�+���n���21֠"%� u_�k���u�r���M��sؒx�*>�&>}y�d9�)�f'�;*������^�D�BN��eܾv]{����/�(��/����V�c*���'���6�H�~L��h�����ve[�`>����vW�=U�dm�������0����$u�6K�--�w��2.ݺ+���1O^��Vu?}C���	b��!�3Ø�.�?�����u%x^N�^�� 9�`E��Eɲ,K�����<3�Z���Ժ�[�Z{����$�<3����,Q%Q��@��@��9�~9�=��$嚪ݵ��"v�~����~��{�����Z:��^9�$O%�ߜ�Je,�����ٵ޽�=}h'���c�ŗ����3��N\�D����$3�����ʥ����%��1��R~�[HW��]8��H���|���Y@g�z�HlN���1�<U5"�=�x�s�/�W�:�����7q��S-����˳Ѕ{�<� b<�KS7�Y[zڅ�^i:�t6��[��&�&`lT�4���y�$�R�[/��D,��f�kV�gp5�Cg����2r�Mk2�#��@2hS�Z��)����,�&4�eѾ�����j��<G2��o`z�^{�u��֯���G0�;�;�����3!�-`t�6�H<~���q�Dѫ�Ԇ�޸%��E�O�҆��U��0���9v�q�%w�k���S�m��J�Z!�S���+�u�M1��ɛ#���wW���E���3o0^�:q����~��ܛ=�C�p�$ҹ"}�1�>��|�Y���*W��T��y<�Z�}�Sɵdɜ��A��B�Q@Ie�v�͘&��=�EE�"���o	I�g�1�ԟ���0�>�G���|ֲ��2�b�
�T���oMb��ĹKc���EtEPYMc`�<���.��011iI�j�[��y��d�&Y�*�
�;��'ykos9c�l��<"<��j�5����u{o��?�%�Y��mr;uX׻��]2���K�h�ٚ���d��p^�d8���r�t�c��S��
�L;�|�c���	����w��Sǎ!0�M��a`>�n����%��(7V?��hc����?I���*nN�ڌ*�	?^�KM���m&S�i�Ԧw�.�cֱu3(�-W��ޝ�̅-}�*:��Ò�q�K�cC(�p���$��O"��4-�&�{P�j8�82T3a񡿷w<d�T�d��"��X��hl�.<�*�!�	3�xN���G}�La�Pa�0i��|>~-���c�E O}^��U�1��z�7[Ua��ء�!�oGO�~���v�����q��`�u^����^������(~�ӟ��w����
^�3�������g`�䢋+	�<}.]�l�� X�J���4t�.O�%ӕ�\�,^��0�j�h,f�753��_eue��:Iy6�0�NI�Y~�<w�����Ur.Ɍ4z`��6C��*���$�v����^�8�(���1��yH5�4L0!s${�@8�v����?�$>��S$����<�0�hx�Ľ��U͋�H��m�G���[�a��Zud��Ͱ���%p9`�^����m��K��$j!wG�AL�]$ ]�3,bpd�w�|�!��./�������d��m�l�!!ނ�g��K_���!B�!��v��<�$�6��ᬡftJ&Q�ۥ��z�Ҧ3�jm>_4�4?�����G�ͭ��s�Vx���Җ1��|p���u�+E��l3��<�~�N/���S��Y�������E6Yĩ���8��Pc�����"b]!�����`[�&.��[Ǳad���!����9�(/�L�~�<���n9z~׻2�w���Sé*#k=��g$-3���"FGH�vb�Ɣe�c!�]�^~�d"�ͣ�,ÿ����Ǳ�����p+�S�`���{�"�=�����7M�%XmY�7ݞ��r�L\T�@�1�G�$�Q��)y�O�԰n�]�u����M�f,X���}�$��؅_�����X"�Q/S�/����w�'1h'P�C����.���"�&�$�U���d
����A�˸V�����нصo/��f�V���<�����xA�M���C�d0͏[��O�o0`�J�Snվ��^+g����kt�\�-�I�jr??�u�W����l<�������70;vä����'MB~�����G��"�{��7���?D�����&�9br��ۿ�������Ɨxv�5Ыʠ����3�F��j�R�P/���mݱ�[w`Qw�������0IR� (�{N�V'W�{Ps4��%��E�^�{�D2�x�N�?�w�2�k��^#���Q���8{_|�k��U�q��{��m�Vnن]�w����7p������� ;�;��ȯ;�	o[�Ϫښ&����25�,M=�&s~7)ݪ`4�<K��zTM)�UIs��y�
�|^7.��W�����8����Y��H��1|�#� p���~�C'01>�B.����o�%�{<����ۣ��l�IgS�%�»��V_��Vy[��6�ZBI#�y�������&���o������n���j��֧����3fכ���),��:W�j�9��c,�\�Gz斍2
����̡k�&f�͵Y1��#�ar���CV}�)�/�ʯ��r��k����3��s?��� ���x�Õ��Y���+WvYL�~�{SO��ej��Z���N�Ū�Nk����>2�R��C��[���k8���~�3o��b2e
���|���D<���>�,N��:��؁+ܓi�%�}ٔ	�l�}�d�g$��II�]��f�Ԝ����4����f�S�)�ߏ���阼~��3h&BR-�9�]�~��L��%b�WD�|^,��~I�_<�2�y���8;6n>YK�`\�~�sKصg��n5+zav�������ɋر{'~��~�XՇ����$���g�psf)Y���w��ݥ�7��;F0����t5�S,���{��.�sO5�m�rzk�jz�1�v%��c|���(�ϵ�X_���f�
6����)õ[�����$c��ƍ��C�{8�������;�k={���Fw4<^������?n��p�)��&�{h�w�[�n5)Bse��r(O��G:���X���;&>˸��g�@�Z�>���c�cO��c�M��%It���坶j85��cέ�|	�4�����7��@4(6|r��UL�-Za)�ۋ�-;077�o~�9d������!�]k�0%̍[�Ľ�R�ŭ��n�����l�?�Fk޷ȷ�uq��3��R�y���d��+���u����T�B�9����
��z\���&j�G}�Ï| ?��}X�����F�bIr̹)6���w����y��x��#�~�
B$Van�M[�"Hp�{�|����[��#bP�n_���^2!��}��ٴYB5Dw���is[�h~v�����᪐Lh���/��]�������s�9��(��rR�P�G�������!�|I�JV�N#��`��^q*!�r��׿�����N��n��������h�=�����*!7��2�hޞ��jv��>����ɋK�x��(Ѫ��\�,v򒕅v_W�ܵ��>�5����	��&H���8�Ç٘�L&��oÛ����/�[�cVY�	�:���$k&[��_k�q�z�-�*�eg$1U�ƀh�#�����ضy�ӷ�zz������3�91D@<qT�m���f����Z�._��/!� d��a�w�uIh��t����b"�\�@�9���$r�8�^A3^m�vsm7o�lrX��}����G����oH���޴5��b� NnpVC���;�d4�8�L�n�8�ζ�虗^�n���mV���/F;�Ͼ������XZD���-�6Wmqv'	d�uƮ��_�2
�5�x�u\8yڲa����o���1Gb�W��p��Ճ�r�,uٗ+��p+o�L&;#³XkU�e���3v��E�q>���5��f��!���)�f�9$�e��I�4_sEl�3sj5�C��;X.��|�3 �؎S���t�
ق��D�������z�l�bm%�����ɏ����Ǐ������c;�ɱKWx4T>l�jժ#}ץ�1'\'ۭ/3"y����Ү��V5W��,������H^x�����!&Ʈ"µ[�����������L�	�\<w.�5������P߽a���V�X�l���D����U���S��Uu7�{�a������$(���l���A8q�*=$��� ���
8��|a�$�|�D+���zL4����sعo7����4�H��I��q��3J`X���^{�5{����n��ډ����`g7
��c7'�	�@
�l߹7'f�&�A�"J2KШ�&�%��� _�e1�p+���>�;��.��S���*��2U��6\e>�2^{��+'_�s�z���j#>4ZG2M��N��yɐa\�E��x����q������گ�ݢ�Jsu�,���GrO�j��T��f
8'�a3���0	�����0zI0e
�d�Z��ݺ� �?� �w�c�1x��rff��k9��Y�dR��cfe�Y��tK����D�|V9��l�@b�;�������(�x���G:���/b��=x���{ɇc�8��<�ȃ����{ӈ%C���w��K���������{l�*@U8|y�:��k~����?k�h�����c�hM��N������a��{�|���]9w�rމ�$�%��T2�>�$���/�s舶��{���!�Dv2��/��g����/[���qFg�K�'���H��l1�ꪭ-4���xvj9�$1P� 0��2IA�]Gqe������d"���l��6�=�Lq_�Me�1WH/�t��v�ϦВǊh��F��Ն���q�����g/�'��u�0���y\�t	�j�=��9�~��o���q�u��q�-�d�g"�Kٜ?��W����#�Z.�5���'�%�ke���׈D���z">�koG�`{��4�Y���7��u{aHɧ�fg�J0߳T+u�㚩�&����4����ʱݦ�*�#o�Ra%�N5��H�����w�v$�	d��C�@B8��ƭ�eL�&�h��[��M�;-�y����gx�-r��\Ӷ \f_�m���%
E�%�XJ簕�� o~?پ�IBR����ŵ+���V� h����b��4Ÿ�x�
d��>�,�c���-�n��B����1!���癿�����QޞYo:nWk��S-��L܄bI����x6�o�$_��YB���Ϭ6̓�볤t��ub
a�"I��*�#��#|�c��K���V��<pj뮖�Z�Ƞݵh*�ϒ��ڻ[Gx�0v媩)t~6�=�G?�s����̉�x��$J�e���5�;5�6H��s��n�h�DmM��8z�m\�q�ح�(|6SSʓt��d�L,�}�{���4nN��ܹ+���ORP����9��9�,�c%���;va���f���p��~��g%W|R�ʎ|T��q�W��	Z����/n����Q�u�[L��x;��lM����~!�FJ4��]� @�M������]���De<��L@�Y%9�bb�����/�r9�b�zj����C��p��z�4��m?���yӀ�w��6����{�(>��EW(��T��W�L�P�UAF��~�@o��RnU� {��޵.�z͍9s�*ܤ5����:���f�5Y�>��
�\�l]%h2�+��qTù��_}|#�h}ʰ���ę�x��Gx�<�qo0v�*�\�\Q{����#j�^�Ï=��c�s3�;t'���=؏�˗�@'$ ��/�{���&k�,�U	S���q.Os��yݖ��$7h��YNY�%��j����߿��ky�dLm���k6�xl� .^8G�V��7��8����?������'����4���yrZ(:�%5��9�1�yJE���\����˥�V��ϼo�����@p��3�N���p�*��̔��(�E�ʋ��A�M�#9
z��6���𫓠���ל�V���X8v
��]8}�*z:zpkbS��f��g�޻_��'�8��;�܏^�����~�m��7O⣟��Ix�y��	>K�01���T��>����ԯh�6�3�T$Ǚ{�(X6G_+9��PI���)�0����x��Wp��I�>�8س��_�6.]��/~�K��?Y��;�D'�_6�h���gNXm��&o��LO�B"�2�빽��W҆�B�0����yɶ�����M�@:�ā�{q�\�t�!�t��}��ªg-��U��Y�k���^e@��Ԁ]���;��v�����U���A���Z�\���
����UND�n\��}d~���=����Wn����P�����Ͼ�%4
;�^{�(�c=�|de�-��,�E0\�,W B��F���'0��h���5���P�;T�<>oR�:d��&��ZY�1c�)�|v�yy��!<��&����*���\%���r.n�Fl�Α��(�|K~���E`����*	�*���-�[wL�|� ���d~W�_�����Jc+q��/"J2P��3D;;0�N#�3&�^%p_ �W�ui3>U�s�N��@�\Ħ}�p��5􎔰������#���o�:�0kuiUўy�<�(F��u|�/?��p{H>�(pO~����.�!J2�F�X�t�P�2S���Y}U>�C*��B+���j䤏߯l��E5���xW�-|b��@����&���q�E�Q��hU�^�3��W�l������݁A�[G�0N�`r|}o8���ac�3K��j�:����έRi�2p���ƥb�f��l��,�s���+X]\0�+U����w���x{6m�2�u�g㳟�.y�d���%S�hDB��"�9g	�-[��A�z��t�]���u�>=XXʠ�;d�L����2���_س�t��ͬ�	ry+�qs|��O?�F6NP4��ӌ5�>l�c/���dK���7���{��<r5�=��p�C�eu(�����\6ʣ��u?��Jb��o��5�����l�{���w��\c|H���+���/�����r߬�K� �߇����M/-�ٗ^@ li�q�%A	-�-��n���;�Us��F-A#���F�g ��n5�D�H��9\�]�;~�W~}<���}�������9D����w���y��b���ǆ�8W�y^� �{��\����X�b��1����K	D�>}A�|�.]���� �^��j[�d�C��_�W���H/.cq��t���-h����P_W@�-���5*�TN/����\�����6M�#�C��MC�%˭��W%'L�jn	�}ɜa� ��d�WE]�Es��6�]�d���r�	0��Z惡����W$�Q����{���"�����>#��k�����|�p0�5�r��9!I�b�w�?ĘY���e#_r���G!���d�j���<�3f/��l�e<+�^�i2�0�O[����1�3˘W���0>�Pw�纉��9>۠����U\>��
$Ѝp �{��c��ʹ�Y�T(���J�k^&Risfn�/���m�Iꆻ3rM�9J�"��W#�����������*�d"����^X+㪻Nb���(�YE���C��y\�t�%F������M��EZRp9ݫ��Ήw!�j�>��?�g��|����`ݦ8=�^�6���N�����>��!�a7���1<ڋ���g����Y�U]�w7y���V�&�E�J��b�d=C�����);�$�=�|ӏ�_=j�'9Bg���Ufu�Rĳ����<3���2�%���x�5��õw��x��(�̽;b��.SB*�b+s6�G�e���{|(/�����L����Xn�4�5�i�`�_f�-/�1��`O�mc�5����N����w��{������[,�� �����I�`�&}�'ݲi�}�~�_����"�����d ��/��kGl�q|yղ4V�⇟��4g�}���� �y���W�3U�z�f�a�JM�5�gQK�q�t��\��}س};�LS�SpsA2�K��FD�6�DN�`�}�`��38�l�D�5�I���N��B0�9H��P�S�X_8r�J��n�І��7��0�@�z��|�z�-�k���q�a�<䲕F[e5跅P�4���h�|L�Rsf�ș�|[su��k6���~���:�m��!����8��$8Ҭ,ê	��2��i�f#&������"J����SUƪ*.�Y�rܻ�KSh���,:6�M�����Z��R1`��YX8��d���44��g�'x����oRdPM���Y�hT�n.U-�$"����E��<x�lۉwN�1�ps|��i��ۅ��lٺ�	�N��Y?�ͫW��?ƶ;��p���q���I����A��}���Zck6W��	[ P� �
���5T�2`�֬
��X���	�$Sn[���
/ ?�o�{:�s����_��̤\��Pr]��>y��"4m�����S�U�%j�Peɰu	��G�s[%P��$
-m�.�*�eC�V�O�*�����䦆�Rހ������s����4?�m��Z�š����$V�~:�Z{XI��$k$~s�eˎ>�@^�$K�+H�b�8��<���عs7Q�G5�Fr�~�c��."��k}���k�j�`���_����&<s��$#�\�t�ic$�s�=-�wՑs��V���FBA�.��#��u��4PTf��5YR������IJr$o�wF��ݚ7�ud�6ǒ_��rc��5I�v�z ��@E�)H,�H\��G�����c�.�7�V��Z#$Wu�a^�%s)�m/�:;\s^8rZ޾�k	��� �V�'��\멑�����G-���B	��_���Kr_4��!>�߫/�D���D7�����~�l�e�3�cI����K?�1^�u����b���*��M����|G���*V]=g|>�[i��L$-����*�ukȯ٬ʈ��ȷO$�wSQ�,���s�����Ao���/g5�n�W� `Li��0�t���\+�|�
T&��٤"^�S��YZpm��>g$A��A���ɘ��/ʵҸ
���D~�u3GS�Jw���;H��n��{�]WFBK\��C_W'<|�	��Z0��>�ˈ�� I2�%)ڵ}���k�V���7�̙3�Ar!�-�6�e�W_z�|�[7nZkC���>����\��+!�lك����W/]���%�/���8W�����w6����M2iY�2f���bE7��uU]�5����)drU�jn����q���Y͛�w*^6��d�|�:�xw��6�B�A�Q�,�,ɔ�A���s��,�%)�$�m<��#���Z����� �!IrS&ّ�[Pu�%/�"�C3sV��0��t�x�q��T	|!�I�������λ�����/�ǿ�f,p�bq�g����W��b����g�����XC&�ǅ�W������+!�7\����)K�	Hv�3yWD�$�;?q���"�ً�*�$?�5���y��n��H���Bu/��Ik�6>�2K�1���X�B�!_�ղ���p��
(g�N	��\53>k��,fʩ[1�洽�9���ccd��`��l�ʍ�y)��:{�1�q3�Hp���c-������f;�Q4�yx�$nK�eKJF�3L�[�?Խ!�?zz5�g=��N��x�m�x���Q�5ܽ{�%���%�qTɔ��'u7�f���p5�Т�f��9x�ǯ��7�Y��g���)Ȓ<SJ�����o:�)�4�ZI�1���Igʍ��W�Q�\S�����Ǒ\S/�<Ƥ�KSsR����[� ��Q���Sq���*����\g���<�9t�u�w�Q���@S��Y,-�ۙ�"Hɩ4�N��d4�M��@e���$1K��J=�I�,��bZ.�)S�CQ��.�Vz�W����~��:�������$ֈY����'��D@+J����(�X
��۰�Gwta3�Ә��i���Yb��;?���,����Y+�x4���<��^�S�f{������j _P[Q�Zq�>�A�!V�8o�`-
� k:���x� Y�r��b��
&���s$�F�����zG��}v�
�X�������}��ւ�¡j�k�1��R��l�M|l����K��u]d6D�`[AZ2�J6�ٛ�0l�3F����<97/�����9��'����<c�%h����.	iZU��EW*�N�C�l9n�F�c4M��[}<@~����z�̱��ͦa��E2�@�u�D��W#�Q�A_SF#��g0����Lԇh��0R��~��l�=���eą۰y���O]��T��*����8����� ie��|]e"e7>35���7����jy��FVլ�_�.]� kzc�����Y�[�"M��K���nؼkv;d�bs�t	�m�����oO=*|���5S���u}��wm��#ߺ�=6@��'��r�?��o�3����u���
���T�SUE�ە�2�j�1���I�P�/��]5g��o�>58Y~�����n���ܥ�M7FG�l���)��i]����>0���v����l�Q^ ʂ�s�� ��=�}�rp��5sQ�|�7,��ٹ���a�A2�+$��$6�}�l��4�ı��bqj
a�*\Q��h���G�U~Z��O�u1�����6�{eC��N�d�%��>�r�R$�aI�Q��'����g�t�5U)��̩�8{��5�k���-36?7ms�LJȵQP��DO ��^O�w�q|���"��.)K����̰����3��D�i���/"���m~������� �W�{����X9s{z��>f�3�ю6����v\!Ϥ3��ꎪ/�S˼xVlX���W��������hb��)&S�1LL�o���$�c����ϲƋ�;�"�d\�7{�{��v\Ak6Y�k�p!h�y|�f��_�b.!���
8�rI�v�#��zi���1A����o�&�y{��$����d�j�F�8#]��W���b1�Gc����]�Xz���s��B �aƠ&��d�r	�SeEkɆ�	���8���3��x1+���p�*w��gs8E���%~�'q���O2��s�� 'I#��[ݟ3�����:;������;=1n�F��|�g��WЖȚ�����VIh��J�2�l��I�Tt��,֧���}�q�e��R-Z�Zby�z]�A�? DM���i���K%���0��$�m�3<O��T��<��aZ�^I�ik��EZ�;�ڹO5;/��C�ֶv���ԝ9Q��"�s����܋��!�߰Ѫ��I&]��n��0��lH�$�٠߃4��L�TA?s��I�kO��C�K7��ƑWQ,h^d�fU��v#����z���{_f%Y3S�vmo=NP)�NSH�	��-3�e�o����ls�:Jl����{��\1c��<��"D�T5Q��/Y� �!����x��~���h���Bq.�,��T�s�f��F2�vw�cr�Z�8�d��<���z����3�7S�(ɟ�*Ϊ�z�>�5!�8DB]��慢=7P�B��\�����5WP&Z��	���jK߀c!lp��5x�[Pf�Sձ�q+2��֎�Yh"���׿�m#����*��q�|��5crɛ5oxM#	rL-�q��U��!L�/cab
����,��	gܪ�+6�\���,���&�~�Kx����.��T��+ ����c�>[�.�ň��I�#EH[� �#A�%oWBG���cs��c!1�4�J�qY������Z)!&@ٴ�X�D�\���h�$�/�%�-�y��xD@����I��^.N�V
�ln�9���������zO�H����yׯþ}L:���Q]��?���i��ܵ��'�>��.��jqj�t�wW��˝���ZHϗ#BU���ʡ��0��,��Dd�y�>\>���I�x�]|/�}:�jב��z��p��kv��ػ}��o���<f�f,a�����%}�������w*�e���[1�B��Kʱ��q�%��#��h�\�����
~���4F�H�����E���c.؎|TgR�JrėZ��{[��e���,�����V �jm񚣬L�D��� E�z�݌�*�ȱ\�o��mؽs:x�gW������Y�&I�&�T2@	�Z��u����}����"
�Ib�B�2�� WjZ2ES��pG��q��
.�tԆկ�����jw��=Y��|��|��͏�;I��7ɭfh��_c����~�c��Dt-����ڞLƌ����ʩ<�a��;��7̭u-%�QcL��>n(	��8��!_w�dQ�N�2����\�(ZD��1�����4[���K��廎Q�〮�&[�����Uz�Z�j�LeIN����s6h�?/���"±n�_w�����' 9GM+U��ɒ������4�6�Ve%g�l+��iNC"�8�[�P�&@P*���J����TU�/g�`{:�l�FY;�ǧ&qau��!�x�m�Ϯ�E!	�Dܔ��λ���#o��ɳ�t��Z"yE;HB�p��{~��XNߚ��V�����s�0AP��|�z+]�,~.�BH![���@69#qQo��s���z�\FuA�ZUD�z��L���s�0������$�JK�װ�8gk�1+v��z�u�"e	�,l����m��6����He3F�%O1���`�h|E8��W&J�,w��Hs����R0W_����ոY.{xх��<\�N�Qgض5N��۰m���/���_S�h(�/��W/�ov�U�/ �F�A�b��|Vr����D&?��^��Lf2�Sa0�祬����(I��F�$�Jr_���6���X�F��ܠD�	P��^dlT"����bRÚc��ҡ�i��>s|�d�bZ9(�K�����YU=���,�d/����^��&��JR���J���F�ыd�&���R�[�;�^i�w�A��zC�{��W��첮2B�i�Luu����]I����q,��H6����h��_�u�&׿���\#�]'�����bߡ;,y�/�mf�*���U�~
�/D�7�ŕ�5�5K0�Mq=��I��&@Q�[dH��U�;�.�q������Pƚ�S�Q^|���L�j�3�QbH{��E�dN�3UF��]֔�4Y����ϟ��sF��.�x���
I �I�_��*!���UE��ܕ���FC��D��I#�Ngڼp}�e�a��V&�q�y�^���~�錑M�&7W/��hW��NrF�3��wܼ������9�����Mg�g�����s�����k8?;�9����%%��}�ӒG��(d���X�e����o���D
i�)"jܸ����+\�@���əd�/����Q�`�w�è\{�<���h���߼4g������6��zXq]���%�U$2KH&���D�.��Ld��H�����f��m�㪏�qU��X�x�k�%
`
�;գ0�I?��WU�,+����=�6T�1Mn���9����8�x����=w܉];�X���7	Z�c��(z�^l\?l|/��#{�Gv�Ξ�������k����)���I�a�t'k�����(�lټ���H�z���$�M%��ν-&.���^Pq\g��6��j�i����{��#��,�<6��;�|�⁉�M�ǽUu����5���O�Ϯ��9�����B2nj%
5?LD��s��/ XmA/��b&g�I�Tq�H	�[}����,��F�E��l����]T��L��岑?I����]��u\�yG�!+Oi���M[����صg�=c�?w��;on���o�G�x��Ώ#/I(�ե<�޵�F��{,��bܰ�ΐ���P^��e|�G���d0����3��:�y�(˅ѥ89�$1"���,42����q��
|6�a ��c���*�%)o���X�&�'9�WL+��H����!aw�uɭ��\Abn�d�w��Y ц)�gA3C��<�t��Y���{)�)�^T%��Xn��u�A8��/չQg��f��(O�IV�Q���E�GZ�]��P�Z��9,���<��C�d��4��������L�1�ۅx2��;v������?O\�B�{"E�֔����6�6	ݡ"�Ns�#�U�I�����
��7lGm5���a�w�b�T&}���	����hC�	�ԓ�mT.��D�_�UV%�VKHc�bG��,�J���{�web↩f��g�U���U�\�a
k���˹4¯&�O@�Ԉ���ē)L�]m��I�T(�F�(�"�$�
<�~�J	���%�}^���-.�*���"���п��rfP7�0c���v��ݛ�ھ���Ɔ�޳3��;IoLN���Ï���}��9m�6)�"��C&����P��8���r�֟�>V�㑀�I�c}�'Q�������,u���fr���r�Y�B�Lu��Ū���3>�_�1�K̼i��o��`/�Kx�巐]]Fo�+�$���c�t��,6�dt��ʳe��b������df3��
?�So!�ՙ[���6Z�����$1����O��O���Kn7�޳��������X�ZMB@�	���@�,fqs�R��l@6�3��u��4��-�A�a�KtE+3d��<�ʀ(�%8
�r���]=��D��>73�H��mU�ʤS�|� h����Y����OQ�9�o]�*Kk�e򘋧�4,���$f�X��or���Dk�i�-���}T�'��=+�(��`�)�b��BU��/�	)S�&Xe/�I��@��A�|���T��ڀ^U?���b�f�A�Df��Iy)��۴.�����<HA9=��7T땜Z�y�z��_�!ic9���-�!��#/�h�e�e7�4���H�d��Vi,,�l�j0����Л7l���("�d�+�1�D���q	�Ν���-^^2 ���ŋ�����XR��4�_�u˹4��u|�p�$k8wἓ]�^�3fS	ܼv37',�$�<{��R�U*O�$XA,��؞�Lՙ��7�w%�N��j���@��C^�f���z��#ᩦ�Lީ�����
x��V-������p%�BU��U�u��PR�^��3U��5����׭�j�	�:�3g299���԰�̝�d=!��^�{�1%\7�l:��q`��ػs���kW.�S��R�}�>���6�N�u�N����9�g��>�I�|Kv��^�����%LO�X��FA��yF����;���ueŞ����o�P�"�|�j&.E�!�!���J�!�T����4�<,t:w�i
]�>�.N���� ���XA����	&ق#�񪥓���,�W���H���%�<�$D���=��`=�Z��F��"�:�]��e�[{X�	ҕ�S%����N��!�P�����*�}�g��T���5�f�#��$'%Kzƒ�۷�1��I$�|��e���K�q����'>�$.����X�Zɇ�[-g�<����)P��?���k�����e�*���Z��HW�z�	/_8gҰ</>�Y��[l���zJ��]S}�$�J�l}�7D�Ve ��Y��Md_.�<��EԗV�e�����Y��\��\��U����)d3�$$q�ޜe�]�lJ�*B���<ј%>"Q륩��c�#�-;�{RoH6�,��6Չ��h���~L�-@b� &���������*�6���.=������aLe��س��/��z������^��P9�>3MIZ��d5U��w[lUf��1d�(���A����5�_�9lGG�fƯ#+9��*�^��Jg(�)�"�=<� �T�"�-�Z���r�&�������B$��S�f��t���x�$��g�y�.�.���q� uyn��%�=�;HfK�����j��oKE&Sܫ>>7�<wԩB�܎�z��k��&�F��J=c�VDUM��c�������W5�_�$P0 �OP���h�G�ߒu>t��I�����~t>p���~W���|�����+7�B�5h��P��2a%�&k�#(����Qn��u��{X�$A��k��qv!N|R�d��WՋ���<��kUJ�7ܦ`q�&��ߣ�Y��Y�ȟ�Rd�����;6�`�u��y�4�}a�*M^:���4r`�
pO��L!�8w"εbd��,����H%1qk���*c{�[	�I�Z��Fs���M��kI�5�O	�	�N@r�z���%��I�*'oU1���-OaR�	��X��}[[�$z1l߱�Μ��/���}O=�!�}��̞�����.�����Y��H���Ss���wYeL~�c�af'���4��n�A�ᗋI"�Z�˒�fլ�G�X�����k��xy�k��x��?�~����/A��
�oڈ��I�zu�VW���~�����ALLMc��:��޳aV�ֈ��ཕ^^��w�]��c�����r.����^�QmX�2fNO``�0B�|jf3ߛ���tڼ�����q������}�<�ۘؚ����*+�V�$�}�XMW�k[3�,�ή��,�~�(.�s
O<x���CgXDT�"RHH��qe2TB��i0�R�q�Tu�W-� ����5�rG�a�����`���B|-�EV+L����DV�U�e0����Uˁ�1P�<��ڦ�����G���޽s���t�,����/��bo����@��Y|Vs~e��ػw�ݷ���x�i���Y��x��Y$SwIiT�������?����<�}�A���Y|��3~��Ж�DS��.�z�����)��7lN�@��M�B+�g��&��˓h� �������2I��	�kW�%�䅤"@��%]9�,�u�ڷ�T��jߪ$Md���Ī9ڕ�ꗓ�Cò�s�+<<��a��1�m��(��1FB')��]�҉^{�(N��h�qeOU���h.��*�z��6I])�'�%��:;��NܴG�4�����=͐�x����I. @U��ȩt/�`k��&�i�͡��R&��\���8.z_j�&aS3kHs��i8���r�pz��ԭ��4+��9�	���%�n�~;��h-���.?�DeWU�y�F�,ˬj����o}϶�{qם���Y�����w��7���c�9${رy�w��yxV40��G�˺��do�Fr������!���+�5O��ۍ�Xq#gP��J%�㏩�Y�g+ʤkWېq���3ɲN~g� �*�r�U����]T24(T�������"��O@#��;=g5�<dVlX��oJ�H�n�2Zg�3ײVd��i���ty)s���q%$A,��fb!�Q�q�˗��~�z��v��X�E�X�s�T�y�=N��|�<g�d���݋'�d1����^,�đ)�q���Ft�Lw�؇��/,}�2��r>T?�dC���h������g��A�@�Y��`O�IGff��WU-%d�XeF}���)�wt��F=�<X��lzͲ���ɸ�]WM�8/�$�ۖ��]uzK���$?!YI7[�C^��*�k��l�砆�~2�f��f�g����"��N��<�u'y��R��E	�0J�+�&�O{{̞S�����>9]�R�&�4M�������n����]�ì��]�܇}�o}ےH�z��$���Y��{�|�qܺu�R�$;� ͹���,;s>-��=��\���6�V���K�e&ky�7]�>�7>#���Ar��U�%�S���h
�D��9�
I4	J���y�� �\�~�yv��EP$�1{��M~�����
m �8�����2ޒTgז�\X@.)�����4����g��\:K�&{1 ��k���*i(����6��n�ϪC�@��iL��S@&�J�d��-�+�P)o�4��j8����`u����5ޤ#����c�D���� ���������bL/��#����;�q��8f�\e��Z7��ۜ*�r����Jƚz�һf"��~k�A�s�������ևs��ik�����ZUY�_��S"S3���%?�za�F54��Vܨ#:����ON����x���x{�/<�<�2�j�!��j8��X��1���3�<[!?�l݄m�6����\/ޅ%}�8�]�l��"���Ht�.~����y#�OyG��x(c�hg�{��.@���=����z��`�vp�Cg��w����"xJEy�����/�ac$?�û����8����~<�������<<�_��ϛ�ӟ�����1#i���E��
r�,�͉��b%o�T�H�9WRN�:cR� Ҏ�z�	.y^")D���r���0��Z(�8S�(�J�#@_�9���"��~�[2���C�����5:��o.��h�gD+X��Ȧ-\� V�'���D#�D8�!�zw�q�z�4�O}�7�'095�g��]�29�W��
�:�(Jm�Բͯ�#��T%�+�<{��;�
j `�s­�)�#���W*	�՚�h�jcQ��� sa�2�y;	��p���4nܼ���>�%�1�n߉��g7cOG/6m��;?b�습{;3c���ιr��a=��i����9Uv��D�ye��� �d��i������G��yw��Dg�����m&�XA��~��-۷[�W_��]�p��=��_�(���_���=�Ņy�Nv:�1�� 21�(�݋;IK٤Uwm����ص	|�?�����.\�5��kW���~��Y�8�1)K���{���k�}��*| ��Rp���h�T3*�����?�kڌq�f��j�18ϝ
��]����"c¶m��ܔ<\
�B����ږ$�T?`$�`�b�
��[DId%�(j�|�����������J|i���&#����ly
n�E�R��XH/�b%���{���O>�Q� Ų��[GF��>�������ayn�$���s(?�X����{�ud?����c�F��t�6�܂��~�zο��H��h�n|1����E�QW�?��qȟ��Z��OT��!h>;�������{-�<�d�JMP*=��ʌE'}���u�V����J��;���>�2�l��� z�.T�JAa]��.�$<̠�ȃ�	��̜�Ȼ���p��E��6>q'Ϝ�J#�ߑ��IZjjЕ�+`:u�ԙ�Y#d�������Ћ�[J %,H���-��IZ��kCh�Y�g"�g3�?��T�����)�����f/�L��<�X'7:�[h�Z�IM��*�[�*����A�'eE��S����3"��Q�i�^6��2n32YP�N�$�6n�n�:I�iv�M{#}�e�$�U���++�&ke^5�VV�"�����x�s�X o���#|̜_��e�<��G1?;e��[�|�4FG�ᩏ~o��
�_�b'pn=7A�ɇ���f��v�ko7��u�&39����[&U�#8�ʌ�{U��9`�z�}���M��q�X�����$]�Ɲ�D�-lr�Z>�5�Te�YfN�2L� �R!�R�/�\a�ϛ��zg���-���p�ߓ�f-��s�֐y��=U�5�Yr���i�@���QI�4�XRA����ۻ&�?�)���\:i�@�jѪ�n�\B@���`��_�>�p�}\Yz�/?����/���S<O��E��x'N�m������q��⭣gH�Vm��:����DD]	�N>�`K�ժ6�w;M�f�� �D�98�l:k�ʭ>gP��?_Wok���jT�O��ΛM|ћ��²1Wo�ˌ�ʈ�u�Tu��HJŮͣ�+<.�k^����q��ƺͮ��tm�̪�	�wc�dutx����e�V�/]B&��Fp9��4O�i�@��ۚ'��.����V�@��������g��E�3w(+�u&c��6IF`U�d+��=�;8���_���	��qσb/���#x�����MH���lF�J�,��2P¡����pDd$�W�9�^^��d��岦�������3<���۪ruŞ��bFL}�r��:�I��2����J1jк�����ES"�I��G��{h��FO4�C��Ͻ���s�L^����53(ٰ�z���rK�\�:;�m�&�ܽ����s�ӿ2�����_���8�Aݚ)��*j�f\��&��4�h!1py�V-���p�@�d�n��h��z��X�� �@�A�I4,8�/L c����æ�\���rK��	�ӫ�\\��>�~��~���������c$�n�*�(h#������������u�T2�����Sn��F��B	���((Y�m��h,�Ǒ����9����b�L"$T��+��C>���`�νؾg���l�bQ�ؼ	�$J|���q�^ɭ`�Z#>d�ĳ)��*���g�����F~e�k܌}���=���/��[G�����^]Bh`،zį�	 /X\�<Y2�RCg�@;C����J�I	��X�A�dcx�j({�`//��f���_Z#6��=��~��t��m�$�3��>���6�E��/�,�>y��ZL�&�MI�ռ� aT����K�5缩z�'@��[�0��>h�o �@����E|��Ym8��ٱ9xLw^����1)��\Dbe	�5;voÿ����[FHn��^DO؅G<���|���'���q#���jo�~�WP�/��я=��߃�Ͽh�����o�~<��gL��������
<�~���[�(#s������N�����c����o-����l�P�����9��{P3):*�4��,z�}�	U���|˶mև(	�];��_�,�V����119��m��F��}*�z��`�}/��kI%�M�N�9�z��Qu�Ѱ9���)���}f��8]3y��ܝ�fL����݋�N��n�槭wZI�}{��33�S＃Օe�f|?�m+>��������ן��'gf4
H{��I	�z.m��B
?~�;���{�@�Ջ����>��c����wF�"$b�s�ش{�ͪm���y�*@��T�y���0�_Ӫ���P&EWI=#���}hܗ�e�|�+t��捐�����aǖ�6.dp�ߒ�7��p�x�ޮ^s��I"���^�H�b��>�Ìٛ���l��R*a"�����VŘLÙ�d�ʆ�j�H��֮�:OM���n���~�r6N|������O?����x�x�0.Ncמ���/}
�?v�S<�ܚ��M��ie�;�o݀�G��M1q��[XZXF(�q�y�!|�`ff��^FQ�1Ć6�#s��O�fu�!�M���@���2m�n�2�PE�&��qo���2PU�ɬ�M�}	�	t�R���vUM'�g&ZԚ����s7���i3�D*[�E.�<�9�y	��u+�pp�>ڻ�����1� �m�?�V��l��$fM�J��{��;�]�nX�*���0yIrT�����JV��^v�N?H�FX5�՟'Ҧ�0ɓ,6��k=u�\�]mVfV�P�!�.9�I{��:<���غc;�]C�7�\�I�,n�ঢ়����!��O���� ���%hߴa�J�1�iԗVW05=e���B�R��0b<�!/��ih+߳O��	�:����i�>��$Y`�zU|~s�SB�	q��pg�U�t��T&r��Fy��X4��^>�W����4�� �C��|����%��[�@r����I�����_�1� @��5r�ktF�ه"jf����*c�^ ���I	��~�ڬ�BU)�%�9��zM��U�cɞ�㶹n��3�H/?�׏�}� �n�䬬.b���7'p��e^��c$i��6_ò��Ēɥj��A�6�ݵ}$�6�U��9O�=�k~s����w2eP����s.�4����%]D4A/?cņ�J�(7RU��N]��r�l6�>l�!�^_�Q��~9]0"h�6ɜ���,;X�d����	�4V�����-�`u�@���-;M) Yl�RtF~p�wuD���$"�J���^?��L��CN�aڼQTB�w���s>�c��lePm�C��|����rH�̋<�7X@���{�؍���-��%��p�cN��ő�_�k�4�d��m�>33�E��}��F�q��I*6���c=I��{��W����~�����5�]F:��s]$n�<ԑ_*h=}��IB��T���hS%F#j��
Z%!�s��h�{ç�
:xFLZZ(�r�k�=\��mʴ�Pj>���X������3s��q��	�e��9��*L^ǽQf5Q�^�9�C}�$����gX����3�E���H�蓚@���U5W�*O;c�����UB�ϧw�f3$���%�9x�ܰ~�
͢L������O}�����~�?!Y�w�zԃ�KϘ���`p���-�"��.���.�O�����ן��䬝�*�r��m��4�
?�*��j������v�(�C[ �v�1 kf���rU�,�9d���:�!�8#J�n3A��vo)� ��s�x�����U�[�@}��_6�����y���g��m{���k�̠,_pO���R�$qo�Y�Io@�����Q!�ΨY����H���*�g�CAO��EҤ�)��i)�t�JVိ����v���J��<��a��XP┱vz_����a����_��w?�ыh�(�d_<����bv�Z�GG�G7"E"��o3�V��!��a{^�=X\s#�����zG�����Ԕ���x�������M��pk��I>_Ű�7U29�}@�CG<»�gh�m6�����v�8F�j�����:x�A|��Gm<A�`��Mx��K��/�>���g~�X�B�'Pi�5/駋�cξ�eo\�y�	~�����aH��Nq7��HQ�V˖ey�e;�t:v/q�]�N�����J�T{&�T�i�N�Nƶlm�Q")q�w� ���{x�~�����T'���
��-�r�w���w8R�U��eb!R���b>���rwM�a�f�8�0�������,#GvQِ�u��)��e`,�w>�R�O�^|�<������'1:<���}�م���������~�?�����I,������b&��ా�nlټgϟ���Ƭ܁��N\[r��%|�K_Ƌ�}o��.��F�[������A��8����R�:�<��~����U���\g�	k4gQ�aE~���b��=��x��997K8s�,n����5��fr&�U}��&g�)�>�ݫp��'���������z��W��~�\����3Q�_Pi)3�	���6�jNݠ���J�Ќ-����.�+|?d���R��_����ɒ�]G��V	��{<1<���Ƽ�>Ri'�15|[���/[p^7^��$�]�h� ��3K�[�A	0|�y��'`�jkmV�х�M��ڗ��m��᭏N�9M�ה�D?K�/��+R6]���y�Q��{�0!�����tG�>��,�şU5�6#˒bۨ��ù����?1֖�9UG����3��f	d�̧�̤ �)VUpu���{���"��n�z(8��>eW�`��1P~ǧ�c�OW�۫XE$#�U���=�v�PW}?LR��neՌY!���G��x����7��+/c��u�b��~xL�b����+�m����������Ȟdf�}���b��h��q}��-�S���kȖ\<��cؼ����ĵ��x�M�vF�ne�->�����]Q�z��"P�+�#|5���fD��c���M�>.�@.UP*�&�*��WJ^$�~;R=�Hр�8t�~��LՑ2�$�ffe��Mb����Ŋ ��.��Ԥ���Ϡ�c�V��n�۠R��))1 k�k�(>�{63 +f�*{�O��TJ���e^v�5������(����O���La�x���d�8�Kb�ZA���߷O>�V��ylۆ�[��?sZ��J�����K���T�B���h���|�{@��dS�f�3�<�\e�Лb�o�-БT��D^~F*��j�lo��B�Eձ� ִ4ql���L��<�GL��u����a45'd�ڣ �Z �<��&�/=7-�{JT��/�v�ٍ�{�mL������1#"�T��$>��� N�F͜U:B	�t�V�l;��$f\ A�</����/���.�<ư�q��:���d�5�M�A�J��'�|[w�0��⼂�׬�z ���Iq���څE�Q��O�aql߶/<�Z����� =�e�l|��ś�L�KNUE9����H7�R�C��[`@��r��˒�N$�zO�)m�^�"� ��b%U͒Q4�����Ra&y��}Vژ����mM�6l߲E~��N�2ǎ�^T�g��vq$R�#,�Ӟ2����z��.s��/n�J"�*�\�6�mZ��|Ѯ4���`��~��r��!1a/��`�)g�5!�3�rǩrWȊ���(��9�[�nCF�4��JcU������|�Y9O~����3ɠ<��,[���ss�t�t᱃)e9����F������H
x��O��������W����U�H���Ύ�S)����BVA��������r�ęe�{�bQ��H��AP~����+��FL�v��g�-h�ŀ���2�֮�g^���l.��������7�������_G:�ŕ[��7��P(=.i��ѠFU�Τ
l��'v/���H�痠���4(+ս�y��bY�3c_�v�#j[漒*#�$琊���͈M���蠯��)v$��WoJ���2�#�av{������7���G:ǩ�0�������W���V�c���v�
��\ú����� ��w��/�~�����Pe.��Ź�MX�n&8/��5`I�'�[��/TV����~�:F���L{.*�A�<�PL�њ���_��oi2��W����
�\�p._3#.����o�y?�y�)�y�!�����vJ�҇'�X�	Uy�X���D�fR�;[I0T_�j�Շ%��Uf*�-��DtP3�W��J|fCc@�L�9
I�"G&�*Ş�U�,�ި��(�Z��%���=�˔��3�iC?�ܿ�����ӟ�T��Ӝ�x�����K_���"�8�F�%��u o5G�l��+�p+^y�8�"b8�:�0��;��~uw�cx|�Q,��њ`�|Ylu@�a�����byP����w��?�[���2�W5�|*��Q-
�hn�T!�ř)U7�r�F<���:~ᝣں��ܮw����Ki|�0qg �||�V��s\M��mh�����*�Ոq��5"�b!Z�/heO�Ј�vH3�Zʐ�ݪx �6�2��(0�i�����J��:YI�^����%�"0���@ ���Iď���$��3fO���_</~����T4�E>hK�@���oh/NC�`�T�k_��x'��/j�8�c!�(�~��Sx��'Ŀݧ��d<��� ��H'`�ة��5�M����:ŧZ;�4���,k�csK7ľ/P�X|�d��օ��EG�������թ=�,b,��e��q���hm�و�7�h�B&'`��#�_̠��E��rE��
bw����Ӿ��h}@��YV^���j��L��?S֒��j���H�A���r�k�ddI�k�j9�v���5:|G�b?֬�Ǖ�1<�QLS���R0�5�"���rh��k�8;����ڎ3�r������wJ0�6�;øu�~�k���;7�G��D:�����[��Zb�c���'���ȉo�Z�
����ҥ�sgT���cM���o������F���oڌ��##~���[w�m�{'�`Y����*|�-
�ZZ�G�G�Q|^[�&�S[0�����(��*�S'�4�؀�Ҷ�
��z�6�̌tG�Z�.�M�������iAu���h�� $|�`�B1/�;���rY�FWį�"���8�Ʀ�����ۂ�8?16�����`hd���6ɺ�����i�/)6�a�݆��	���ϑ�7���G�Q╫W�h���kO=�G�n���i��v�bF1_�����5/���O0v}���x���7��ϭ�☿I����g�V�+[��E�l�yd�-�c�2 �����7��[�a��0����X�B��1�C���8��T�,��B�0g<�Ȑb������,�\�d+��;�y�3�KiI S�@9�~#�����7��M ��ڔ��{�w?sj�B�8�Gi��5�����z(�7�0���Q�B_r����>��o~S�ڂ ��� hfbB�䃏?�z��8pp7I8S&O��tJ�x���'��g�Tja���K�0*���w���ѩi�s%�l�M�鳌�!gܱw�с��iE� 5É�������ug&顎7Ӑ�L*H^<wZ��U�B|S"���@����WUɼ���U5걧��/^{�N�Uj���U�K�_�u Zr���Z�'B
�c����o)@c#��,���YU^$��λ��eg�O/��.0�C�Ɩ�9v�~�Sx��}�y��U�J�&��*�O?�$FF�0#��'������ٌT-�}��_՞��ǎ��ހ\��.��n�W���x@@���>���1N�Zc	Ce`�N�U@�p0����Z�c&���C����9U���;ǌ� 5�{��� .j0Y@9��.]tVj"�L�X'br6���`��~���7�������G�?�����/@j'�߸���"�mPQ=�ff!�Ul� WO��g��,���C�l�h�+�fi	YMUP��θ�HHKg��F��(6o݌[��sU���*���. �S�["W�ؽ�~y��q��U���M�񜂥�K__��C'&jعu;����O�sܾ}��zz����p��y�;wŨ��f-��4ҫ)��s�d�
�<�FTb`dP�RY��Lj�ˎ�-�פ�d�R:�*!�9hG4�}��q���C�$0(w}��}���'@��n����(h�*Nk��!�)�i��儃��VG�oHjrK��]�=��+��r@U9}z��p޺�dkU�}�~e�T���yP�d*�Q�d���Y�Oɖڷ�-��WxJ@in]m���H�ouz7���O=��~$wU�cyI�B�{b �������Y���~x��:B�ϼ�Yj8w�O�w��b�s���h��d��cڒp��	t
p̋m�@�	���nU=&��=)�m]h� c1��s5�?���A�~F���V��f�r׬�U�4<:��;��o�����kEL�e�h��o�η�����6�.><}E{69K��%��I�綒��R����A�� n~�8{��暙Æ/`���j�o���F �QQ�9jd+�#��X�!��}gN|����'���نL>���=���_gN߲,wI��r��v6+�, k��Ӂ�����9ʉIH���/~���!�僣)6x���RȦ�꼹D4���/W|<ߗ-��sخp֛`&�t���`^�	g�RE�o�f-SE�X2�Y��  �,�22�rՏ�<'�`����*�޺~O<��|�!��1	~�28"���]��o��mQ|�{?��\Z�WR�?�xFs�*d(�����tt��V��Լ�Lk�fy{���\�G
��:G|0YF	���Bʫ���	�nIP����k�@ќ&���˸z����5�"b�J���]��-��m-���4Qa�;AGk�|�]���n�ƿ����������+8� Q�Q�/��Bږ;>=���Ol��V��6	��z�}�g��#r���޽�93⟆$h$y��aug+�v����0/6�;�����2.\��\�(�+�[?&�R�S�=�	y��Z�/~���6L4�]]O��`Z[���C�\�i��+�x�'#�Q3=k��ﱇ��T1X�}�l'��Jo��]	S�sZE�G|:˲��c3M��|��3:�c�V��R�Y-Hp!�;O��� Z�]d�Ⱦ��s��Z�-�]��Z?������_�ھ�h,2+g�CW��)�ܑ��[�b�j7����k���Zl�S��t�W,#$6r�-(�k���؉����K�$�}���X+����Q	���*�z�
F'��Ͳ�§Xd~�������"�_��@1��"x%�=٤VS�/�4<�!e���n)	����ql^���w��䯸��C���9؆�J'����l-�3�-�P���.`jt
�M����J�i	��Z��ٍ���k�mqt÷�yB�<�{���M����x�³bG��~��ف`���y�p����b;KK�������>�l�H�������c�{bD�*��wݕ������+S���S�3J�ŷ<�� ��+`�?��MF�*S�3s1(we��t�)���Ҫ|�i9��#ߟ�2�����A��W���u��)%��+�H(?��q�ɧ��َm������Qյ��}:*��,�e�n��^�����jdi�]3닥���k"i�l���?iV�5�E���A���d��)V1jz���� �r��[{������W�!%@���j�ԩ�^խ�ȏ|T�/�ho�vE�E'��n�,	8�-�~ݺu���Ż￧N���]���G��Wo�N�
Kլ��&����:(��֨8YR)�6���w��ӿ�Yc:�NS}�dx�<P	xZ��.caf���IyM����s�_�	�V���'ǌ����yl?p_z�E̥%xJ�i�6�V
9�l�$�P��Q=1��$<i�zɜ�=[)��gFX���-����	4(fj�Q�aA���6·��!%�lJ'���E��1�O?���O����
{YS@�s��X*Tp�b('��֬��]{v*%��:_�ү�O<���p�0q�(z`���k�~����ub� *8g%|nj-�m�ŋz�+5|b�#���ਬ��[4��Jg$й��z=�hM� _rp{p�>�I|���$����KP�5x��Gq�C��k����[J�*7G;��b2���ϻo�$�&�c�Qϼ�4g���_�k�X�!���<{�XIG%��>�^٠,稊9�2�ّ��0?��U��I/����Μ����ғBª#����=]ݪ8��ڊ��.��&�'��'�վ����:d��wΝ>�NW��=Sq1*AGQ��� �0{�fmٰKKY�M.�2���WE�PLm���P�{|����`�aq��N[�U�_���$���}��������|����#�:0�D�*����Cյ
�������kr�ȺGH��;�Z!��m>P��-C�U�<��8:�sU�_��x�l���:*�W ���?ǲ�!��U���G� �U�|��簡�_aL���ֿ��o�>���#T�&��ݴ��AR69�ի%&ʘ�єlFF�����f2�,��پ	����dE1[B8�P*ۜ=��}|��La��xt�nq���66��/}o�uǎ��ؾ��X%v-�0���;��@����ϱe�:����p[����7�������M�w}xZG��&56>'`uJ��2n����s�]��38u���A��U^cLi�u�Ί�r�q�N͋��e>�j��JL:��ٶ�{�<�IH���4:"�V�*E���4��U	��1�<�
��Ҳoܺ.�{Ll�#��oDE��b�T��`ʀ��-�cTVf�+�F��PvG6�Q�7��^xA��q�}���s�����U�0�ֳ��Ճ��l��䄎�y��=H<������7p��MM�bI4���#�om3�\J�0|EA��������8t�&�{���e9"A�쪑§}(���qg
3?zYlj���.]_ބ��{2Y-'�+-Uk�`�i��]�X�jkR<�/u�����	z�"��^Q�W�x�u䉫*�5�d��e�s���'��[�]��̙3Jg�t��`�&���踯���֍LFOK`7��H��+����t&eF��y����_�|Q��/~�Z}ֳ¾|2G�)�AeX⏨pN[Ї���-?�"VT>8r\@%R�$���V��
)���oX�Ͻ�4bWʂ?mI|�ė��	�I�;*~��{Ͻ�H��1B�pL��E"R�)���>��>Y�������Jv��a��ku<�>έyl1K��/�PۀJĚ`aɕ������l`P>59�Y��3Dx���-�OY"A�`�~#"G�x��������rr��Ki$�?��\��`�?"AVOOr���d.~�E�ǎ![u12|�d����l�b`L�<�9:�W��^�j��u�����E|p�j/Pm7�؄xG'�E4g��J>;2�@.����i���Q����3��B����������-,!.����,�J�b��dTn����r�bz�]�t؊^	<,nbt��?o�.�<�h���^���&���^�;ʐ������pܯŉ��n|�3/j���hG�����3�~O
�e�b�mr~GǦ�>�l��`�q<�/|�s��f�%�S�?�z�7A7+kp�ֈ�fPO2�R��@�poT|�w-/I���/q/e���Ӹ�I�/�:��o1jJ���ʣz���A^6�+�*MR�M�D�Tik�0(є�ٮ���R(�̪�X��**�C`9��P�7�A��fr��JCs�Q��A���x�d�ȨRذy���t����<:{����:ï����i�q���-�`�ly��5��]�0}����ڄ��]9u
`/@ql�G�/h?�G�U�tP��P����*3���-�ŉр�>}J�Rh�;��}��o��:�����8;$���G���	I��P��ϊ�\���~c;�{����}xA�rW��EBg��9]���f���V2>:�
_��l޼^wV�����ؗ������<%�׬���w`����9d�z�m|���#!�gP���!�8��n�����O}FB�3��$e������y{�����u^Eín�\:������0 �s�V}�Y%�����Uk�'�5�pD3<i9o��Z�����^���>9=��g��tĎ��X�I�,�o�`�*�o��*��%1+Ɵ�˟���5~���\)�[6n�`$�)��J�3���0�*���~|��)\5�ݻ��Ħp��c�t�&�;�}3b�Y1Lg�*�R��ކ��?���naˎ���������n��ٳh��aﮝ8q�82����1�;*�q��&����x��Y����j�*��3lo>)����}�[{�[c��wQN�p9f/��٭0�z�*=��* ���y�P��� 2%����R*��"ucL�ņv�_��̡�}`홻us cc�ړpF����Bj	������SO�ܹ��R�@Q%x�o���oƢ��W��ޔh��_�
�����k���>�c�� �=}O���ڋ�޽|&�	4j%�O�}M��/=���"��n�OȖ�������+l�ҏ�۷�"5;�B��M���r�^󐬕8o9Cf�C@{�X1�!��R�������z#�ƚ^���Y�;�9X8ޝ�;à0�	�g� ��U�Q��e���A��� ��K�x��=J'��LN�#ρ�d��(�s�&��*%#��^Xĵ�W���^���~$V�y�bo���s���PF� �$�>��JEc\?�RU��&����ױ{�V���ط� N�8'�'gV�=�ЅFyΒ����/~�	<�{7�Ůoݽ㩌�r�Ld����]7�3��Ɩ46u�W�{��ʨ��&F@M"�����Al��޽Jz=QV��:z��'�����;&�XI��CjD�c�أ���J��.g����3���/v���w�w�Q@aH>G$vuw���
r��GFtTP��%��r��u����۔}��c� ���y�lވ�_`�s<l�E�[�{����P8��1���ص�������|��1}�5#n�o�rM�e͖H�Öu�X�Ո.��>zP��bU����Z�z��+���8&�<`_F��C��ؒ�&R�*4��j��8�,�U� �~}��_A�ǂA��"2�N)`��$�站�R�w+F���\2�d-}��L�R�`�٧w��sW7�o�z���VƋX%���]��6�{�vm?Μ:�[��g�P^�|���~U���ۇի����19�B�믾���Oj0�`�QQ�r���`;@�+ۧ�7��EQ����0���%�_�{鲇�#��>���;W�s���M�%�gEY�b�)ΕNQM׈����K��n����a��!�dU��L�qu$�N�%�SU�=�t�gx���Z+���ͼd%��m�>d{m<�Zm��b/�g��\���h�;P�b���yo[�O�졌Hp�e�&�)ϫ�K��bKKX�~���e��g?Ӏ��5>6�m!--I<*�����������q�ޛ��.���[�`V0Ck�U��8j'�x��GI��u�����n|����ﵷ>�� \K=��Ɯy�D�|ys���}��ө�$ �f:W6v�md��o�)榌�{��PS#��2Ο��*��D�m�I0�+{a�w��������*o�j^!��[�2[lXm��f����a�����Qi;�8�H0��><����s�{����m�����}-v�ީ#?�ɂ�3����q�#���w�}<��CxH>._����/H,�e�z�<W9�M��\�&~?�P��n��!9ߤ�VU��$�H��|�]��ǽ^{�����ؿVR���e�P�G�,�1,����,O%��]�
P���.n@d�jJ����J�cEk횵��cR���gP�d��=���`h	-�8�$��~`���}p�=J���G�\�rM�2niU���Ȃ�� ��P�q��P�oۀE������G���]/�`q�[(�Т�9��(�uc���%���0�8����N,J������ԘP^�O~�ctx�KxZ hgg�^z>���A�-�qU��z�"ZZ�b�0<<�����={wk�}Tֆs�6oߥY2Ε�rƔ @�{�53Fg�E5�̪ц���b�%A��-�(�Б�g�1�b�%e5W�B��	]��D���=,A��;��q��Si����LK��Jx���$T=��r����C8{������$EV���Z�"PW�TZʿ��m<��n���8��aY�j�]��U��^"�4�\�1�P;^Q��~'�!*�kq~N������-g9.�+�w�zqq�pL�U�dI��ޞ.�d�Y�gEkzjZ3�<�T����Yxm]f��Gye�vD֜j�� 
6�S�P��8�^|���I�r�e�����ęK����fD�;ũ
p�`0�N)�|��g�o�v I7�J �ʯޅ%� ��Cok��lefvB9������r=�Nk���ݣ��g�mx�h��5k]ϴ�  ��b��B��^�O�ǖ���Q��O:��1{� �ٶ����(��崢]����ĉ�Ꞇ����/Uq���Mz�H1��e�Zݕ{�07�������GF��С�p�ã�x�_.+����`�I�%�S�3�8� H�{����o|�+ص}� �&�;{AA�?Ѥ�_����/��bqf��i�\�������_F-X����12t]�[T%�`��Fv~m=�T�Ip����8��ܼu�p⑄:֚ ^��� V]w�z��n�-�H�A���^�WS޹�7�z+u�kf�c:,�R��gQ���`��ʂ���6&��GjY���q�~۶mF\@��˗��G�1=ΰ��[��w�_�e����}��d"����~����V�|*��+H �<�(A4��(�4�K����8��A;�2<>��$җ*�P�,AFV�=�'N�ƏԈ�~�%�w'���95��|��X�Q�BD+*\�Bfe�Ȉ]��P!�$��+N��EU��3������q�(�{����׿r��տ�*��ʊY����	�/X:���U(R�X�g�>����Z.a���>���/��D|��-�Q�{t��I�M�c�47���XC��ޥ	L#�o���t�ǰ���8��!N�UT�\�(�q�oЯ�
�ز�hY@�ܓ@�R����"殈e9WT��5Đ�V��w��L^Fj1���ֵ#7.`||��9�b	�É�,���p�"�ȧ3(f�d�h_E���v�:���{?�`�@1-�JH�x��|�,�EbF��^^�V(����&�QZf�):��A$��ʾp�*����_{9���[�F�T�="v��׆ٹi����3����������5V�����D[Alꪮ�{����GJ)f��--	|���#��Tȋ�|L���BQ8r�9�)�Ф~��7��o~��
ȧ3iL-�`��)=-x0��٢��xSR&F�G����$�U������g��4���
({僣#�J�VV�"a�̖��랊���,����c�{�����{�:���t4�g�TU9Y���̦r���5�_��,�L��`F�UG2!�Z�/�b�r�.g��֎T�R8�sX	��[�7�?N�eV�]����s���7P��U~����lkzz5aq��YD�7�H]�\[V 9@u>l[�-�3E��-�ɻ�ۚ�P_l E҂�_G��D�b^ޏ���6�x�`�W;���q���8S���"X�$}�ْ�����UK�����-���N=鹨��޲`�$�m#<��� �K��5/IF�
{�%��`�#�_a���)�<���s��~��bdxkV�ª�LM��߉����O�]�+�3s8~��
$19.�gΞ�w��x��G4I��Z«���9��������|<x�b3�\�/ֆƶ�h�X��5�(�S�H��� �����S�O�Y	��^�� ��e���^t��}�~91�TyL���P�B6�)���E�������=�4����J8X{@��11���v�)'��:TG=!Ab�o��|O�)J�xs3i�@1f�	�9>��/��n����\JS��gf�����U�[���#�)�����ꎴ^-����b���hhjf挊^�:������E9d#�Q�[�?R���t���t�rx�dz��5�%�m�|,���'�}��J����]�8��.�j�h���-`7"optҨjV��`O87� �R���0^�p��P��>���	�~��_�u�"{*�),�3�˽�
x�k_�o��o�).AϹ�e�`��hn��jE�θ8��!�����Z<���O��77+��Vv4#mZ�M�[���9��9��V��N�`yun�O+N��P?�Y!ǔXy�f`���pr&Ha��y�FlۺEAK&�5�����6%Ɓ��P����ϚJ�<Fߪ|V֔}�l�f6s��mH4'��?���j�܅bTe���?�w��/�T)KpA���~q֑�<��][��s�JP#�M�fS#�
$�	�#hd)��ux��U���{��Ҍ�����˲�4�"e˝���c�i��� ۸��X)�PQk��ް�W�r��U��6T�d�}���}�6�`�F�n� ���1 ��(˹ۻ�=�$��c3�������^4�DyL�%�����I�ڹS+w���
�����g�V���� �ݺO<�R�X��]\�'�|Be�/]���X��Hp��3D�S���׼��HhV�/s��������Gp��iY��Jyҕĩr��#;�ņ�L�0�CC���bQ�e�I����1y��̎`��S	��m��XCJ��f~W@{jZ-cP�v���S۳f�?�vCe�
�q�N&ۭ�\�zW�/��k�)��e`X#����z�̭O(�@c�%�9[��[�- gZ�@��ذi=��o��ｃ����>i�T�W.^®��o����d9z'�Æ4������ٸ|钼�<�P�`Ψ��"L`Z�4�D4��+W��_���_���g'$`�;� �}P���X����vo�EK2���O�v|�_�R��s�b��!�YgࠊGm̲;�]]zv��~,K���nQ�$��ewM���za�w���Q�%�K��u�3d���鬕���Um�G���B懥#h��y�	��n[�>�E�W���v��NY���111����'`Z�j�����a4R�R�`|avN���w�}��q6lX+粄u�6�,ؿ��Ø�IǕ��ԡ� 1F�bƵ�(Ʊb�gů�d�n�N��AwK��m`_��'��U�2��Y���6�8w��RIW��ױ5�IMI ��/�G� ����_E�L\��o
+��\��deX���gUҩ2n��*0��C��:_�^�0A��G��Mj�7 ]�_���Ŋ�;�5� ��s��"��G����ym �%# �lR:n�����nm}���')�T[����;���E�d=�D��4	�Ǡ�_��hįTS��]-��ַ�݇P�����TJ	���4�7>v
�>��`�&$:�8�N���p�z1�n����(&�����;Z�'e26s��I�c���sr�ݘ48��l���L�&�t�z/� ���n���ly�"�K_�����F����l�I�\�
k��,��ۨ_.��w������H <?;��ܝ�n.v�yY>�O�#�N�Ԗ�+viu��\ffg7*=�TaRAً��w��y��e9:Fl�e��mMq��b'SWp��u�=uRG�Ap��s��^�q�i��X1F�+������%\�Ʀ��h[�]�둯؂�}:�*��X����*�r��%ޜ`��p�dJ�SF�Jyl�ؽ����r%�onl�b�m���X*ȃ_`0X�M����W�E�FjՃ�:m�+ 8wx�yjFY]�&�	:�d�����::��-�2O�C�*6.���_��M��0��8\"]�	��c,�>߹3b��r�Y�a՜���7��wߕ8(�|.��g�bq1%�%&x�I�U8&A���
�_s Ҍ��ڂ�C���-�w�{�d��GA�?��n0��{%Jy�Ԏ�-z��{2��r5�S��%Kq��,e�I�pkE���)�u�*a_�����#C� ��\�F�Z�0��ưXͣ,��$�y)����-㲁�,��Fዒ,:��8w/��#$�G\.�`A��K_�R�h*U}�+tXǣ�ݭ�}��J�N����-7���N�[�z��R�9������A|�aX�#X���H�(f�t(5�@6�rm�՚.V�6m\���T�p̈qX�a�>�%	ܖ2Yu���X\*�A�"+U[�C�a�u���j�ና�Z`{o��]�4�%�IE7�r�qē�:ض���� )��7n����ز�>	:�kc�t��2��c�,�@�+��L>�q���A�k���ez����a�7���W��ăeh�Z������w�SUڢ7�BT���p_�2W9�Tg��~H�&G���zg;�q9S�K���޼e֭_���_��e	���c�kdl@h��9k[6mB��R>/��G�^�?���)�6y6nܼ�B&lj 7\g�P�Y�xp�:��a���Ӂ�=(� �[T�N��ʪ%���ѥ̢!��sr��?F�ڿó�~J��Ҍ�V�e)�|�X�#_��:|N�����%�7�w]�[��b������ca(֖g3,���������I�"y����x�\n\��x�U3�ɭ�}U:K�|}^d2٨=�O?���]¦u���3�(5�/��=\�k�q�^��e�� �4�Վm�Ui�����=��ҕ��@��eM3��>�h!�{�Y���p|���s��z���1-F��f�JvY�"a�Q$�.���E��г�vݏjq	'O������1�Yӧ��Ņ<Z�Cr�%���$����`VU���6�2���_��훡�3��V3U>��ܳS��s�p�U�\oo���Z��LeP� @�����h�>��[�Y�N�}ܔ,-)�{� G*�1 ۰a��tcV��)��}�E���B;�{�וH4*�����oV0�g�>��}�ܱ�۶��W��YGN�OP�,�s�9|>FSc#ҷ�p�L��7��@��������އ�hJ��}6ʯ�l?���~�Dg7�l���x��w��_��}{�=�V{�
s0\�*1��T�UZ&����cJG��-11(�/7v���lz�op���>�+UM�y_[i��zIHW���j���D,ae߫
��̾L���ʠ	N��V�Z�I��k���͛8�,����{��[�ی��b*r�>uΝ�4���KQ\%%�EMh//\�(`0�2���t�� FF�������h��z	Lx�y�V3���V�a��g�����شc��(�O ����r�~�cI�ʖ3��\�>���T�#�ѩ=����1�: �q�_����\:V{�w��nzU��ή�u����3��Zg"}쏵R��Yf�!�,x���]�|U)�T2�X[�Wᐵ`������,K`�9��l<�c���Z,�s�VLK�A�C��]�qM��5���hWgƖuvq@�cA��g�(&�Yc�5燒Bw��;ZK6%tT���8Ł���5( ��:�L���W�7��d������H�����Bl�SD*WQ����;��O^�>�"�m�(�/�Dv�#��Kb�"���f��ѦVM�h����z��A��D�z��?�Y������(Y�Ԙ��TἺ�3�d%�UY9����؎|��E��9��լ��H\��=.��21(̒u�Л��LqA��XIÄ�3�H�AeB�̻S}�+.�����MxO����
�Q���%	/]�-����(f%`�S�/���[�	�#�&k^ƥ�	�z�F�H��>7��媍y�z��5DZ���=�?sk[����sN������L�۱Zņe]�y�,Ț/�L�O1�{e�F���z�	L�bY��1�i�=xa�^]�ͪy�	V&����ς�Jw�tg���I���L���L+#������;�/q^4�D�q�K3�O�B^{�mM�1�?.��تY�
E9��KK�R�H|4;3�x�쵒��b&�r>#��$v�ǈ�U���6���K��||m��?~Hf���������tئg�VT-#0`�����eG���4 �Lmڼ��M�č�AlٺI4��A�5L��"M�',DC6���Ҹx��΢y�_�cO?�=7�:6W3��*_oI/�Υ�؉HT��<\
����$S������yU���[����l��Q8�1�'lao%�{*<��ظF�Ɲ�_R'�E#�N�I�A(�[�ڕVB%�"�\�sj��ݳ,�Q���X9llG�\�,�Ν;�#Q.9�O�H�#P(��3�N%�-3#��T���ǒ�ś�q��yt	�a�H\$R��FDZU�r�c���\����RWT�E%�`T���Ԙ��Ց�l�N(h�c�Y1��!͈��=F:W�U=;��a������s����������թ �D����*�"$/���0�zx�38�/g18p�8�(�e�s�1 �#(�K�eR��fA`̙t
U1,3�Ә�KZT����8���&̈́Q�Q�Rn9�4�
��ٱ�ǒ�Ա��t���U��FD��q1o�;� x�b�9~�=�P�]>��&���c�X�~�^8�S�`ݣ�������|Z�L�T�8�@�`�Y'���zvX��i�]U���3����,��l����+\v +@ԭ[h϶�Ca�Lk�~��~Z+�rx�V��1��j��V��P�4[�}�~V�~ T����4�K*x�d��T��ɖ�޹��E5���7mP092<���{O��ܱb.�X�z�qDH�&M���B&���5yC��%��x�~�����۸3�/�������\�PS���@��>dp�}�C<��Sx�SO���i�}bV<	�B�<�#<�W�S���N�4����i'}�ApL�7秪�+�4������`[z���
1yqo�^��L.�n5���݆}uZ�q��g�r�#N�V�I�������+r'��d�8���ѷz����+�=8<�6�ϣ��nL���H�ܵ�W���?�)��٭���%����~��3��a�Z�ԕDSG3b-qUg�H��3�����Fě�8k���ؼ�A��~�t�r�
��[5��ƚ[���q��,|�.L����K_�2>��~����[��
5*G�nV�|(ڠ~��&��ưu>����V�'s�^ Xs�����̿U-�f��ZW*"�JJ�6�,�,R�G �͙��DC(g:��رc8���R`%prr���9}�ܻ9�@�Z?% 7����3X
� \E�����$�IPX�z��&�k�6l���V�)�ψ�ȧ�s,���_�LlO!�L�`K��˖��[���I	��,���̊r)�
�q{�!ܽ?��!��f|��_��M��0`5D4�E1�%�;�X\�Ո�M�裰���ؿVQ��:�j��������xPW�ӧU&Su���:+Tk3Fī�;�JU��5�e�;P��N4��J��j��p{ � �^X�Ԃb�W^yUi�Ll�'M�Lb|t\|vYY.��0�H
l6�LQ�q�C�:8���K _�M�A��]2ٌ1	P�L�I`>�O~R�6�'&G���L�1�wN`"WFA�7E�s��<����]hj����ر�q�s��t{��)T�8^j�
�'�$h�(Az(ڄ`��&�9ϯd�,���M;���d��GN���{�z�����yv����T�o�Tq��{Z*q��:�%�t.�i�u���d�?��H�M�m)	`;� �Hl�b0A\ՙ�>]o�q)�@�e��@d�eKlez~�bSoݸ�"��PX�������
���)]|~goM<8�[p�S	�I�K�ރ�K�9���i,�l��w#D|)�bllk6�l�-��$�,{�>}E^�,���`�J��dȠ���Ok�:Z�_y�+&��D}M]o���)Ѹ�+��!D=!��d�'p����7�{����Tt�yUۺ�
;x��Ĵ��򙄏�a�3�GL4p&��-�^��BZG�D�w3��7	��� ֪%}~��Q���Z���ز ��w��*����"[F�l0�
�dp���/|����/UA�!Z1�l���H��*[��@���XiP���Y����QX����eU����?,���֬�����/����ߊA�)5�)T��F<֨����tb����9˘�`iG��Aߦ��K`N�(Щ�B�����iد�G�S��3.�ʃ�r���|W�+h����5�+�O�c����㕕���Y�Fp�Ҙs���52&;d���˱4�`����%��y�&.\����e1��s3�\=W�:(g^��t���[X�߯3bxPx�n�9�ͭ��^�KZU�74-����+12EҶ��"��e(���fv����?�[({���X#������rYK��u(�[qg�:&f��~t�J�붉�oǔ\�U�,:�8����>9�-;�)�`�%�ܬ�Dt��9o\��znU��	
�WU�n�v�~R�s5#�������1�����֞Ly<���kZ���*��l($B�JaRo����НAUD4���:>��9�����Rr�ٔ�Oq�3b@nݺ��y�$RH��� *q�L�r͞
��Z�0���\���Y�>�G\ǶM��#�j$��%o���AI$�����M,��އ7�;�;w��}�@��}c~���G�g�n��D���t�A3f��'��P$����,��������^���0`��'s`y+o��xm�7��`z�Z�}�$`��ܱ��GXqF�4��%0`�k*�(S��ԱҰ�0��iT-�S�8z����)�=g|��Oh&�*�˅.]��F�f`�ւ� �P�E�U�̒W	��� ߗ���W/#/�iN@��/����x����|�����8PO_?��p�:v�9��m�����5hhM��L�*gN@����-66o�%��"�]{T;���%��  ��g���g4$kE%:Vg,����T~������S���<4�����-�D���Y#P���w�}e���ʝEgf�j.�r^+aU���a0׮]U��'�_��6�sӺ�H�"�W�眛�S��~��G�'-�СC�|�2FGG�k׮]CsK��mnj��lZ�X��� ���ҴҔʥ����D3��**9Mmx����˟a}��2�O�����]m<Chl�Ƥܫ��,Z�v��4�W�:)�Ԅ={B� ��ñ0Y�e���� �g<��Sm�L��&��V�(��O0+���-�wD������z��V�/�cF�������[�U�kL|0�$21E5]Ce�� d2�f�J ���e�$,���B*��Q�'#�fI� ��*U͔[^���=mm�M�M�q�%$'0����RV�_	]�m���� ��t� ��uXZ\�Zۖ������Uex��C��]��r�S(4�ɝn�2�\b���ŝ/�\�W��H�.i�I�ںfƆ�?6�u��d�(��>��rM&&6i�5Y��b�Ԏ��Ú(deXiid�Pa�f�}����1�V`�3��Zy��@ys?=�^�s���y3
���cOY^�;�� ��bE��`A��p|l\�.�9�7[��g����f^���#�8��Nx��O>/�`���J󋨅�kl� ���R�M�c���m����G����א_��/"�֟Gm��\h�r�[�D�l$�=E*c��`y�7������2��ƛWk"3W4N(N*S͕l"ٷ��[�Vg7��#� �������f|��o*;jǂA7����ڰ�,fHl�#h]�W���Gr���=e%�8˭��<���}T��̒�{�-���bSj��k��&'�f��;\)�T$�w��˄?Ǥن��o�*+H�KYEeR�*b�S�=ϴ�:NF�Oǲ4�6��17��EUє�� {�#CF�-���A�A%Kz��3��b�z֬FDl)1�J._F��02�Ҽ�a�
���>eg��zYϊ�ֲ�ʎ�����d�e��hk�qS�v���z2�����lYQnb�~8рX��0l1h�
��f�[�hټ{%ӏ�֚D(.���6�4���ܬ��R��� դ�.��T	���F��-��ߓ�8��mzs�evy�8V�$.�*��vE�Ħ0i�^8`⚆PPFe��yͶW1%�[�;����B�:��ja)ߥ�z�uYp����k��{�j��{TE��#�,K�-�H� ��M,dp{|�Co=���vW1Ѻ<FH�G�@'нJgf�A���V�������GX ���a�58�BQU�9��}ałAiR����\�>h�k�*��֋�2�V]�+'{ʓ�.���]i&V�[3U�z%Q+M0�{Jat�\-�9��y�oHp��V/��l���e�ٰ����I�&Gv(�N.�)H��{��	���"0m��3�pgxD�9���K 09�����
�$M
HM���iB'����%��՟ӗn���9rI�G紷Ee�`�J(��V�Y�\�:�ڛ0/����/r.�MI�V���9U\�:6b�OX*�S?�+IۀJ<ن.㚠���v���C�]QD���4̎�ewj�����g{4f�|��G�՟��U��'����j���4�CI���iw�>M�x7�?u�8o&t)�#cȈ�eՐ�/�MokoSEɲO�j��&��A9;)�R�f�ձ�BU��$�+�����=�?� nM˺E�w��ɨ ��xk�Rj�]����9U�]�����!7`2%�=�3�^���N�Q���L��ǰT��*:a�j�"�Y9������+r��9L��IV{]r�Z�7V�vƒic>��t�ҀS���Z%��1�#���r�9F�ڕ+�-\.���̪��r��l|rm���߳b���D���_�~�e|�v0�����[7҈��1�@�8NR��h�
df&���@���Ke|������kw��V���l��6E#�\�\����)y�DC1LI����	{P�{�[-�=g�0v��VN�2�r��R���7�DA��9Us�����M�����1{a��f�^UR�i3���:����A��ޤ���I�Q���^��ʠ;���L��_��B�ɷ�fHY2����x�R"+������sf~�Zp��o�j��߯f�4�-�X�� �g�(Ljq	9y^;�@�n�^���}�$��d�D{��:�h{�����x��%�>wCWo�*�";5�tk+�z�(��'��	$`�|�Ȟ.-N��_�+oG��K~��'e�˶�҃�
���BL��O�<)-�a9�CS<�#�_&��H�#�ӱ޸�Xi����c0йc�V I_�ϳ�LJ��
U�z=(��:UT���4��'%��s��gy�I�,�M��3Fۆ/����L�ɖ M��'*]� �e	Ҧf�1�@����ZL�$4������w���+Dg��e9C*y_Y&��W�E϶�Ȱ�pvN�l�`�՚��H�NbV���#�;��"{Ŗ=}:�჏$�'�К�7I`�M[�3�b��2����o5�C� �sM�X��8/�*p���1YEj%����l_K�9�:̯�ܽe�����`�0%dhr��z�ިv�lD~(
� g�fpQ��ݫ�96e*������<�|�����Zƽ"ȥ�%PW=}톆?'lɷ�ω{*_�P�j�Y��k0=�<�dKrD񆜙N�����7��c���1�'g1��5	#�
�FTe'�<e��r�G�rꛢ��W\�`����yԦq��U]\�)�6}%uLAFQ6�;o<��c�� �mtJUӫ�{C�`�g*D��ؖ=�f�^��*�O���A\ؚlFgK�~W�0?3���	Mו���*,/��������j���<������s��0*�B?Ge[x�����CZ��r�Y2d���bI����3HJ ��։��nd�,RyT��� ��QP0*ذ��NliF�DE�1/n�gy^&|`�16|e�Ӝ/`�CZ�)�z�cb8oaE�#�w����t�Q�_()~�k���2O����'��1)I�U�̈��=H�󩠏V�e���߾�� f�F��q9�%	����Q���͸&b������T�g�X���%�3#��sR��Y��
И63����q���Y�@3���a
u�cMZwqR�/r�ER�zm���2�//��ǆ��r�0VM�����)�U��О�����|fV �3/�Rf����� ѹyy#���O�.�wV�-�PH�0k�!*�J��S����F�F��N#�&�҉�XOIoW��*M 6�&H�iul�+�#/��e�:�k��]�]��%�G�5��>{�]��%s��5D��K����޼�Jk��r.�Y��A��}�^f�\�Y^#BZ$i�� z�Ǧ���=�<�,y�\&��ׯabb\.�9��"�~�����s�� ��K�W�%�n��� ""#þ8�=>~IP��\��;�D5W@jfʜ.��Z��9�1N� +�#' ˞�#rXȏ�+�����9���^��YG�^YosB�I	����Ӹ�1����}�L��V���ʾhLi��>��Q3
���+x���`S�q�L��Q1Gڅ�U�1�,�pcG��2�l]�ƭg:d�&�)>1��$ �VZ�J�2��@4�C�;T����	'p��8�g�m�%�j�����
��Ov#&�e"U�O�� ������L�yxm���oA:���� {��������p��N֨і.8�)P*qP����1�p\�a�^s���ꩵ���j�px��� �[���0�(PN=��׼�$�U�h2?�7���âmm
�SоGlAUޯ�m�T��ՙ���E}����X���,Ts�����i�`U���-�.1��=J^���&�0A�]1� &3��V�Q1�Z�T2K�든�Wǒ@��X�b�[*�Ν	B^j�pKOM˞^B����2��,v��h�`g�`�-��kU5:���PG�z	H�_��Jf�b�k�M��7">�$ϑ��Z��^s��EIU%��k)��F�����~=�׫��Y��ɲ�q��R��Lv1�N`�l���؛Yv_e��޷�K�[ef�U�J�}�-�Hț^���f�1C��t�t�3�=����34����6�y�%[ri�}ɪ��}���s���{Ye]�������-�|��|��}�������OMLKC���VCb��m����GU�3��`<OF��[a\<c��sH��N\������d}�7�E_����8{�&RI�45�m��6���M׮�G��I=a��C��*C3u��w֤��`ua+2>{�(8�f�c�!���}ܖ9Χ?��t��ET�q�T@c�£XzS��L�
����sh����F�<:lk�$�z�Q�F��a��Ka@f�.��&�iP�6��J�=�9���Ү�HI����%c\Cц�u6o����&�  р7L��5J�b�� ��N�,�
��7��Y6?$�lF�P_R���瘼��YZX46�X}`��P�ڐB��u��)Ӝ��p4�i-K�\��[7�'�%�E_Y�ɭ6F��Ǥ�[�A39���o�ٿIut�hG���̻~	���W| ZC[wM����9��m��L/]��� T�P0준 H8�� ؗ FQ�6DP,Tt�}	lҒ�5}���ţ������{��� o�����-���I8/�b�$� &]���=���oH���5�tI�Z�fc���d2�l�:H�tm�	�w@�#:0�+32�6�S0]�@��겨ё�l�c�Bz��S�EqY�eec�4V�dC�O�ޑ�SJ
� �.��+n����0~)����!�V�t�lT.���
���5�j#a�t'��ca��/�I��<G5W�,!�b�P�����.W���2a i)��ghA�
TV�0�=5}@N��v��g�*�z��9�Ԇ��s��;��f�26"�܇�>��i�^��4ȴX�r{�Ԩ��#V6z7���C-0IIX��B�۪��Xە�gfENN�KZqdK�F��A�'1��څ�+Wy.�ѽ�P�%`�.L�G}a<�1�^�
J�!�cQɳ��w �Q�V#�A�_�T&jF��a�` �X�E}��LA�&��9����t��{�i��|�c�N`���(_�7���RiGV���F].�V0��wQI�m����;Q$�\�|��)���K�,E��H(���;�5H�'b�>��q���E{J���E�F��<7`42`��*���7��`���X�+Ǌ��*�?@;,����X�E_g� ������-a<�����5��lꁂ�dJ��*�#;���ʪ�S�+�ͤ҆b�\/1C�s���L���0��L*����vY!4Q�k��m����
Ā�1X�F� ��S�ل�
�����^B(����g����A!�T�c	a Pdȓf���\eV��!3V �8�0���:��<<�v��axb�Nf�����RQ��� c�PYc13���U�ҩ�4@"��nn����w��:�=)'Wy.�j@�_e`c�a�լ�ہ�Vw�'��hȠnX�_@�m�Zm�
��>��3F͎�4~�#��)Ra*
3陮0��Po���6�Fj�R"=0��Ȥ���FoO�`�oA33�HO�zZ��SP���̹>Ac<A���E+�g	�H�k��3���͝����$5@ ?<�)p ������{$H�p�QI'���Pc�D�k8E��Qy��F&���3�k�9k�])��Qp����� ]n�J�%sC�[���I7���Lu8�R���>@�{��B�	�{l�M�
��C1#�N
�iĠ�5����枺���_=S��b#�����;4�u( ,����t������w<V2 k��G3��!T�����L� 3i���1�]a5=lH�����Z�e�����
{0�#�;�w������'uٳR� ���.��%;�e��h�ʎ�Ͳd&�զe�	����yS�e]���%u8����!��$����ܘ�G���t)@b.�w����Fq�H�1ؓ.�7� i��q�
+E�4����G\ـ�
��?�NS�G��	P Q	�,��\	$�����E��
���lz�E�p��<���e����zS��]>[V���{
}^�F�
����p���Ȓ���=KU�ߠ*�,���LvH\�kmݷ������{�GezjZ��_�����!8��������=j"��htu�HB_c��1�;8�|w׷d}���K6�'�	�{�W]/�m7��h�/���F���a;�=�9��UB��i�j�6	1�Ce��v�K|�6��B���1ʺQi)�ľ�����@�.�0l8���R*X����{�~R��/ȥs�ٶ�`��	�H�ext��j�{m��c�/# 	,��� A��WcA{����E�
b\�@?��Φ<��ɓO>,��%y��y��{��Y�J�ڵE���ax��M�,����w��n��GqGgwG6`��~��=Ѐ(K�v�Fv��tY��'uk��6M଀ "'q��1��3�^��mGp������;���WT�=�G����F<j芘�d<���׉�z�'P� F14���#9)�=�Z�qU����J�+2^l�����4C�7��f�V5�7�17��C�UX�d� 7b)���DL`�E�^�g���-�ʡ�*�����"�Kץ��#ۑ�_))N'�4tm��w�t�Ӽ�;�����d9�����uO�cU(�1,� �=]`�\>����@��z3��k`�-D���#���
��p�o��U_i����f=�X�$�(	��(4-9q3�홤|���Q�Q_�Xa?!@r��9��lPx	ʒ��'	L"���62t���3�������*_iATO�,)G�7��8��v���.DjS���4 �U;Uq{�����mл���L�LȨ�}�D�m��^P���1�7�X�80OQ��:E�2��E\�^�e�/W�
�����h��O�p����(/z���=����U�v�6{؁��wI��bĴ�j��R��R��p,��k
$!�G��+�կ�w���~W���ƫ��ͅ�t;�(Dd�s҄��8;l�a;� �,���M�9)����*&C�o����	Ѧ2�0i���V'c�V��:S!4��ۥ�;�����i� ��n��\lYdУ�ր{ʷ�C"�7�����	�м�K[�M��
2q�(#y(u�u���_u6��D����!����T�}-���{�L�A��R'(,h!'���D��x���H�I��Һ��#�O[�G�Z�3s�6���j�.X�6�d��	|�|j�A�98A�>��Ft�`�#0���ü�|-�������ˬ�<OI\�.d�{zH�Je��=,O��Y�����:�����r���.���W��3�{Ek�ɚ$��R(�9P�ꥇ�A�����N �����c�,��G�ċ�R��P)��׎a�!@��ۯ:Vx·F�Z���Qwd0����&F�@����t:F-��%D�ĳB#��\[t���ɜ�}ƾ0Z����A'���2G4�淗D�e�N*�f�,�~0���4�H�CyT\���ݸTZpl1��s��<�ַ�۞�JbEzϼz^����2eXs��"ݤ���o��
#j75P�>@
&*'tߩ�eKrS����aҶ[�f������>����'�F7Ġ/
Yc�e_T�4��V�J����?�'�Og���̮X�}qLg��Q���BK����M�	��Lu�#�?l�G���ބ��N=&��%6Ǿ�7?転�zߜ7��!��C�,3t�Q�ß��^$1���q�AT8�	&[R���R�*{����H~X���H�C
�W�KfBf����6�N�R]���PCرYJ�2R�&���*�*��{���ޔ�+Cc����٩� ��R ���
	����g2��D�@��P�GҸ�諌`n�o�L �B�t�\���~������� �/��y�*u�k���V�����Հ
i�ݥ�h`��;��+�tM�
�GF��b�G`Ǥ
(l�$ԎE�]�;g�"�� �n�e��'�&�9�YMB�w�Tk������č1�ݲ�/,JS�����
Cd���NKg�+kחŇ���Җ�XC�kVmb���cs.�0�׮����gjW�*g%��dx�����]�1���5�;�ۡ*cvL�e��F{�i��0�	�V��;a�@o4���Og���ٯ�����L&��'F��?��g5 "� ��V[� &��n�
���ӝ���-�-�PU����Q��~s�37VV�9�x:8V*��Lm>3�Hxi�;��5���1Uu��g�@���0T��0����(�!�l��'4��HR���W������#e]��7��Mf%��6�/�����V�9j7����)���������G$@��U�A7�*P��6n|('M�8VM�lZ|�f@P�L�	������z 6U��Z����V[:%�(~j�X7T�q��307�8	��VI봀��k�Nh@iԵӠ�������7�@�p8l����rmT�T�Fe���%�����H�[�4����bv�(Tԧ���łY �0hb~��q2b��������z�ve����
��RY�MK�L��]�W��ڊ�4�]=�:��Pd�]��3�v�ow���\�z�46�$�� ���~�6-B�3)��a���F��7U�A�G�?�ar�"���7a;臤���d�� ������lF L���j����կ����� �f��%b�C�i
F���j/0�7�*����-q�c�b�e��ꡥu�6����K%M7�� �v2�t2�QG^P�|�a����&7Q9�+�����0��k{%V@�@b��5���yb���P}EN��oK<�笲+�Қ45������z_��v�@$|\��AB�ԶT�� ��5B{�v�+��xF};��0�!�4D8v+���}"C��|���X֣c�	���L�Q���3I�\?U;�L���9l��V�(����Xyw��6�rMkl/�G��xT�!|�u`�j�ӆ��_�2��1�:�����?���� �9V��ve0���H�{��A㡭�X3J�js$���ɖz%5zuf�[��lm�CT0���Qc���x���p�O��Q��KF�;�2{P/$�73�Ч��`�+��ș��cV��A��h��H���mE	��cE����
���md�תQ��gw(�ϔ=]|��*Hy����S\X� �AP��Ci!=:Uf\ǂ�x������\[�4ώ�22:&�dJ�;,�7`��d��e\A���h�]�\1#�>�0i}/��m�'<�K%6���o<��O)�JH^Fx�<�
�����6�h9��� j( Jz��P[]:�n�3}h����_���r�����a&DǙ�d�-������Dȧ��r�c�d��{v��B�`Sm��q�`%��뚟	�
4��xڻ��J ���s�����U������/�����o��2�޻��v������yy��Q�slALA�i��4�z�����\#duϲ��k�����ʦ�mT�W�ǈ��}@�Ň$8��籺�B���tǀYPeG�.�sg�}8d�{�B��Tq���?��;����1I����g�c��Cf|`r�!۳A����iѣC��F����t�������A	��p���Y�`�i�LVa@]�J�������j�-#3�x�PCV'Z/�����������O����$�q�z�חn���
�\<u|{�S���D�H?��͜�G�o]��Ά
��
�
���.��Y�>MPa��c�AWjL�~dL�h[�]�$�A첢 `ǋ���Ű�>D4"A[2���ii6���!F%Z-�$���03���%8��5YL� �Ձ�+��%��v�(���^�U�������n�ț��_T*SP;Q���.��W[_��l�WK��2㱿����
Z+���J�F2��H*0J�P2=85%1�Ug����:vR<�#�M��v��A�#U=!ݝ=O{�Aܐ��:!�°>��`�ӺQ��˳�uk�
����K��c`�7C�QU@�4"T�@�o��,7+��UV�q�P��(Ff��H���@)���L�́����/\Z��e���?yF@�9|��!Q��Њ?��J�"`�gb?�ջ�x���)Ѭ��(W�wYn�Sd��D�^!�#��SLĆHy<}��o?��$��L$lF���QI���� �枠@�H\�?��z��l)HlT+�u�o+�\Ss�z_s���⹃�AM���l�C�:��C��.��r(g���f�QY]Y�ju�}}��	*�5���E�/�d�b��'�{��'�ՎW8ˡ�Ȯ�7�TP���A�ׯJZM�X�VsL��'տ�c!�$P9�+c�V�~�5@E���'�ɰ�^ߌ>p��>n,�v�]`��1�vO���G��s�CF���ÜA@F
&b�2�J�{��=K�N�觊�vV�o�D?�H=3�6.DQ���a�N�h�[�%���.cz24=êf[� |1R�0O�1��n��w*�e���|&�5� ^�+���X��~��Ԫ5�r��,/-�b��ؿC�����/S|�2A�	L1�CCL6n��2���A.*P	Քsv^2�]�-�+��i8dk8`|�U�<{�&%(NrɆ��&��t+l#�-N�m}#ncZ2?"�f�%�1 �Q�v�ßA��J(�?����y��W)k���ݝM�齹yEd����N�B8e�)�o�-�87=wP��]OF��?׫Mί�E,�3��#�%#���5�P(��q��_��z�ʻR��Ln�X������g%��S���">LrϖT����H�FՖl��n�!񳸢���f�gL%$�b!̄�8~	g*�����dɠ*h�
|����.�"�:�T��Z%�ְ-6x��2��'YRu-�'�>�Z<�pl��`��kY����,���:z[y�����q��w�:<�����P�|kLĖ�;^��9�,��j+@�TT-�HW��*CT�,���Թǥ������O�'`���fբp F�:f$��хJ��sG�![���J���t��4K^C��g�&Յ,8"������;�k6���&�c4g\K;5�``e�����(�(���`�Њ����!����T�Ө�bC	@f�}ӗ p$�-��h��G Ř�Cp�ZK�z~G�4���� ����T֋�2��������������ݲ�-�������@�b�2�{�\խ-u�-i�m�i���+�OKF�Ȉǒ��s�$f5�)0�����2d`{S���ʬc�B������?��(��zf��`��i��A1��ǁ��)� �� �����)��Ml�>��b�L�@nP�#�?H��(�66��Э�����;~��f>'�Lm�,���W�)����T+`�g���k6����m+2���x�cՓ�ѽ���[���a��H5�����l���[�;��0�S�Cp�7��(@��VCU��~��^�~;��,;��  ��IDAT�c4� 3j�8gK��3PAs�}�%p�R�q���g�æG
6�gh�T|�fs� #f����2.��Ы�s
��l/.Z�w�hoUՀbx�"af�{
�h�z_$��;V�u�/��e�{�`x'Iw3�.�w���WՁ���韖T2��C����zܒ
���JP/K{sYv@M��R�@/��I$�὞T��&A�&�֪lC����!=� F��<H���34��V7���!�3��Hb�#�o� Y���{�Y�����d�y�c��Ւ����N�4�c	�V��$xwi�@��^�� 0�J+X-p�"+��P)��-T��5 @�j��x��_��U�vM�r CA��k�ry#��DFG�V@�T�����}��3ḹw�9XUB
J8|�8�V?T̏JJם���ۘ��R�ґ
�5)`�<pHF4@_�깭�bp�Z�!�DA�nR\��'"����/�n6��FcF`<���|\�	��tu�j�`p�Y�뺕�We��eE���25Y��?0��}a�d2�d����e)���BL�&DE�<���%JD�03@=�gS��IӟA�ب6�����0�U����w��+TD8gP��rd�F$�@�J��/�óGb	��.��!�@�I�0��!�Ğk�i���Du�;pϠ?	40h�%���$�@��%%1���C=�Z[���Uo[Z���/�ψ;� >+ٱ���)�3�,/I��k������\�(ټ��~���#?zd�%�A������Y0ۗ�$	��(��*l��136
"c�.^PH����<S�'������������_۰~tm��540�Ou]��˲~>�=���?���Y΍�P���Z��� �����nLRB��3�D��PA�ǻC��M&��@�O�Y_��A��5E�ڨ�5?��J�0�#� ʤc�A�u�'��D��L73sK����}ݧ��M��� *�ZzbF��]R�7�/�ݼ)^�=���G%��R�~#3T�5���ߒ!����9>�>t�(�����F(2�|���}ۛ[��zz֎d������;����F��;P>�����#�00� ^m��vI���oʍ�5z�+j��H�"��3�?���3l$��,E�b!ߪѣm�4\��ݖ��s���s�j�!F�l�64�9.�8ILK��=]�.ƍ �D��JM��X�#E/ɄJ�T�5$�5�+LLHjh�J�{���wRV����,�^�a=��h�$c�ڄ3��!������x&"�W/���4��fri]g���o��kkRS۽���ֵ�\{|�=��i���8 ���d��3>s���3������l�W����dڀ�W�h����O��n��Ij1���2�[�I&���i�ld�w�AQ�"J�o�:��4�����[������1ǘ�0��*/ѭ6}���=�cZs�g-���``���q�����Wo���/	��{��A9Ш�0�4�M5�[RVG�Pp��d$��Iq4��"���^�D��F��+�$�4b�ڻ�g�A�.i��?�n�P71�������6����4�X�� "@�@�56�%E(Ԉ���jpÙ,���L�8���(��{�)��j.K�a�
������X��}�h�frL\�[Yh�^vd��V�ݪ��֫5�����	�F��d�*�7n-I�Rg0�9�#Q8+(8&��&3��
K�Y�����Q�\կ�0-���
>����@Om곥ԉ�u}w0���O�Z���5H����
��gi�{%��l�#t8�	Z�t�躣��5Q���N
�/ל?8a4�ùU��c�S
R�� Ps�S#!@9�-�V���Lo��;�)l�ξ�f�ALƞ�e�[�p�R��o{m0h+Ѡ@� ^I���c��T�R���G��ӽ��{��p�E6t?��!��$��3=(�k���S!9��EA��Q6$Ȅ�h�v�oQ�b��afW=RP��ЗFU]z��`�Y��TX��0�٤4��� [J_7����n=`U	������U:?d�ٴ<qLW��t�	s�l >�p�ކ�����b�1wGl�'Ι ���S�$`5t�VMm�c:��q��ڍ4<���E~�u�5�{�1{��D�[�����\Nb�4�[S�-�����+�@,A��M��8V�k ��х�Nel>���:\d�k{��y�L������T2���(�_��@T�\�
X�Nn�(�#��.���dz,!��ޣAAD�YE�z�2��T��:�:3���
��jSl1|��_�)]=ǁ�!=G3w����9u�a��ޕ<���	$��d�"+z+��Ntt���,��˭^w�����F*2p�*�g�t�0�T=#٭�In��#��%l��%��I�Pbd��Ybv��@9�j4�|�,���VP�V{34\���u���ؐ�?�Q]Ø����6HvtX����xP����d���V ��OHHA��ʁ{����g�O�K��.Ҏ`��PJ?����Չ&A�X6*'�|X~����m��'c���I<H#�w
-����J�+����|��_�յ�ɔ����|D�U�?�B�\���`�-��8������q}C����rV�;u�d�p|V3��kT����e@i�M�����IʩI�`$�]����%��OK]�gy��>Ҁ�z!^���o՚14<N5�Zz��BA$b�>'ԟ�P�m@�ZO����*����l���zcA�jG�Iج��~F
3s�P;�Yz{�=�%�)XR�p��{eD�3�LsDK:�%���U$����N�#�?��~&�z��P��fF%=3d�U�Lx+@F�vg��l-_�ݽ��}?xP�zFB�Q�+�"��sa����~�!���q౩�9)�n������$��`V4�>��aH��1��(�����y眨�p V��`r�G؄�,���t���c-����OIs�+�Rc�P�ͤG)�C������T])�ں�)�	�z���]پy�酱���ōpYnrR�^�#�����.[��PP/�N�=v~@wU�P����sB�2Q����R�\�,�t^�g���Z�s=@n6Zr��-]Î����D�P�5(|I?۵�ߓ&z75���v��r�&�C��u����|J<&#̼�چ4�/�m��*�X����
UGQ�"�ƀ2��c���营!�?P�Jw�5�F0��
��8�����W R&���A[Q���f�T�H��/Z1���{:��oL�m�v�~F02����v!�g4�~#��ЭnnJK� ��mO�leY}QM�ِ�>`�U1��O���'w��|���@r�1V�V�.>���G
E�΍�u�5�1�3Z�����T7�������_�U��d��c'�s�n���e�80+�}��dGl�ܒ���l�uP3F�oץ��H:P}�=�������y�Vh�{�:ұŶ���;bp?�J���rϷz����z���X��8�Z�;pL�n'Xf���0A� D��b�?0�����_��i�\Sw?�	�9n?Xmtl5��N>v����:��F�B��Lj��-}�j�k�Ó�
$���edz^�Dd��14+����Ucғ,��\Ӡ25ٴ�cDCK7�� I�8>&��RR9_,H�R6r˘���G�ʝ�L����s��̙W�ЪJ\�c���#���G�Y�0ە��&u,@��pyn-ޒu=x��������!���}�h������5F������x �B�s:Pz�Lf!0CJ{� r4�����<7T���^�
�b���5
:����g�I%=� M�Ht�f[z
"<Dax���9	�K��6�z#�`C6���=.�BD���vt[0`���z���$����C�:գsc�M[��,CC��Nr��6�	`���n���E��g��})8h����'�����Ǻ�b��c���������I(��8����\��(F��\@Әz�G�/E�&=Vq9�vv�G�t���ܐ��b?0X��o��[ށZ��ء
5�V�R�p�9qQ����ּT��
���*K�\�h��rM=]���j1�[V`��J���ٕrhQ�/��YIf�$=�w�Ӡ\6�6��4���ޱ�y}���/&:��h�P=Ե827%?����`Õ���2T"��N ��A�z� �F��������8���n]�.��3����r����!�B<[�;\�����.G��R����?]�6�+I��; ���~�~�(�ElV��q����fV*U\�8d�]�G��7x�⩄���\��6��� �T�|P'�EX!�����D�y�+߫7�`��l�z�B�d�)@)N#jK�{l蕸y�ui5:2�`6������#E�rzǮ�1�-KW?�쉻i3k��Tt= �
�j�I'���_�����7�R+5\F�ץX���xXJ��ޓ6Y	�W�e�rb~N�zfo\_�����������1�굆�1u�5K#�9�ol�(�x�c���� ����~�t����*`h6z<���޿H**�� ��=V�l�LH��ra��h��")024����uh��|nP��\Q*gDa���(��@8O���B=4S�)7�(�~v�(�g6�e�/"}�S@���)�z�0�/_��"����k�ȺFv��_�lL �?|H��9J�.�h�*;RY��HƑ=��\Bʵ���IaVq�8}R��������g^|A.�=��:*�?��U[TLD�pU�NC����˄��6�@�T\Vv�e(�amuc�I�ś��}M��&g!��qOO��2>6)ׯ_ֵ�d��s������k�����'�ު�#B�
?���m����.a�n��$��H��
us�&�2�""��0$0�.��՗m��ҧ�^K����@�١�q����3I�8�2�:M�����Md��ǥv�:�)-ca��0�NO��H������I���{;�7KR����tJ2==+]�,��=��_�Y�D�*��������O1 :|h^��$](Ȩ�YT���0�P�VemeMn\�&�Ն���ڊ�,^�,��#SS��w��i��N\0:>N�o�K�M������S�s}��T�����~yV� l�n
��E�Pe�����bUs���=��]�B t��T�~!h�&*Bz@���GD�=IňAj��0�%��G��P$���%2d�/�Ð���z�"��8Ä{D����e��۲w�P����ҽLJ]}L���2h�Xc�[��>�V\"��2$�B������s�UU�?��?��Ǐ��{g�_��\�r����Q]�����'{����h=�ͪl��$����nE�{�%��ڒS��/�������_����$S��G�������P5�~��~bC`��j��s����@-�kA��o�p۠��d���ozQ�d�a�X�n��S�Ю�:i���Xz)��aS-D2I�x��;TǸU�QG�V-[�7[u�_G+e���Ƣ�*f�?vR�hR�jw��W��%�J��G��_��Ոm����Q��8����,�ξ)��S?/]�_���T���.�����Gw�Yc��SC_���QT�0�]�����7�X9r�${��@�$~϶[��h֫|�D�h����D˽���1:�G�7�GVӂ:*X;��@��5-k���}(���������޿���*�����LK�	����5C�;�ª��I&r5gC��M��������B�9��^�����w�\�&�|x9��p�4��r�	q��M@��6YV�Ô�<�HU8�͑�X@�7:1��&�Rė�N�AZY�h���
x��Q��
a�<T����\P2���S���U�Aiq��s�f���w�����$�ՊG$�`������]֋��&��ܫ�cbz�=(������f�X��	� JP�<>*_���w���)��c֚^���0�k@CE�*'���ʀ�F�w�V�<�B醬X�OE*����g�4�aR�}�Gh�̮�@���ذ�a�ר@�Z���%��H6����u��ށε�/�~&<�z	���GԱn닢	U�f�$�W��k����W0��葔��֧h���~�<��r��o+�ؑ��U�l:*ɃӬ���@"��,hj��x�kR�y@����
�����O�ۂ̸�N/��4y��:�=���(���k"=�o*Ddz�YCx��Ў)�{v(y�6�sf�^��	��ш[j@4�$��>�!C���i�V�u9Č'�fFja����Jn-
/fF�ޛ��$�[Jy
7�n�>K3�Ik�/j����7W�Q�� ݿ���VCn���,mZr��qy�Ԝ�����ҙWXy��#z��C�����1�=J/�rw`r���j>���'��\��
�C
���F�	�h��Y��"3�~����r��	�Ϋs��&�� ��#@��z~��ç8E26	T}���'ɉ!3/�r)]+H�S�
 W���~��D���T�e���PPˈy 3��N���D���KK���l�.����ɹ\�Y}TK����#;>����Q�S�(hhh���� ~&/C3�$���qRC{[+
V�R_�%��T���4`ƌ��}!F�'{[7�ÏKk�,�ǿ�yy酗��&�U�����.�k��Ȫ"x�U۷���w�̞�X:ɞ&��|��0၀��)��ꤑ��X���-��}�>��>�3��g�n�K_:FM�؇aP�� u�X�xB�p�th+!0�� K�H���{~K�QJ
�~�:�e��A!o<tF5�N�-�s\àӝ�Ȅ�FPs��u�q&�j5��t_!|��Q]��7��%����u��LCF���ؐ��v�4��*�ݻtYj�KR]ّ�ܸ݊yQ�(�%��}�q�j�N�T�T�_���,�^]>��?)o�q^~���%�������{���r����.;
�;j����1��l|dd����Xpl��;�����Wοy^��s����|.-����=���4˻�F���j��`:�"�s�wc�2TPr�,`�������(&��`L��J��I�V�?���`�6�3*̠s������4�Ay��P�Eu-�ER�����1����m��͍N��Y�niK��u)u�XN���!�J燧e�ߖ����XZ�}o���9��5�J�_GR�IJ�,^]����>y�٧�ܛo���eglD�?"'�:I!���k �ddtB?CA�G'	H��ښ���o����o��+I�}��g�?�Ϥ������_�����A�睃�Y.0ö}R��p8�"`吽�}+�2�^rL�/�H����I���}.��gp��2�k��l��o����#l04�,�{G�:�7c��R��>/Q鎁���eX�ى$�YQ��r��t�d�]�L4 ��U=i��5��/HE�YS�\gcI�O�d��`px{Ͻ���M�wu�9(�~�Y9{I}���L�7�N��O?%�N�%;{�L���`�Z�*T����I��b��V���ÏI�\a"�l܃8��TF�Z��/l����$GmU�F�Bwt�3w�7-.aV��� l�" ��@�v�IMw�]@!�o�]�q�>���<���Sj���g%5���x`*��A�̞DO��BN�7z�Kh_hz���d�������O����b�(׮ڦX�̃u5P�r��z�;�
	Bz/뻻���!�v�|���f��6"*�G������^zY��i
�C!����O�_�*�JIz�A��{��������(6��o� �+[S]���J�`��AD���m�`�z�1-b0�a:�ed�k��`yP�"u�W�5����&B=��?�En*�1h&��gƙ�mSh����&�eQ��Av2U����}�dc�7c�]�³��� ж.Ip�f?�۱㾊���z���%�����b6r�?�2׎c�Ǩ�E�+5
��m���67�0Za��LL|��i��+5��;�lI�fL�[�dh���0�ɩ���ڥ7�>��4���F����Ӊ��-R~y�єZ�bx؜���|�K_�����J��v��u{}�����=���;~�i�((0�������z��8�9��:4$�����)^�J��Lp��^��@P�A����Bp�3�Dv#��Ȍ�#w������k�كo�wl�9�U�/7:B�����F�ēR�B���pd�:���l�3Š���gG�EPeԡ.��_?���`j(/�������T�R���_�7�duu��	��?����n�n0�d�<�l�}��r��5^�Z�������8<,��sr���u��?(?��O1�k�cJz���� R&ճO�
�����'�g(��їh�A�`x9@W�8Dz�}�g��=���).5T<�N!̆��go���Q��N�����*�Paӡ`�>��.5<A�M�'=�=5F�҆�o^��~��aE�
J�z�E�[��+-�\�,1�A��Zz���;�-9ydL��������WC����&��΋/����>Ȟ	��Tm�$q O��>(f���_}^��2���1#��3��?�#R���W��	�y������0�|c�	�f�im���$*fB-��ƽ@c:����/&��3� ��b�ڤm�<�/�Y3;�� �~�HC�L~�o� �&)�p�z�!��Y#o:��۳<�����G������-~�~eG�t��]=�L���2�9(�b\4��ke}���ݺ,{�Nf�0P��jv%�7%���%��w��uS������_���Q���oJA���?(<p?�M�/��\&͑6�.R[�eQ.� <��M�ٖ�μ*�/��f�S�����'o�~N>���tɚDTm��e�_U��? o��]:��|�^C/)���;�kD@���]ӻ�c�\zYҖ�H`�:!`�j �3ZQ  \\o��C������� �������b�Asiz��[1H�YЄJ|5F�df�%�[����rMz{R�A�LӚ����KI'�Jg3+!oTmܮ��
��|�
|��V����P�vb�|�_���������k����B2shR�������#����Q�c��p6��@�I�5��7#g��]Ɍ���o{�|�'~\�8rH��ʗ�8�^[�+N�d_�
�qP����Y$��{a�=�5�8�/��q0���j7a�AGr,�>-_(̲�y��c/@�;����U���B5��j��۫��U�Ѣ��'z�E�a��1ԫ}�1�&��.Ґ��ǩ�I���d�]���/�W�IE����e���>˓�óRJ�L��t-J�m	$e5p��݇���ّ�UTP��Yړ͝]4岇�b��N�#�˷��~��ט�O�;�ykьn��A�*g����'�p�!����.���C���w��֖a6��<�ȣh�7b���B��!ǰ�p�=�
癊f BI6乬L������X���=�~b��}ި��9C�t;�5��@.�$�MF_*�t$DEU�"A;���b��g�s�H�Ov���K T_*��ީF,�;�x�쮬���{��R2<T���qI��&�_m���=����=C���qSX}��W.˛g/���MS�8��`d��ge����~�O��Q
A edxD�h�=f�FK8}�����d,�~�.�]�_����g���F���?�h������i�c��ى�ံ��a�p|X��YT7=�S�����A_��7H�XJ� �;��?8D���{�U��7bZ��bj�]�T���dme�^��b�O���]�Rۇ��gΞ�����y���tᐞ�y{k�U��U�;wx^��\_]���eV��@�(�F}���/���G�&�Ȑh4rp~J��(�:�={N��w/ʑ#'4H�rva\״�W���m��'O����!9q�.9{�~oOVַ�\kIq2��O]?��R
��z�s�`gfB�s{����CQ2.(��5��!���:FC�-7U=W͖���u������4M����y�qx�?�@�7b�Pt��j�:���wRC���q��gF�����/ܮ��F����������0��)��B�3�%
c�<fx ��z��[�zYZ��M2��S���T[����o��\:U������:3S���^����y�ɷ˨^�^��\[�!!���W����ܓ5�X5;�3S��\C�F	|�UP �]�����[����˙3�����ktd�=p����BөtM��{����Z3��L�(UD��:��fh,�娡b��`���4TC���C�a��߼�;����$�_C�������HETʯs��=N	u�#2#;�T���Fa�z,4����>���,��h��޼V��Ny��Ђ<V�<I�gO�%r��Q��-ݗS��}�C��ߒ7�����?&Z:�6U�x��F���3j��?�
[���W^%}ٝ��sr��A����m�quOv6�RW���~�� Fd�M��ϡ�����}1�?+do����Vɬ�c������X��oT9��ɶ*�����6��b6�t�`��+�L�����A�����n�J ��-��x���e=oz��� ^$6�z,E�	�40mU��Z�e�9@s.o2�Mڔ�����������j�W���,k ��=x��Oʁd]�n����2+kHZ���Ր�LL�ҽE_����-�����ϽO���Iy���^y��4�{R�gX��VJ��3����e�	�&z
A�wdD7_�b,��K�1HCb����a�z��Ee=�:�A����r��
���!F�:�a�&��f�+f ;b��]��-PG�(L��aG67�� ?е6V���䪓�D0?��F�����#}��9hi���dU�:�ߖ�Ԩ$!T��V�7�I&9���Y�0�8���=%�=���li >9�d�F\Cy�}ó6�:|�_����:�ᑢ�>}�><.�Y�CP��;d�qO@��X**���Bu����3��8��5;6TCT�1ө�A�}�lս��Rе*)�.�7�J+����~KjЧ�.5u�J�e�~����m*!�*Jd�Ʒq��3�>`��s
"�{�+)����wɭ�=Y��5��}in�)`)Ɍ��:�I]ɏKL���ٳ�X+�B�+P�3$]�Q����@�T��î�}���I�_�,�l���:kͲ�93c��K}涮%R�Ǻ�}���(s��|�A�$g`�w6��/?�Y)m������>u�;�{�I%�3q#�V`*�0�H�������D�m�{���
]?T�PD�6�k�_�Q3���P�	�8���}3ߗ�8�dq�F���D\& q;�%��kpK�$��JJ�ᡙ'd|(+����ە�g�N�]����܄ԑHJG��,��n=��f���Q9{�)gD��"j����F��稲����Y��a|	>��ڪ|���ʁ�2::.����L��, �K�Ҩ����'�N�׿�u&-߼pI~�3 #j��G�*h"Q���YL�?f�{���V�R�$"ꬎI��!�p@��m)FU'��B�΋��r����FB8<Ffļ��'XLv��-��U����Q�i� �Xj�RѢ����6Dp:��$By�[���?%ݽ*���=��׾!1�Ao}�cr���q92'O<��$1/T�d.Bі_���UP����U�R`{PH�hZ����my�;g���yx�Q&0rz�fL3aq���ޙW假����I�2)j @�p�ڢ��1	�������o�W��5y��g�]�}���� ���*�K 9����"}��"z�}*l�M}�t��T4}���Cӯa0��|��)�h��}P���`L�@����V������S8�?���L0�V"
2��\?z�<t|Dv��ؗ}��A���9}t^�p^^<sM���
iI�Ҋ
rhvN�8*+`���d�'	|��T6/Ӈ�JSmT���~�*�ӻ;�+JS��J�F�~��ݻy��σZ���.�p���[��W��|qXR���:F&Asx��d
�D�\�UFD� -Q�|a��Ƿ���B��Q��)&�q��6IX�>��,����B�.���;��V!��?}^�����@����'�G�����
�~@�Ə���',�s���16X��66�q� ��%�2����}�6�����Ɍ�qz��b�E?����j�a�a$d�����D������'�� �uܐ�.�������裏ʵ�ט=m5[R��J�1�(�󌎌��'�捛��׾&�~���������>����yK5�C��nWP=;Z·�An��|�oi71l��GN��i@Jr���Ī^ԽSZ�q�̱O�4��E����i�n����Z"�C��B���<�>/I<�`�oP\'��+�C�@/O�A#����.Z��!� �Qu�Ó�,u7�5��T@�J�j5�]u� ��w &��^33�2>2I~z"� ����'�c�q��t��.ɼ^�\�
��j�ٙU��2==-���W�Vnɲ�!�n���n���~+"����p07F$����Â̶:V���M (�T��%|{':3�V�k ���Y���*)�v��Q������C��H���DihB��~���!�珱c70�bYqu���P���粣	�%v���kj�і��MY�=�9zD���] C�uޞl.�5X���)����u}ww��;�6��v�T�-�r��e�ޛoRX!WնdJN?�
��~�˴ !)���"��`���)���}�iy��ȍ�%�������uy��7h�񺐊�A/��s6�{�g�ΎaP2Bfl��5�wC�u(Ba3Ԝ�f߷s�b���y���o3�}��-b)i�5���H��C�����X�/>�1��<8JH>	�}?���6����r��!�j?��R�~U�K����C225���S�Z����!��9vD���\�v�5i�dhnVʛ�V��^W?k8ˠ�3��r��u9p�g

9q�(龟���*�._�i}�ͭ-�u���A�Ҷ|���'�|R�����׿�<��w�=������R%�*2�xd�ɤ�-�ɣH��Jq��� 9a��uD��c��S(���(�u����b��ɴ�z�.�O:���$������GG��QЃ*:���<��ޒ3�z<7 �b!����P**�C���{���+XA��������D��'����|�=vL64�\U ���z������t�;����y��ߒf�i��%�����������_�<�\�=,�r�(��<�#|�ߔ?��?�����&�n���F�,O������P2��o|Kv5 <��+���_����1y�[�*_W��&	8K��F�v����v(�`o*@1��k�w6 �Gq��
ei �ga_!bF�x;6���~�k
H�p��ż�h`�y��{5δe*_P��`�sK!L�y{��"���Q���`�pe5���= ?���hF�Ð�e�"��?����-���?'�G��o��Pp��SRZY��A��������ӯꝪ�OQॢ���gk��!��ܐM��
4G�^��=61E� �3z�|�!))�8t�)�p�*��Hr�*G�m�+q���7�yV>�OJvZm�+A�8�g�rPp���?u0��������(�+����p#HքBd�t�h�,@�>���g�w@L�y@�g���Q"���C�Y�I_0/03���������C�#��4��۶>�e��@�yZ��������M�Q���<'kKKRH��}o�G�W�����2�����C�t�\[^�b;+���K�j���Ho74 Mf�8wP���T�-y��iI��ITG B������ �#Å!y�����{�Ӏr87J��f���g�B!A�I&�e{�q��uo���xn���LZ����k@�����~v��X �I}T��f@���uX^3�5
j��sKm����0��k�y���p��'�"a��z�T�ڙx�s�D5�b2�h�#��;<3Q����׿���8vT|�Y��,�#�'�r�M�k�K��e䮹Iy��]r�฼~iY�آ2�A�o�4���sdlLJ;!��y���ѡ�d����O����%0 0�y �E�V!��T��VF�ú���V�s��f8��F�-L`����0�֬��e^�~IdOT8.	M�����SB!;�6��l�A%���Y������������P<����-z���m������{��=���E���� ~�x0�A�*ę)���B���28��
�&o)�j�Fb�qicU������q��K;eY�|C�[r���;y�� =q��"�:�*�$5�W����˭�5n2:�3�2�Aü:d�+�.h��H����_p��CU)TD��]���8� �AK}�ȝ�pA^?� !��p�X'0s@���X9�(R��:��Q�B��[����%���8�D���i(!̄�0pK���fqq�1T)���8����۰O�L��A�ٮha�q��4��j��5�]'v�Q͚������{O(șae��A��K��k�3P�4�<v��T��p�,�.��n��q�b��\W��˯ȅK266-1}���hqD������E��� U�;�@�w�z��凞zJ�#�r��Q�'d�76�dwwKjj��m$�x<Aي�y�ł@�wSL��BE��p�f�tMQ92J�&ف�h��`�-��J�A���|Ѐ��Q�kRĄ�Ԩ|�j'��'�!f�}R}8gÍ0���,9 �%2R��Lǩ�J�ߒvU�NYN���ȣ˞��lF���>�Y9zp^~���Y,)0���_~A��:&� UX�ǋW����β�UC��=�  �a]_���%�N�}o}\F�2:>ƾ�Ri�����^���n�Ï<!�\Q2�{C#�K��qN�����ijp�P�h��ē�^`Ӕ�K3c����a�z�U�q�8/ĳ:(ǀ����޲�4]�J��wR1�o���&T+5f����qV݋��ޔ&�$39��1cg܁!�	��
�ۤ5�8�!]�	}�z<"{��Y��PV>�c�Oj��"
�������Kr�SO����ϑ��sv�7�?�{���?{䨄rChD��]�E���q�,-�ȁ�qu��)3�C��իW�����L�w/��h���w�q��L�Rf�|D���-���}����C��<��wɯ��a�sHh%C�l R�PQ��H�Xi��x�%����E���wI_��AJ����D2�<�H��=�u�R)������9�����ls�O�Z��كp����/5�R��t��&��ډ
��M�c���dD�����.92��^x]�><'���� ��S����O�y�{�O?��rUA��G��|�ú�����|6!���������z��$>M:� K�a��a�=11!���)l�AEMOPy{�=G?��E}]��U�(���4���W�B�z��J�<=9�Y���y�{ߧ�z^^:�:�AM���y M���-�zU=}�Ɗ>T��\d��x�z�� 7�NR�#*�s	��Y;I����Q�k5�ATipO���j�d�����|��D��v�e0����'����~!��*m��'�Fe�@Q��>���η?&����7�hxґS���s���?;;#Cs�孧�w?�C��#�'�NO2��~�R�/����}�Ob�!�4R��Pb\=�'-α��*���X�ư�/M~K��ʪ��z[��0����U�z��V8��V)ԕV�;���C&6�S�G���%�&i���6�B`=��ۗA���Ʈ�����.�����������0�z&��?h3PT-l�K쇲v׵C�C�_b�ѳ��C�g����P��g���ߜ*�ꜻ�eY�-[Ɩ�I�a��YX�s�Y`v8;�̞��3sfX�6`{����e˒�
�-uNU]9Wݪ����y���-�ð@٥�p�������y������?�y���a��_�%;��M�~%�����%����㶾�%ݸF�A�٩�&{�w #t�)�y"�+T���f�;�cx\���BV$VL,�$$�̖���X$�8��Z�N��p[vAcJ��3$�7��>A��Yd�J�t[�Ѐ�1\.K+4��i�i��!��(D@H�1A$�౗�¹f.�����gk=;Ib'��N[N�B<�!�#��ш��p��,�9���3��NH�l�Xf���2b��^%�dA�p�U{��ߌ�yծ�9e�{���7�k���!;]�oZ���}�K��u6}�aE�,y8�OB�v�Z�ykW��)�!-@<��w9Ĉd�����#F�b#�"������� @��]*��a��������5�W�{���7,{��X���,-O�G^�t-&�fS�XB��%ٵP��a��n� ���E历��N�p;1�γ:]?��ސ�����n����?^��q�ٍl2��*�?��Rt4ؐ�i:�ژ�t�2b�V���)��lY#_�Ӫۑ#������9d�EU{O������ڇ��N͔y8�di�=��}��������e��И��^���aLuu�8�	jS���X���Ӷ��j���@�200�M�B����E�$�߿�8`il�H*b�}�8������-o�ylH겐)���	�NG��i��wq���{�	g��aSU�n`��]N�s�#2�Ѡbq����AQe�Γ���ֶ�Dg�9�-s�������PM��P㎳!��b���چ$$H�����%B1K��>Ċ떒�F�dCC=����ÆFmzn��>;t`'ͬ������ٽw�����w������ЕS�h�WYe�cL Y��)�X\�M�c 03qm���	ǰ���������n��9w2isp�/#���C��R�H�,�a�#�y��g��MG����f7�Zn8Q��P"mɾ���H����ȠG6Q�� �C�R+����dM��j�k�аQC��<�d�s�%%�\@v2��
'�d0,N"R�-�)���0U��IF�P��shg�$q� �Zƶ� X�ݡ�h��Җ�a{��G�(������{��H*�����-TU�`������U[��m�:�䨦��^�h2ŕ�5��xB�v@�O�[O_������֖�Ck��,�menޚ���^�ec��+�"0%$���ŧljf����!R����;�C熱�t~�)�pK��o=u	�F�Yl�>�N=D\�f�ZN����3���6׫!�-?�����,�l�+����ZynP ����tlî�&�+�m7�N�"R*��R)]H6�Ǭ7�ħ�e륬:�oC�Vذ?���lw��F�����v;|� ��^����7�s��/~���,}��o[�U��R	{�g�z�+H��V��%��F�?7�D2�Q�ϕ�筈���]�Pg�u�OdF�l3���l���[n��{g�D�=�����@,a�ԙdwwY����2�Ŷ�h��T[N��Yd����G�VMD������R��%���()@h`HU.W�ϖ:����2���2��X�/��LT�"����6\���ʆ�vC�-��E�	�J��Y2��D��ů<j��7�f���N����x��|�}I|�;�ãv��U���}�μ���s�-�o�Ϳ�}�Gkˣ
���+��lp��F�U�asG�a��l��s�����۷w�f�{�It�������rƍA-;�L�����-9��[xF��c����m��7�#���Q���E+��2Y��e��|^�Q���BZ�3�p��$rFF��b��" L4�
�q��֔E�B6�����`�g��6�R�qP�^YM��d+��Lœb���v��E���c��~H]�<����G�iG�vYvv�F�b�~����>��m�?u^�a��u9A���9fO��V��$֋%%�į���$�v`|��Ӏ��c�"�#3v�X����v��KS��YE����7MX�Ù�m��4���9��b�SIɔ�!&6)�	�h&MV�u.�������!2��Yb"U"�Z3�1�[E��r,��p�$���!5�T����W8&ؒ
��YsX%q>�p�V����C�|�~�a݃�q����
�lk�`	*5�֭J���u���`,ӝ�������!q���#Ρ�P)��Q���U�J��L\-�6����;_G����PO4�#���-Ơc��$Ϛ[Z��+5�Y��w�W�����F���KR�4���Zjz�|��1	W���;������m��N|����m�2�5C�%?Q5��cb�e "s�;�t��ڶ��X����eE���{�ޏx}�e��6=3c�𩅭�����9��u�ؽӖ����I��u�ú��7�Μ<!��'��k2m��!ަ�X1���U%������b_���1����m�Di��Y��wr[Y1�����e��M<�|٦�g��9�����-�� [�,�@�Lⴈ���j��ؽ�q/�n��6�����5j�6��`���f�I޶���`M<���D;�����v�4����@H};7�^�)��������l�:�7T̄<'r��?:ɏ\,�5N,�M�B_�ܮM	��ހe8 ���Ĥ�փ��g�c�_z��}����7�ކ�v���'���!E�߰�=;T��bQV�:pw��kwYnc5`�Cf�9aպ�%[�ݹc�v���`0�L*����&��n&�ҳ���}�����?���?#)���`��M��C�0Lv��<����p���N��v|O�/���/D1<�b�u@�d��Y��ۮ�(����cGqsf��Q,`�����k+9�������ɢ֎�ME"_�6�KU'mׯeln������;j���}�~��z����9{���Y>�j>�A���<sʮL���5mǡ�H<�7,���b�B���ܖ	�ĺ�YU�DP��%�oxlT�����+�x�TR�D�@(��5��W���r�v��'���'O[�0W�.�!I���g OamQ~H��*�<7��i���Rj����3����@�@h�,��n���\#��។�`��d0�2Ț=�գ�:2��@F�φMCbcǂ+�>��lz��H���p��Bi�,�7'	�j����-۷g����-�����s��c�w���UU�ȃ���H*}8�!1�"V���g���`:��L�(�!xl��M��C%������F>s$�]6��h?���Ą]y����˿�){᥋�������U�Sw���o@�K�6K�E������3�`�*��p8�v��F�	x�D�XJ�����y%��}h���T�	]�:��.��� iK�E'��&LPZAw�:dN|>���Mx
�6�	���|�ME,��-R�bqCA:���ں�x�q؃M{�o��,�1-�aK���.�䉎�]���5����X���@����+c��|ov�Y6�)�>M!�=v�ȗ���m�G��X��d,$;U�}�C@�30��i�^={�%߇����'O��ۈ6d�8"CB�$E�s�c&���V,$�B�Bv�����#i�Hb��]!�BŴmU����"R��~�Ev`�,�J-�DK�0�8)h�U�	�U���K��.d˜�� ���l�6֫�B:`%$~�zeW����K��p_���^���B�������mme�.�>me2S�f|��B����.�AR�����s@�gd|���/�V�mzzZ�,f0�V K�$2\45 )�b�j�3s���0֐n	��n��	�龣h�'q~���H	�7�m�^���s����rs���,|Rsr]�Dh0�'�x�����D�4qF�G�t:;}M�����;���\�^�l���2�)���8�����F�*�z��a���mut9��u�����9f���G�-��c[H��ff����B��|u�V����1��ȧ���Sv�[�#G푧�#��Y�:so�_El�����m���x�/^�d��"���F�)��glff�)m��K���&cPN��z!�r���6�ssv���V,������>�uc���lvfɶVI��Z��јXD�?m��$�K�u�z��X�d
>��r�bfM6�-�ϰ�X� Y?�S|n�Sܣ���K��$��{e+�*T&D��/������-X�/��V"�B�)hwh��!J����j-;|l�~���
g!iK����r�6
9�d�`4p�ΟzѾܮ�������]�ۯ��/��^�N]<+�>\c
�"���[�����ۍJ�/�j�H[X�];�����T�������˶��ߨw���k�ktv�$V����M��F�Ο;���%[��$2�n<�v�d��y[�L4ֆ��p\s�<ӍbI���ѱa�*^8��]�\qs;g���>%�w'�.o�&aP�	���Q���h{iI0�+v��sNͱM�T�bH
�)����|�i�c�v�2�;콽��!�[�M��Ɉc�<q⬸ x�n:���^��flph�aDŀr1g���݅3gl���u���m�w�ޡ1�@سO	 .����'�/�h/�u�w��,�C~?O�~���t�2؋Ԇ�4*֏�!����F��հ����)ᴲn�W&�����������s���lm��#�t�ST�N.�]��P��!�a'���� ��ޙ��
�a����NDs���N��G ��ָ�v�/�i���^�)�XI��#�����aE+�9e�@�~�I{��I��=��-�S<dw��8▭n���ի�$ԅ�J�V�x߰��-�UE��H�fũO��I�A�pR��G:���u%�	^8gH{�g�F���<�?lݩn+��rk���� 3�sPs-<t0���f��3��б�]Ŏυf'H��&�ъ���Z�M'�J�?i����)B�_�bY�	n�X�q&��û��p��H���{Q'�@�V �N̵V��U�z`��U��j
AWֶ
�v��e�p�$ֳ���I�c��_w�}�c�Sg�ۉo���p��V�����{�D30,[�[����IF2��ca����[�_|��\VLTd	��9M>tᨓ��k�3@�T655GCB�Uy��Z��4���S�_ܬk�u&�a!z>�Cj6��"��L@:2nx����v��v ��� �(��_;7��~��S��F]G�]	vGZ~D�.�%ĥ�P�� �"&��kW�,$t��C�*o��N[�{p��HD5�۝q`8��'�λ�/}��!m�=8Jb�K Q���Ϡ5�p8o�J�OI�:��@���������z��s�3

�q��PȦf��s`��s����ܹ�
�GF�D�R��� 5�]j_r?��'��{�%���
k$��ٮ������2�H+�1n� 6�3��d�������}r��	�
�90&[!R"1��4�9�E��%�)}2 ��3�Bؼz�fꐬgb���aÐ.[�}w�e��)�Y�"iN�.$���v�w���s��l��G�g_��g���v��o[}+�ٜH�lC� ��)�U�1�m]����6��{DU�����㿏?��xzzJpa>�K�� HI$<I���V��6��SgϞ��Zrz�$�a��8?k��n�y��N��Ȟ
[J�4gx��G��[n�s/>�૥u����}E�W����;3�}fZ�cGo��YYZ����<p?���F �.#��Y3!k��6yuB�'E����5]�$K~����Cxc���(Ƥ�Aێ=D"&�L���L�~�g?j�{�=6֗��^>n�'.Z�8�������̢�m�n��m���)�E�0=;c;�x�q��Ep=3�.*I���o��<IDqAM������gY��_�~eRNhn�0l��������[�Bׄۏ�Y�:�M�����:�LƘ�r�����5���WD��t�Z�>�^���i�����w���~�榱T1+���
�C�FWG�$���u$��q����5�&��V���s����g��뿄g�Z�YuS4f�y�m|B�U���I�\��L�'B"��M����0��|�v�m�l�hܾ����<lY�zc�`Y\u��N}��q�j�foz��v�]G�$c3'NZ��d���aJ5l	 �Žo��6qa���I왼}�?���Hw��.�Y���LSL�J%v ��9f�kQ���cv�O��������p������-.X2�e�wkټ5�ܱ��[i;��	B��H�
��]�[�b�HX�i��j�u ;�QG8Q��S�$S(Q���5-tII��m�D؃�O0ۙ��?So/���1%�/9� )��5�n~����m8cV(#��(�MGƬ{�m�l����7����|��={�>�U�e���{�45i��E�c���cփק|Ki}�����sL�~�]:N��d'������˂���,0��}��:������/<+��^Q��?�I��s�/���V�Z�!�,�w��Mk���G�1��ǹ1�>�,&�\��{�a���Փ���Zq+���<%3σ�����ٞuwp���_w�c� y.=/H[�߂�2���:'�Zx���,>�8�_#�D#$�Y��^��ǵ_��n:����]{l.});|��޵��mbj�>`8�?M����Č�ccJ�(	�� ���_��ߝ�յU�8ǉ����f��K�$�bq��o����z4�{677g_���E���ܼd�v�ݏ8/��%�:����QR��uc��NzE-�Q�i��J�f�ٮ���x$�b��7ݸ��v����zh;��B�NO��C��&�k(���-�'=�{B4s��M�v�v��a�7��v�f׿��*�����?�Cl��$���X4ǐȌ��c�
�m"�a���J��Y�;o�ú�bw�r�������4��p���d|�{�_�[�rɆn��?dI�I)�f�q��=�2$��)I��a5"��"��Ԓ1V�I���!��&�yl�ՍU	�.M���Sg�̙s%S"�I���Gp�`����mU\�j;7��興���˦���}~��iUU4Ԅ`I��!)�%�9���v0�i���U��'�%�Ѥ#�i�]\��"�h��!���	��\8�d���m�p	U���>�㟴�w�K����W�~�l����+���G������7ljrRZ=��Hw�,_���?p�J��0�db_ ��YU�`�E�yj:��<?;��wD��aH�﷐�K�c�О��s���b׮^�!p0�U$�5魵DL �)!c��+L�k"TiY����\�5 ��~ �憆�4Do�U��nG���T�f7Z����s��m<ew�5��nu+�/%���;�S�hFCn.-���9_0��F(n��A� '��MG����3?m����~��翠��������x������8y�6�q�����޳C�9�9�9|�v��j_1�
y�ʚX8���e{�;O��A�ڝ��FM�=�A��9./.�b������ǟ�����	g@BJv��+����%�-u I�������5':vs�	i��Q��H��,���T\SB�� �-j/n��8��09dµ�Q�A��H��f�
��Qj�}"����� #䐰VUC-C!��I,k��"̔���G�V�zV`{��w��]��?����1{�ѿ��?k��?~C���ă���_��Y{�}��o�?�I3�	<�T�j_:n�_�w��kl��,���Ěe�Q�vZD��{|��d��ا�2M")���6Cn�"���@@�������B���}�M�a���k,����f,�lp"�Μ/��}{��.Xn}Q��"���A�9��.r�M]��5�K�kk*�MMM#٩��"�0j�eW��G�i�!��a7�A�<�H)$��HEx��gG�8��DP���fC0[��fWe=��E�Y���ѝ�%�^��W�p?>������}�[߰�4c�����������_lA:mQoڳޮ��b>������g�������øQ������\��Ͽ"X$׈�q�~�̈́*��� l�]�Y|�[�
;ж�~���:u!9����!��\[����hSD�$�������Nk�gddvnM]v����hd��髢^��E�Aҍu�U�Gٹvyݖ��r�{xh@���+da����#c�D����1�а{��A
���s>��4C�{����5��^����!�x���N����V��~���7�m��n�#�v�cv�-�u˯���7E^����
���V�°�Cݒ�h�Lb��b��#�ǟ���g�1�M��P��~��i�c�)\��Ȁ�E$F�o^�|�^x�%;��I�ي�~'��[æ���cq��Hb���ى��_���qZ�լ�}���\���}�G��t׮]6�sQ�ﲹ�i77��¾�ϡ=H$����&J;�$��+�l�?�X ��K�S�.�uE��"L����yiB���-_OF,8�4S��+��g�P�+'����G�\�}��ld��1<*��=ox�=��Q$�ث	�ɟ��}�}��3�a��+.�{���K��� 1�-JRy8O����l�ڔ`�])�g��uر�}t�s�G2��r���x^�}�1��y�:uI�{���ɿ��� 9A�������_BU�F��_���N������"RB�O2.�9;��aWO!��u�zcw�k�A#m�C���*��Ż`�����1M���H�^����l��7�NH���kS7�`9�jv�J8��sSv�ꔍ������!��8���ؽ��=��w����]����y{��Wle#k#Hs�u]/�vh��ݒ5[X^G �e��D���gյ���-#�$Y]�����Y����%[Z^��VN1���q�ֽ���]5N���W"�?��/�NU�v�Pܡ�?�ϧ"�z����qv�P��rf�6X�"���E#�ɾ`���K߿1�`��q�ɘ��|zII$`3`��������@��50R?�<^��vD��I�����voQ�Ā��\�k-Qj����	�������0������G>���6�����0�'�$rخm��~����f)��,6H��A��0��嬏�5�ܤ�A#D!��)'ǹ�-lȗ_~Yb�4�� b��Mȃ�����K9��P@@V��/��T��v#��X�e�R��a�|}:�J:���f������*��2!��e�C�+� ����^@j!�Q
���z�K���6������O�J&���ӯc�C{��-BJun.�-DB��bD/&�z$i��!A$�F���"�����þ��/"aX���a;��	���}�~�'?i���O�s�?fg�g-3<b#8t��-�h���|���d`��l"��ZϪo�_��/��pyeICU	�������hp8�}A�>�5���z�-: }�v������-����[m^S�"
,�-��or̅��䓌�A Ѥ3��~����Ź	��b��~����\g60gF����k��mñ;gH,��?����KVk#�Zy߂��a7��jRF$�겞ؘy�nSq/d��,m��/ۻ��!{�-o�/��W��G�J�h!8�-��8��DF���������ܣd���K��s�-��h����;E�#��vAu$��򭫧G{�ܙ�6}�ėc�v�ۛ��.^�d�=��:r6�೿y9C��?�.Ahn���X![��u�\��/��jI��f��ZK���Lr:?슱���sdd�~c{�E#
���OeHΏ�'2�>��8�\�Or4iN�S�3q�G�"m<��V����(4$zm����_��<��}��>b��t��Ш��cw���=�8��������W��do�F����mz�;D ���e��5��9{N��|R��-��v>�K��9g�����g��=���#vl��W�¹�v���-��"ù�V]P:7t��Ĩ,:ն�\�|��g��[>�� �����\'2����o�A�O�d�[6��u>;v�Y����;��Y�p�{u�[س�w��l]ec]V�,�^ JR�5�џL|@r�3�,}#�m"�ErXG ���^8�����S�}����v��;����͇���;o��seK�řk����>�l�_�����_[�ǟ��fi3��
�jx�9$��rQ�r�dW�N�����n���s�Go���
NKH(;{�DR�"����F@t��)$����gԙ���7�/���n��S��C�T��V@�AFE�W�&=�F�Zt�:;uG�A[�����Z0|��н�;SJb����c�S��Z������~����#�B�e"_��<!��Ӫ�`�~�C��m�����,r�T�kJ��*B�
��칋v��W�ɠ���C�l��C���Qk�bv��ؾ�lqv��p�S3�տ�+�|Ხ=��'�+¢ ��ID�&������-��Z�����}��O�u�_]����E�Q\�,���epdH3\��r�l���cW䩧�r:�x�l&��qv=ɬl+'�@�uF��+8lǒ|��./��-����I�۸3��N,:��b7���{{zTpP��E�=�cVW�a3:ǜ�e�!�̨H�gRR����i��r��siqQI�/x���\�D3�������GV��mf��������8�`Y�}���Wlsi�ʭ��p����65�lC���=��q#�i2�+��z�)��@"Ȃu,/_��gٸE�Dc�b����"��
��"��5"�p���>kW�iu։��*�k8�ߛ�-҈\��.4�%q�+�$�VER��U�h\K���1��i^����uvO�	�>��{�!�1��!�b����.�9��0�&#�
�9[%���u�(a�]�a�ކ� �����_�"fΎf/^�S�&-���ZkAz�l�4)(�鷳�����"�`��8���1�N��I�[B�PϘ7�A�7��M��a�ǭ��}��Y��;g�H�����ē)u������f�	!<x���������Iq�a�`7�sY��o]�c�kHd)G_C�	�u/+B���<6H�!�dA�(�L"%�ڨ�o����?�� ��PP�n��}tr��_������_��"�$ɠ`��������n}I��H�6�x��2^/��ޑ]6�^�������?���<8�{�{?f�r�Va(��.�X����Y�0@8���h,x`��9z�^m���Xq�����i��v�m�ة��C�d�c���㡡�Q/�)N�\���i	Y2��P���=|	�3�a#�@O�e�)���+p���J����'nsU}�z9%�rv
	�`���;]���Ga�X�sZun�EzZ����w�Z�*�z˖0�'����d�{���ٝ�#!�{�����Ε6�5�:m��k�����]8u�N<��u��sd��[�z�������M"���t�&��0ڵD��8t	�h�=64h��rL���+����$�n/��;�{�.U�}8�J�ębМm���,��������8�^�V;�o�� `%9!īiaV�+�[Ǚ��A`��!���Q��0Xgr_�m��NU�i	v�6a%t����5�kM9�4�L���ҷ��񰛵����H;-R ��%=�d'v���kS�=$
i��1�He(�Z���x��ӿ�m;�wك>h���졌=��#��?�c��c��x}�¬�r� �Q�m�.v�]�݆�e͖�fmmqI�lºn��f{�;ߡٟ����h,���3Y���s�������W�|y���{l�;�j��_����qЇ]
����w{a�����>�Ҍ}Lx������`n�zƙ.��*Ϥ���L�:��~'E;,�@�ŝ˲��'ґwW�~�g�P]s �pRL�C��0X�!J�.� �ڼ�C� 
PJn8cQiRޣlgNO�ī���>�E[���<	b��A�z�~�>��˷{ھ��w�+э �d�즊)����d��W/ؓO>����^�X�KbVcRO�Pv�ؕ�|t�1�2qgWw�|��)���T��H�L�����Hn�$Xe�09=A(�-f�
(���a-�n�^x^��N8�22Dr=*��a��x!7F=Q&|��Ŋ"�T�]%�	od�T�㬚��=6ua���sֲ���'��������9?G�w��;���1�1��7-��d��2�_Ö������ş6f7lc~f;��o�������E����]����q�]�0�b�կ�&��a1r�qN�s�e<��{��--ZAd��P�l�x��^�<�|I�&8S���wj}r��L�,��+V�孫�Ϧ&�����p%uԻ��a7(#C� �l�Qi8;m���SB�0ic�Z��a8��p�f(�-Z
4.i�]�	��FvU�!��c�Jb���%���\+��:eH6��
��x���F���C���ȿ��b��%k�	Y��r�{��ǣ*>\E�{�䫶�8���W��5�F�C�t�������[��*��
�)�[H������֪ �,�4��C�)1c�|��9u�77V,���w��c�=�k�kla+��j�B�Ik#��N7�ڼ�5B��NC����槦�~�wTt�bX.7zB���ʁd���Z.!�	9���T+H7���3.61ۆ�9�A�miH��3�"(#|�Ld���{l`�ߞ������D촼�����ΰ���l�l%������v��Θ������H��dP��-ui	g_mZ�d��F�ʴ-M�5��ؕ3�x�����p�._[@|���F��ԵMaߤ�3�Q���e�Y���N�3����b���M;y�e;{���+cVW��:8S*��\��4Vw�V��r�,����?�җ���s#k/��5�Db�����D�%;՝I�sw]�2v������QG�-z'1�;��������Pa70`w���0��s?�Ψ�.��V ی×�t�[A��yo���Y;�;�&3��M��H�20/U+ol)�CuZ��˗�WYkc��R	��|��$�l�i��$�S�8�S�Lo�>�fѝ�X��x4��;�g��ǒx�-��h�HG6ߨB�&�%.I	�g#%��n�`|�>$�V&�k<e�$��9�,�1���O��!i!���^��}��v�;�h -������:R�#y��+^g�＾��؞E���]�qq��$��D���7���v���h���Xx��pp�-�0��U懟~ў>��Uq`����خ�8�'m}�f���lmuE���=��eW6a�S8��ph5A pa|gg�q��k���C��A�����,ӕ٦?�-,,��f�P��YqHxtl�I@2L��8�^ �h��z��˶=4qզ�j����Il6+AL��1,��ii=�X�`G*,>�����N�񴠒 �2�H�Ǆ����!��9�D�E�VK9kб�ѴQd����yX=�C�2!�2%i�58�������ǟ��+ۡ}{~������7���v������S��ZP�V������SF`0;3#*�+�W���,Զo�IiUY]�\
�5I	n�nT�X~����"蚘�����y� A,��}��U���h���Y�sA��y�QP���������Y�lMs�a����ϙIi�f��Zwpz�&v茶�Q+q����A$<��5�h�*"8B:�.z��B0�d������f-®��@ԼTw:�%a�I��I��Bεl/����V7��U�G}D\��?�8�����IӪ�訆����g&��,a�y�q������l��	�|��rL���oa�Up���4�G~(#c#b"[^Z�� ����=������/�7&F���u��I���c?^�.���*�	r�(OC��3*�IGVB�]���-à�Tr<S��ęcb���,X6�3��D
�(�ZJ�+UӼ�RZ�O7�׬�e5�f�J[+��Hs��iy�%i�3!��{�?='0�@ezm����s�U�,����c�싧,�赕����l?ۓ8_Y$%�;F��:�g��������ڣH.�\��C�!8����d�d0$hYX\�E�9V�"�Y�to�;������+�9�Fp���o(xhhf"�� ����\a�$P�&���Px�b������H�,�x�=�|z%��$���%�i�S2,�`M9��V����p�X�g��ē�-ז������]@���6�c�`��ϟ�E��6�"i�8��*xF�W���K3v��',4Ы�ᵩ�6��)��Œ����(gl���¹�A2�f�3#��,]��P��"����]i]�W����ʫ�m+��M�9csW/��ڒfM	�
S���[���u��͊8�����+���֕����حb�p5H��B��H���d��x��7i�Y�⸅�{��{e�`$�	LBҰ������$S���v��y��2������#?V��V�EK�q���*��M�҄b!��,,lR;�Y�V"#R�8 "{V6�'i��KY���D���^���*p.��'!�N$�����G&ӭ}Hm��t	g۲�����!��� �YK�&&�K�?��ӏ&�qVBBH�q܏il��q}L����a�5i7^YXu�1��[�]ߒm�E���x�*�N�*$7Ȱ�<�_1he�JD-�C����4;AaX"��;�^`=���g{���X���M'�.���ZD1x�܆�)fq�&�B$�2$��Ym9�?��Al��,(��+� �]�\��#��#�0�f4�bQ������E"a8W�׬WJ�IV�ӓ����씊����ELao��:��eGbGmn~��VVu��fH�#��줭��چ�74���s�c��M�mׁ��'o�b?�(���G��=M	���PF�?��#$�ŗd�R,,;�숗k�3����Yg.�:y�#��p(���S	��Y]�0R$cAǳN�x�[��<S�H"���.!=�=Ju�O��{�ۧ� ��G|�D��8�K���b}2淂��H��B�^+�9u��{|�Ww��O�~�n��b`�HpV�y�N��h�K��|�lkW���#��̷�w9:���d?��݈S�����GG,34b�&�-Wh�?���x H�߮s�Y�����]B=;��E�d�6�g���1��O���u�`���۱d���I��y�u�����}Ё�^����݆�H�;�$��8K��5�(rM�(����d��'��k[���?/�Tj���cO�H�0����������u�̫6u��;����X�j��q ��/Y��i�p颭�o�p]�o!�-���)�2��\w�Ƌ��pb�*��aEֵ�Y��#a�D��>N�`��:��nЃ��ۣ�2�Z:UZ]��Ж��Q��S���$#������7��Q�Ϫ��:�҅c�I�#nelt��<���kg4���bח�p�k�V/��FS�O���j��E$��n��b�VC������k"")���矱���H~��o���A��0�9�Mb������oW/\�G�S"�k�[�:�E�k$�\Q�A[����8_Hh��L�#0��BV������K�)�`�C�ėS�Jb� Yy���Nt�do}C%��^fN��X��e����Cd ê.�MLL����l���vJ&]z����n���ҵ%R-%���n 8���ش剫b���u���Sե2sw�N4�T�/$t�j֖�\�f{���?���G�4�uBk�o#�����0�祚b�|��o��Սd�ǽ� �?w�X$��4�`Y�t�>A�Ir��]Je~�1L����=��Sv򥴃��,���mp��fg"n΢钂�Sq��.���-��y�l���'*��AB[g����IN�3Ex(ל$R���~�'�����7�I�WkxfI&�pZ�VUs<L�����˶.�VD�F�%�&�M|v+�� AڗL�񹸑��lH�Y�X6_�&y���V6�8�}�R��#K8�$o'��)�ЀMڲg���hȺ �֐���4�,��rY�I2��kE��m�i�67m�RQG�v�^�(i	��mvzZ�L��c��ZA�ι�U�/�=
�͂H*�@�,�^���sb���5���	K3*"%���m"y!QSY3}��y����%L Th�d���#	I:6��bBe�,m6��bt�I�Pw�F�w$t)%��6C΅&�s�/Ԑ�u�$l�Y�c�Oገhڴ���DPB�/{`sϏ"հ�$UaA-��XW��mn��}*�
�@P lT��0�͹�w�o$��M���څ�q���M����H_�P!�9������hq=�,�g��T3d��av���96cV��8�y��7�PkP3l$�O[��K��<�m��u�I\�P[؟�y%'���ɈJ�X��l_o�lE�^�n	���w�'d_��;�D�� @���s3ĥFG�s�/g5���p��	I���_�k�Z���T�b��FP%� ֨��v�����|��~��O��m�/qD":��|!/6���A�*r��M����������y��v�����`\aq
ϖ�8�%�*
_3	 "a|�;	��T�l�XS!rI4
Ļ�zV,p������#ܬQ(@n)l��p��P,�[uh���W���q{g=���y٬�hMv���ּ���gHs�,ʔ�qYbCø��Cp�(��U�k�8V���{&g��UGNd�12�J+A�f5��X�ə�9K�
�-��F�U��Gvڧ~�W��zӎ��^���i7�OK�2!n��|����o?.�B��;��q���!ux{�]������X$DK�.��Dau\Grp��D�`�櫈=�;I�ş	'Z*����v�Dۉ�_�� �f�T��Gw���S���.��`�5\"級}�wz|&z�>��e���NY�A��JY�1�xn�
g����P[�!�Q<�4�L���֋��J27ؒ(	}X����p�6�g8��K�u��-�ޏ��Y>bc����ɝ��\g����岥�������w����������݈�����uk<	I6���̂]�2c��KX�W`��	%^$��Ͳ���x��gp����D@i��~v�#'����y�J�׹$�W��h�x熟��v;	�v����?����N�z�{�a����[�vV)���W=GF��pv���y+�m�V84pb��DH������zGԍ{��Y8�.A:C;�;�'\�ǐ�`8O�g��,�wl�Rӳ��%P��!�x1^���!����;*è���.��`�LN^SE�ƃ�rR���r��e�yB���Y�3�rN�u]V���H�<ɹ8�4�i�Y��'u5��Y'I
���g�=!����!���#�G8��s�;z�]����0<����r�9ύ��4+ʖt�{e�*�CQ��v\��"5&Α�*�ZF �\&W��!.Yj���	%������E��}d�!B��f�V�X܋)#8ίl�*:������*S<��]�o	8��&9�=��"�*b�D���/�tY��#ˢ��*;�\�@���TM,�V�����?��o;X�����Y�Xj#�|dU�A2��	�%�g}�8R鸺���a �m ʤ�g`��� QM����>����|�P��5�)��>S���u|$�zB���he+d�x&]b}�Ưs�p�3̥�d;��NX�y4|�T�m2n��`/�>ulH��*5�M>/&����]���m0�k1H�B
�9W�`%1����/N�L`�yu���Sօ��Aa���g玢�J�8�=7ϥYd��@���C�:r�O%	�'�~���0�DY��*_W$)Au��ZGQg�?X���F"��J�l�8i��G9�I�v�_�Oq��F��/Σ��ݲVؑ.�G�`���3Fbǹj�j+��9�vLry�����	�Jd�o����L���[9]�k�-�!��|nC�0��9$��3���_xQ��kI'ׅ���׿^$\��d�[����2�Ab���d��-_�jñ�E<%��Kh�v�۵]q��Z���բ��Z�$n�m��րm����0![K������F@:55iݽ}R)C�Q��R䳎��'�C�E�=�7���]�"mV�׺R�� ���Na	k,IY"���3a�D]�&��4�Bvmʤ�3/���,h�z�"���F) ���"ƙ���vا~����yΕK�)�B�hSx���H�l�������,�ӣ����S��T0G����\��T7gzm}	�9j$X{�R��� g2�`T�Zdm8&�y(�IA.����m]�1����lҪk8�Z���c���� �UU��Pow�rH�:BU���C�=������u��*;�|�
|]�;mu$����H���e~���˕H<�
w-����o��M��b��d�ک��� ��H'bIǠ�)+�L�3H�%���bζ8"���G?�	������,P#%�1g�RqA���k��g^�W.NZ�okRY����Q{߻�b=��f��8��/�p_���:(�'8�k�E+#>�\ߴ��=���\A1�64�ٽj
�������(�V͖��x��yNo.@9m�Oc�p]�����n�s��1$*[[�8{���t��<bˍ�pv��)��9�
�<t��qf2b,�҇��
Y(@3q�U��6r�J�z-���⵶%�N*��T��XET`{�\-Qz˷�/�"���SW��V��
9�$A�߮���Ϋ�6*"N��zld�8w�=�7}����/��Ħ�<}&�&c�J	�yJ�$v�V6�o�^%*M����X�����,b:JAEq�E��bOu����R�sIq3P��N ��y�5_���I�5�6:�y��Ab�g��BQ[��a��ޮa�GBD'�Ӕ����6�읜M���sޙw8/�x���&�5[����뒐'�
q@�:�!q2$x�x�/� ��faWq�dmuI������鷏�~'��47�Րl��ܧX��3/_�j��\�𼋊�إ.
rSQ�>j{�X��E�*�r�Kv���;�n�Hقo�6q��F��mvk��W�5��$�c��t�m���]��v K�~7��o�P+��u�{5���Лf���S
��`��xɺrS$?,tl��,_U����*?�FX[۶��iwG�z�3PH'����jk������z`p��֭B��~$=�u�����E� j�7�	�2we��/�x�!8�,	�������0sf�c�4'R �|���ޣ%As�؆��07͎��$z{�E��Ci�ۓ�tA����l��{�l�{Cc�����x�A�Y���T(��E����֫R�fΕ�}�.��`~^ 5�+9�I��ÎF�B����H��� �LÝψ�]2蜅�_�s��h����r�]?����hΣH�	�z���I�C���zk�L���H�}��>fٵ5�9�Dyk���2���ڪc
�v��5{�ŗT)�I��hv���9�O{��#�45]e��CJ��$b�O�,a�my���4;JS砩��a��A%�%D�;7~��0��$�,�1��|K���0	��`��S݀���G��aG�,�
��8���D@� �C��<+u~B]Ԏs� V�9KZG�e�����Ż���k���A��nf_R�$��$~��M�cV@�R������?�.�4��`/)"��c�����I*���'푿y�V���P�}h�}���'�N҆G�k87;���E�o���IJ:գNC��F�ie��XF����=7N ���_�tlC���z�N��L>�Ң���JY���f� �v�b"N�5'J���ƽ�=��7<�S�u�� �&Y�)v�iK�O#��D���#�h6���#4*"���N���!�.U
�󄭋e��rt�L��._<��� �r	�ADb����ٿ���KIf�B2�y�nz�����(7��������}�ӿa��8a�1>Ϸ��m�k���H*��� 
�.�:�W6=��:�M[G ���ܬ�'��A,����tŌ��%���)"i�iSzm\b�eE�Ұ��`�٥={����?�ݧ�J����!K�$Yi����{C�-&�~0� 	 <ǖ�������7�l���+0��K���0�m� '���B�PP���Y��䍺:�e�'3qo�G�)����[�rkvmiÞ~��ۿ����w��Q�O(���
�Z���>��@µ&�+�5���LPC�6�(����xF,��S�0#��)�w��?����'l�ڌ�`���\�X3�f� 2c�9u$�`���MKfz�W�r�J�l�esDAς�n���s,\F���,�<?m��Q۷w�`��L��M\A�G���|I�k�	;>x�L���d�;6q�3�;l�ћp����$&�7�#@$Y/�>��=�8����T�뒫����9�B#!W�!�gˏ�5�[F�~��e˖�6=q�v��H��ba�EZDt,Tg�rH��`[�1����C���o��v��U[�ذ����9��@S���R�c�W���x��AE�9���{5c7��v��m'5����$�?����vPo���N;�mۆh��!cs0u�(|a�r;v�Xd��8g?Y���>�-.�5ځg�T��0�c��L'�Ls����}�ᛩ�v�[�r��ma��C�S�᫔`r�3����jY���V���@�u�_<�V@_�����Y;w����y�\���>$�,����$B�H�%��݌��J�7��v���]�2m�*mĕ�}�>�@�p4�]B@�o�lhl\�X��� y}�����V�s�>d�9�5ڿg��������Wg�~��P�c�v=Bq��\O>Ϯ�z�-��8���$��{��Hfs����� ��Ȏ6�b}2�G-�pRfJ9�Ɏ-� �x�,�1O�!͌8	%/�+�v�7�`�M�\<
�u�--�o��B�1��,�`#7-�����d��N<��H����xn��-BD�����G��ׇ��k��ǂ���i���
'2�uÂWj���B�iӅUp��F���ۭ���F�'�M��_S�z�ȑ��N��~]1��\ψ���m�Ll�QR�~��K�ty����~&jۿc�w��o���g�	��"BD�z��ӡ5uD'�"�O�nn_��������9��j��X*� �!����=�����X_̗���k�<�z���b;W��Uj!Q��l�n�n��� ��z5�J�uP+0 �등n1걒�ӗ�+W筈C���+��-�����>����M����)�� �s�0`�Lx��\Gغ�ǝ�7��dhÆ$d_��Yk�ʺ�ۺ��m�q^�/67s�sK���O��DЗr�z��wg �\@�F�8s�1d���E_[Y�5a�#pD	8TI�&@#��X�6i��3i��x�୓�$~�5��N�"��_�ᄯ�d=G��)/KOg���֚����a�A`ۨ�Ԑd��P�8ѐ�8gq�?~�.̯h���u"����^{��t��RAN���Y����T��[y[) l�,�3����XX��܃��H�)�@
o2���%%:����1�vB�.�K���!��e�	Ț�9F�jrv����~�-#�a1��Y�e
������aAM�@�%�0�uK�X�7i��[��q'].�������tq����y�#GS%�
ɹx�{�u���`}�<y}�q2i"�1��g�|��=z��#8�l,�$*���-�&�зb��@a��%���歆D�o�_0���;l筯�~���rgǑ[]穌{������/dS�˪�_8{�f�f]oWrʂ;?ZWZnZ�R*���Y.��6�L� 6�V��L.`�����+Im�D:i��r�� d�pllDLv���v��e�\D��,g�(ĂH�D�зs��i����[i��{���8;�jyFm`���,}K{Q,Vp�MU�9'G�=�
g;#!�3<�J����7e��Ť��/>-�)�z��)Y[Y���l/�za���W�w�_	6ej�a;z�{%*����h$��=���]&W|��:#��]��d3�i#�cꞝ�T��=�����[I�����jC�!��&��-d%&� %���&�a<��u���TPC�֕�(���v�R���`�p�~�$3,�1)2$�QC��3�&�_��[Ś-�1��ߒ��Z<ӏ3j���YK둌�趥�ҙb�,�b�9��
�}�"D;Pި��{F��D�
61w�~�w?�}�y�\�H����ڥ�%����^Ƴ�/�*Zb�0�Byt��v����,.گ���Y:�P��z~��RN��J����b��*��U����ꗨ9�[!u1��Ւ]x�6V׭g|Ć���.����s�G�0Ylሆ@�E��}��"�sQ���g��c�"�,*���'e��l��������cp�k.�O�ڰ7��=c��k�0�^J2L��,�!��`��������FIAX]���vG���v��5�M�@�5��8��lh��;��eA�/MN��˄%���WUH�J���\�mq���{��g�oP�g/k�2��519�ɘbva]�G��iqs='­��E�E�4�v8�Re�ϻ�t�O����#b ^����e%1q�?g1]!��%�831"�A`'�$MH63�q�K�+Qv��K�#	P(���{i$�R���C���B�FK.a���ND(`����`�]����L�2���I-Vƌ���|Q�5�Y$:���v�˹�ر�5u�����pޡ��(������^ב�����ar��V�q_���_�5�,�������G��l��q���0�j�Z�u�o,�1�o%왅�����֖����)��}&>�6H&ޝ��Yg��!#��ձ1��$�	����cƣB<�ݜ���i��1e¼�f����M�-s2�6=�ܝ
�$�!�r/�},�m�zX��M��|��h_��x-�LrD��~�,��!ّ�Ў�;m�{6�%��u��}�ӆ%���,\��^�D��⸐/I,��3.d��0G�Ͱ:�5�p�����c�FB,�_�߱g�H<w��e��3v��i1��8��A�:��t�ܳu�2퀌��mA����A�uC�V|���R'�
�|C��k�\��n񍉡�8��:�ҶkF���l���:�;�4�\ ��A�U������uJ���?�Z�.�6�C��ۖLP[�mkr��e7+de����E6��F���O�e#=��9����[q��0t�p�?�/f�xye�4d}㻤��Y�&6ͩs�t�R�}�Ua��t<�dC�s���]#�bi�B�$�����[5}�pT�vF�E�u}�:b�<�4�lHjS	U`�����4�ͤQ&$�Q��A��p��3�;,� �D�A.ٱ�ã��kE���6�L��X���[ZT�t~L�� ��\#M:�d��^��Cn�.$�ZS���0�04u0	�d���/����mh�/�78k$]]}"�i�3��.JH�9���lY�0w�¤-�Iz��(�ۥ�P��$;FL.�������L�*� �,�Xۄ����tΝp~����6lm��9D�s�.]�,�����<w5�TI%�
A:P�8̷딫bFx*H�M��sE��P!o]���>!�};w�{H��D�.�:���}���I9�$s����!�~0�Aթ���:�W��~���p�����X���bI#�U�S5�|�5�C�3^E0C2���Qk�{lǡA�źW���{����z��3��)��?��;���<{���\�J`/�!9,��H����kY���IN��7'����z�]'>�����Z+ۑFZ˲��h����Fr
9C;���p{��>���@J�}&.��+o}��)��I}̠!�,��Jw��T�Ia��iۀ�2�"G$E�<����+\�Ã���m�U���uzb�f�t}�?=�}L�6m�^�A���u��"�F���.7��P(��i�"	ΏV/Rg��݌�h��`�mC�c��{j�Bn�<�(H`�T�!�<�"�i؞���b�Q#�#���3?z��5`~Cg����S8S�Ġ��P���Q����#��ڡ�kn9/O<�g�`�, 4H�t����8}^�@ZR�� Hh��V�f�"l<X����ݻn���퐳�'��%=#u��jS����`zP�J�}�k�P�ur��g���0������2�.��70[b���f �b�|V)��kA@	Ht�,�	�����`F���w��������j[A,��̗�b�&u�m�3�� �-Qѯ�*���~�@"���A�� !��"9�tV�_ $��3R�I��i���l� ��L��g�A?�q�,�h���$�����h��n#4�#�6�}��,��d��k|B���,��q�6�}�ic���DAn���&�y��4m:$#��$RY/�΢���JJ�6��"K�HH��ʩ���m2�ߊ�P_*�T�<���ݴQD����@��l%�|�A��E�U���~�憈�\��.���>��G�P^[V�����h�ډ�&)��gct}M�r���`;��g�況b�������
f�S̊��i�k�N��:Dӝ$Պ������p�t]p�j)��9����dxh@��59��۲4}Uj���\1�cQ�~�^c�͎#�A�>$`�YB,�aL�N�=���QA&�j�]J$���t�r8��\�ĭWm�A��_�96�o� l�14�Th�)t�ܖ�& $�_�T�M�4Ħ${�)
I�@��d_����"�q��QЕ�"�B2�.ݮ:�XS��50��{F� ���i	��
����U=�9���0a�-��%���֪R]_���Y�3���B�#a\��q��j~�wxpp@����^%aa�TP{٢m
Z!������#��#���@���i]��%�b�a�5� ���S[][׳�X��|I�*�wq����4��l$,�c��`e�m-&�d�T��%胊���hiEj�EJ���K�=����2��I?�i\c�nY/Jc��q�u���b����g���(�鋔e\c�ݻ�yOJ�� S�ͦ�����kR�3��}�+�����~M�
��r¾��9iG�x������ivR6[Ơ̕��Ig��曅����I��|�1���I�vy�`��2���_�F�!1K��9~:=s��}�	6`���!D<�G�m���a;��A�Կ�c��6�_��K�X�ø�+��L�������¸nza�*o������[z ����//��k�8a�@"@��Q�6�Y?6�S��+�3rir�7��4�hF�'
O2*=�p�� ղ����>.	�|8L��k��A���/�5��T�y�� $!Ө#���k���`Wo66^#�as� 3�:2�㔊F�JwPG�  #-��tr�Y����@�\��AdA f��b��:붰�:��[�N�T���N]9/�'/���r��b.(��˹"̮ ���"�����kpW� �����S��� �	�$�d�ȓX3�QD�LJ���\ΰ�p�����V[Rz6@��J��5M{���a]�8G��9Q�h��6A�N���:�P��ݺ��+b T��}�(��
0��pI6�`����t�Q2P�H�n�
��c���d�M����ـ��M�����O���u��u�,�t�
K3���B���0�0lx��A,�����a�F9ŎT��rtV�Mz��/h��^�K�U�S���a�0	����>�B�[辴|�����@߀.g��OOs~>O C��5`I +�%�n����wA���:�4<����L#�%Tw='�3Uo���S�#	1�F�Α�J�l���(�(�mt���L���W��lj�R+�#��`7#�g3ؘ���I=� *�j03���D2%�j�@����U�Rʯp6E���5M�4���.yix��5*�s��$�R,�i��~ILR!C��t�&��|��Q
�!���{�B6�B�����km�Dp��r��i}6�b���n'�D�`�b���Ԇ쓰����Y(X8Ns��H���-�8X���G�ڥ�9��=��myqF֑�%V��	������7A�ds�M�a7d!A�="�$.�L"
잢��5��:����󑏶4)�ԯ�j��g�t@�P�(��ʪ\��(��iI�RF��S��n(bά��miL�e��D;:�lW�0#��6�YO�ED�_�#�S�If@Qtk�� N`�c�4M�&*�;��C�����Z7��X�e]&؀��8�!y�1ݣ�&P�t��.��;��@7�8����J��l�2��B{�(�i�U�4�9^��,��	��9�7Ȳ2 � .�Yh�Ci/��� �� J�-tĄ�Q�wHd��1@�DC�M�U���v�d�&�>g�פxX���k��4i]�N,� ZY-���}<y��A�̫�������O���F�k�.9��ܙT>#�/��g(Ip���r��%�� �h��EIg�є���!�tZ�L]��gN���$`g�HW)eA9�Z(��|�kk���S�؈��i ���a,f~�X�I/�=��H6��񘟺��{F�0Npa_@1_+�y�[�6#,H���K���{Ag.�&�f�ǌC���)9�c��v�&���m��تV�X��C��J~��4d>����{��c��+���X#���p���.ٿw��4fD	0R4"V��x�$�	0�Weii^���ɹsJD��qH00��Ɉ.���F�OZ)�Qr	rX,�q2�u��b,K�Z�WbI<;�u�o��a13M�M��ar_���ä#��=#��q�Fddg���1�zI ��/�.+bȶ�� �ۊ*�70��0�H�'H� ei��߈I&�ɮ����<��ʒ�ӳs��M�'$�ս��%���S��DE+��e]�]�����l����-�,��ރ�y�#�F��?�h���r�K}rJ��ٗ^����9ȣ���3�� M�h�B��4�E<��e{�[ZN��䬮���^E\�ٴ3N��VH�i���cW��2�\\��'�
��|���7@���_�۳���#j���D��6�ÌTl>��.���>6�P���aY1�a�f���s�za�TX3wA�=c@�t�-��s)q+�/K����^��rA2	�d)���oA���0㨾W@J���?�d��F2	t�m�qUy$�!�ٶ$�冼�fT�y�U�=�z�8 +�Bw"�n�;v(\Ҁ��κYF�$� �/f'
�^Љ�\�' X�5m����� �� v���9MT���Noh ^�.H,Yabf{�"0�c�q�����GIc�[�T���(|ӒBGw]bg3��fF����&ݑ��l�����5�� ��k�ZT&��7���j [!DA�0:,q�W�E.0z�F~�PG@K�U�G��gU_w��j��5��g?EM��&��'�ΆǊc�iC�莅����b7���)q ��:Ղ��:����z�3�jy3�^�}W,-�Ѣ��R�*�Q�= i�X�� �Dڇ��Eـ��Xg	o�uy�p�ۡf��������*^�d��4�[_!���2��<f�Ft���j��	�]�ZIb���B^���Xv�jdE=@�4T�e�T�X��/͑�6��@U���4KS�X�{�+Eޣ��x!��$HP�VjC�&OB��f8PV#A���"@d�n|�u���d�)�$,��	֚�� ���ȹ`Ď��VV֩�ԥ)��>?#�4 	4��Ū3��g�9�Hgq#-J˘�H�,��|cP�78M�nU�#�k��1� .��2����*�� �y��<ǀ�Q�������4� ��ݾ}�x��X�ouҖb��b̺��%C�S]�ٳges���-�Q$اV��H�p�.�L׮��M�A�-9闢��ɅN%��Gl�����@v����QXg�BM��c �]_�'���P�<�R)ʵ����ܒ1)R׋K�94	�9�ѳ��Q6���@��ċ:jƘH�G$��|vO��@�Z���&�)y������S&vl�@H���u��6�k�.�N� ���&�Wgf�W_�c/�,K��Nw��3����e�|!p�N"�T����aW֗W8o֤(�<œ_|�E�mK<��u� ���#k����ש����J�Ģ����t]
V�j/�܋�1����FΣ�Ϙ���2� ���`x���)�w��&u���Q��CwB����,����⬬��f����$�L*xp�l����{�H��!ϙpQq�����$K����5�Pz���Y���o�\:�fX�̊�٤��轪���KE�'Ю7�P���,��w�s/m�·9(7�����C]��y��U���SB���k�〇�ߑ'��]�uJJ�h;���!��ԳX���,�^ �U'yG�	�����@fڲ׵��~1�m7 `P��ͅ<�R�&�0�E$K�x�m��0���$���,n��٘/1���KmK��O`��V��X�ȉ�_�tս��,4���@B_%���\�����_��ܾ\.]��sgߗ}��;���2�����K@��o���դ�]xψ����hWN�4�ýo ��W.jY�.�5��H�&�m���CN����;���kƼQ�g]��
F�V}�W�Iֶ���e��g�a�a�U�l`/���՚C��LpۖҶ�����g��\2(z�[��60" wKE8X����Y�|c�i�s�DZ��d*�k�h�VEC�e�I����!�F��u��n��!/�/�����E	$��5�P:y�� �Vi��6�s��I9q���A�V�2���oc�����&�wp��~�]�.[��&S�f$���5��ޖ���ω��d<��4�:�|4tX��/L�!��yD;Ҳb�X|��7��'����~�Tb�~W��BH`���[#.p�+Ѵ��y�3��{�O������d�w�M�z�����;?B�����6�3q՞����S��,dx���A�J�C��Ā7oӀ��'�����C��\6�9�X0"PG�WbF�����r��9#2P
!��ٳk�58���b�T���ѣ�"���������L_fU�� ����w�^�0�c������!"���1E�89�Y��v����@����
�"���ա�\#̪��T\�c�ۛ�K7 �5=�K2�R$����b0QB<�.t���(Ń�LT���qH�l��<4L�+��(l�<$��Lf�Ξ�A ҋ����2�.A�I������'Oʹϲ���<���db|\p��	�BS]���5�/�l�5������笫�۪S 0�_:}n�#l���4IE����5]{Tu��7
��C���LI��@���j���Ɔu�,o�1�����d�gkK��[�xN�UJ�f��m[������y&ΦQ��R7�..$�*��G�0���S��n`('��I�Ɔeמ=2?�̎t���\��3��#�z� ^��g����+0I�ҙ�[�Gv��Av�95����4Ʈ�թ+2::B�����*��~��'dN�s,g�?B1倉�8V�z�G����ҵ�p�4'�U�M�$,����� ��Ơ���\$����� M��3k�aE%�kq3R4?��K�ܢҧ�ѩ�[�D�puΒ�k��a�3ps�X�����&R�@���H��I��n��=�S�<�����EٺmB�@>1y}�輕W���[:�&�5���M���w�=%��q���)=[YI:tX�������)M�2�uT�Z�l<C"nD�J��u�|����coH��M-�FB���c���8�䡳�$K���-ka�0%����M��"�k�9^r�<�g�H��=��X���f<+�V���9�����Hl r��N��ZP4$v���ܜlI3�4q̙�f0�uڙ\����X=�<#�6�:w�T�{�K*?p���ⷘ|�Ӟ/VeU�OWO�i�{��O��J����~~����7$�+�2���b�s�]j/����R+)�g��ٵ}�&�6��z>�"3ӗ��uh+�)�����~�-�C�!<���|��}��;�1#U�}C�
r1� �K��N:D��r�,�Kjߗ��M�K��_���A@�x�S����:ZvLZF ԙ<�`�*$;��%���A,ҹ�#�6�h�G����sy��*cVJ�������K�䏿&gΞ���	���i�&��镢����ޒ��k���*������k�l�;;6��&/^�{�7�>=�_����tuvZ�9��\���m���[�����΃ϊ�Py�7Y,��v`��@�Y̼a܂�r@p`�<��dA2"�@��*ao,�L���s�U�00Q7���
�(�Ap��>�y�X4�.�,EM�a��d@�b�$�K����;a�M�l�dD�M�@UC�S�:G������0��{�w�o�G���"k�U�����q|c�ѣ$��:#��%��j\�*�Z�_��,--sN]��&z9̈k��_��ӧ? A ��lN�m�.k�ZO<�v�n��=#�)Cjg!�N���A<=�� �o�=�u�s������P��b����В�L��I��}$� �B^k����w�$X�<��vɑ��D�a�4A��KFS���I$��Y T�;���t�i"�=8��&��FZ2d\V�LKW<+��GF�4lK�(9=',"$Ҵ���&y���}�2�"�|������l���}R4F����NFe�Ę�� �+�>ٺj6�I10��2)�-���9w颤4��λe�ޝ���r��	Mv}9t�-j�r��ݨ�
V8Fq�Ye3��g!(��I�;���K�S�GE]����A�CD���6��͆��zt�>mj�O���F���a��F�'� �4�$N���x�SxQ�'��#��Äaw��M&.�?(�I���W��S��[	���d����MÒR"j-���̱�k2Л�_��e(��HC/q�'t�@1�VD���1��CxZ���?�(�;�jm\����G_�a���ܡ�S,�5 ���P�E^���wޓ��|J
�+8�ʹ��B���AU��r�t}1�!_�9C�i�5�2S��.�`L�8HHVZ�xt������م �(�_hi41Qc�&�[?�k�����C���[����bTBg�u�%G�{|ϱ���e�pI�{& �4ȹ�����^&��`�|�zq�zqP����J�V�R�5�7���4Ь�Ŭh��S��������X�����[�9D�y��?��V�	u~����/���88G >���T� �i�Ld�0p*��H��4�\� ��K�j����k�k�p�9�3�j/��-���&;�0����4 i+�9��[�7$W���j�@QmT�i�휵�5�~�lE]�j�u�X�]��؄~���)��/�l�$#r����_���E��%G�{+��Ҭڷ��T� �:�i�WJt�g{s4�xo}#��s����(XQ�f�V��&�v��� �p7�`�� ���S���RG��j>:a(���^#�=Y�L*h��Fs]�q�>@��kӜ�MjR��:�ؿ�� ʘ�S#�� �B�� ��c�)~�Y��8	g�8S�rw��yM|Xvn���ݫ��`�]q]u�e��Fw���ň�\pvP�{T��Ή~����ܹ�r��;�f\Y�jhxD�Ol���)���C����U�kq�n޵M���B�/�M�=s�2mSg�KΜy�	��⼬��Y���."q���ȳ�I�@���
�,� 
�ʽ@�k��m�^W�B��®�����:��"�kV��1.��ެ�Z3a��c��Ө���P7@��G@�y9J1� ���$2���4$x�PZ��)��Z�W�eل�W`�Ѩ+{2�4�+I!�,�җź!)��E���oKM_�s`Tn>p�U������x^���8��!<7*=�=jWj������I��� ���M��dj�
���(�M�w���$��w?;`H4XB�I�7"Y\��x��	����m�xwR(z������sB�Y�1Tԗ�Ve�R�l�`�iꙊ��j�?��|	E�D���fg0j3� ӵ(�@�ҳ��J�j�KmDW��u���F����%�m�G� �ikRѬ�Ԇc'�'"L��|"� ~��ȸ�I���Y,���|��*
�w�}�\������?}Z��9�g�$�|U��̪�A�����ĉ���PL\޵]�&��8=3sm�������,�.�7��9��2�I�C��"��H�����MRF�	���qL"p������ �a�y�~n� � �:�zwo�=��Q��{2�!J�T�2~��QHO,Gr'��3�8M��m��b�?1]΀ɠi�!��YA�o6s�	 @�GHH!i�{�Ȁo�b������ڝ$m�g��e�����M��_��,�寮��|p�]Y�����>$��N1fK��j�n3�j72I蓮lJ�;�h?��#Vx��~�җ>'����w��s���5vƒ(���`>Q�2.�%5ڮȒHpf;�ԤWm H�ZxF:�x��4�ָ�B-���L@Er��S�F8��I�5#mCZ�ܠ�%�T�1��t9�?����D.#�ǻg((�r\U�P�<��Z�A$�>aG2&9HFE�a��Cҝ�A�V�(��:�@i�}O�͵�O70��4��]�T6�6�3�^:���Ç����S29y���=0��3�Ա���ݻvA���ʱc'dqnV���

(�$S)�;m6�K�hLT������s؅E��q�|7�ä�f�A��� ��J]w �H��^�ba	#�>�͔�:a#3$�1$����f[����L|#���a�%��b����5q���+x����z���N�:�U<G��u�TO6���0��?c3>����c��Č��V������~�,��ɷNȒX�l���������ɔ�����C 1IFY1�C�r���OK�9I�Ĺ�mv�@�RӤ	zz1=0��G۲u�PC��s?��ז�0�W$C���N`8��DNV8�_b�������  �h�c��CT���Lc� `���N�g`<��L��!iSǆ���4a46@=&=���_q�`~�b.�u�V�}/����d2"�#�X.]����TT���.==i��o��\�|�T�0l��%��$�dlpP�^����M
��_G�j@J�<������`hͤ$`\4�')A��N)`�����O~Bv�ي؁��������Om0�D����ŵǽ��S�Z� sm;WC:d�5:��O�Tʹ�<o�K[��@�%�H�q��琹V�LT\'F��M�Di<`�>b��v���܄063�Ɉ�M��KWI"��7[�
���~0���K��?���e��]o5��#G�,�>O�:�ե2Nux�9���>���:Ӣ��ʕˬ\�ؾ����<�=��/���'��Â��I�����'���N�F���x�ˉ�+��{�_�3�fdue���/�i0Ä���6�����ιܹ��H�[B��_�:@�:�t�&_uY�e���N���c��|��I�Ґpf��mP�hۊB8T�"��l���[&%���3�
��Ш�_ʳpr�����?�c�ߓG��L-,��7��!5��];wJZ��+/�L�Y$0'Ŭ��|^|�::��Z�&�3s��\WNn��,�/Ȼo�)1���/����n����sc$R.A�ŏhz��,� �5ؽ(�ܦ!�mAq6N'�Sny�C�L!�g'�!���Y���w����d�|�`W���OtC���@��纳G��ۤk`�޹nꡑ�"��5����ɏ8Dz1'D���:T��1�1�LũX�b]��d%���$��	�F((���忔v2-�z�r��I�͌wˎ�[�h����櫯�]�7���������#D
���NM_��.h�!���~E>����k�-�����������k�����F4�U����@�IB�b3 C(�
YLl�g���Ѻ���a0�b6[X\]'�TǤ�{���"�Fgݑ-�$ �1� qvB���������!(�v����-2<�C"\��V@�r$�Q�4A���1��r(	Σ�O���G��p���n"��i+?C�_��þ���m��.O?�}��4���4�������M��`���{�9<����� xQ�{�Y9qmR�7o��d��{�m$�9�������dqYme�F$љ�\zh����ɬ	�R1�b2��$��$c����#�� ��F}fZ�f̠�4�@�npr�w����30�&G<n�(�6l���Z7R"v�L�b;@��D���;w�m����_G���0�0:�4Ѩ����(�%�u��r�$���B�6��.�Z����&�H�����M$�	��If;�g5d��5�v.��ҋ1��4�����JwW��ɏ��8�&�t�^9z@~�1�K_�?uZ������eye��!�s�c8<��~ܺ��]M�
�G��^o���Ru����t҇V(.���P���W�U�1�-P�$�ƣql4\6b��x�/-��p�g(�4-�c���I6��g��@_�#�#��e�S�K,<�t�h�*�<	f2��l��x�K��QS�Q������ ֎��SO>)}�L�k<��es_N��o������������o�E��"	�<���8��'��/����ok\�Cy�(��iO�G�<eN�! M`���L��گ��=0+W�{�co����Vm�+۽���ˌ+�i�{���~	1���>]vdA���7�R�'�(e����u����J��Ї������c�#
@ó�G{k�����������z�����r����m�����ϺO��������Z����I���6� Q�Ѥ�R#�9��q����G(�t^/+�b ���g>-�fEN~pB����� P,JW�A7��/��O�����0tQ\yM��J���zX�dqeIΝ=K���~�g����h	�rI�u�@c�d0�.c�y�B8�H8C���ke8�%�aǌ 6lXA+p��z�D��,C��*D��\����0ą�p.W4��:���B49c���:��Gxy������j�
�\<ОO�W��K��b/�X�� �tve$��+S�y�O_�
����U����?x^�zI�h�q�wjB�,��_`0�
X.YgG�U�k׮���%�2q^�� {,p�w�~���W^�K/�z�G-�E"m2�	C��&�7+pH���>Z�u���0c�"�����e}^
�b?c֡e�P���ލ��������R#t(�h���d"���&�����S�dD�=�ـ�IT�ctVqe��n���Fw,m��hDK���Us~$A��4��V$��H�Y�W�<��VLv߼��믿.EM��5`ؾ}5�r]=2?3�F}��M���F�H�@}��CR�u���iY\��m�}�S����o���xK����;�{v���G>������<��֋9b�d,�4��#W�B7w.���8c)�-0S"�a2��<_�`WL�l�N�l�oq���������`��ֽ*���j�-5������n��Iq����7��i0`�I,ys�Q��f �@!	{Ȗ��� H�}��Օ9��JJ�G�Ԑ������//����7�&���$�9|��|B�$��
�P�4��2���R;�̌DX}}���Q�p��O~�����>}U��s_�yJq����uS��׀6��p��1�F��x���
| vU.��~a�0I��&�H�PYG� btr����5�V��0<�^���F	�]kB���@J��秉�HTj�LV��A�!�-���dpLb�^]���0��A!�vUuvg��"�!�����?c�H>��yŲ�4� v:שA@��ҥ���bF��n��'[�m�'��k��� t�#)o���ڶE��v����	)��g�b��{��d~a^�.-��j_�e�j�!=82(w�q�(�Q�L��z�"6�A���|#WBQ����Eu��u� ��]��ws���@y@g����5Y� {��}�23?G�4�:� �b��M���&gҙ��@�u�ƺ�}�Vt�4PNh�Mv����@d�Q����l�c���q�H"Ύ �����A�Ŏ3��*��X �]���3��!�� 0}�ɧ����K&���1����yGϴ�?J]������I�H�<x�=�[Z�q͢��)����k���������F�Ȉ��n^mEXj/�����	@3�8}��m	��Ȁ�� V���o����׽c�I�}?�����l�<��`0G����h�kE9=�~�H�N�t��&٢�O`t|Ml�d�|�Ԧ.F���{w��#c#�,$]��,W4Q������o� �y.]�~�o5�����/�c�S��l��t�����{�[&�I6����Av��x�M�ַ��$Њ���.s:�	�s�.٧��3��׎�oW�Ԑ��}���[�#h�� �U��m�"@�t�/C����j��H
I��əlH?��)LB�4��v"2���pZ�5t�}�@� .@�ngژ��� *���g�9j`]�6�ĺ���M�3m�T��'�&B`1OZ�w׶a�ik�t%�RP{���9]�����+[wL��Y��O��^����AI��XXZ�k3k���+��p��}�/C�wrRc�D4-[6�ʾ��e��K�A]�5~���2����÷�Ν{��`M��Iy��Y�]"�d�چMjw0�{x��HV��bD4-Ih�E�[_֯�_+�W��v"��+��mU��"
�6�`�|Cӊ�&�f�����P) bcJV:�V5��&���H����DE�q/����Ѻ���,`�腐���Q�/ך��6����0�	�O�y���͍߷��6Z��
�9X}��b�·��ziP���1aD��!�4`� Λe�����<�ا��$���<+���hp��Q�m��q`�:�r�� C�n���"��A�>1>&��7�;M{��-y�פ�ݤSER �>�Ś��Ȉc�t���u����p64�$!R��F2��'(i�$��q�y���O2	�`���r`���WI}�^�[�p�h���HJ��D���� �V�7�1���&�4غ&k��5]���G/`O �X�/%t�����4��HN]j�X���[��G�W^~Y�z�-0R�y�ڷ�b�צg�4H��>�� �Za��`||\�����ǿ�Y�{�K~�w�����5�@H�����z�%3ٛڎPƳ�D��u7�1�0.b=�I ӝ%1Y��Yq��[C�:�Qs���: �$(�4x|&t:{�ԟ�lV�4@Q��J������#,B@�\*��CP����+�h��'��Ŷ�E�6��q�AlƯ�fM>�� �VB�d.�+���x�X4��QY��}����,�+�����k�Jv�mG��#B��\aR�G@,1��fI��M����Ǚ,f4����~���?�J9�Ye���h`��TA:kQ�/��z��p�<���x�C�zn�4��%DA%u�F�S��1��(�� �aG����0KX�rg�]W$�� yd5QE�]E�B�S�O��l��ǸVQ�O%t�<#ab2Ȅ�c ���V��l��z��f논�:��56:Uc�Mh��fs4�=���6�LN&?|_������P*�)��i���ɐ&�c#���K�ȹ3g)n�_Ya�{����k�� ���C�+���23;'��>)�v2������$pN�'	Hh�ֻ��V��绩6�o�fz�J��$�uN$f����Y_[�4	�N��8umN���،�ޛ��a�$��C2���氰TV��C(>���Hhө����?K��2�祫o@�K5Y\+K;Ӗ�P�ET��RY$v�U� d�X��lӝI����K3�{M���Hd2zƶ�����gm]�#ۣ�M�C��A���a^�w~�w4��d�C�Ӫ4��Cwɷ��y��WȰ��������~�������: ��o��pN�>�����=)�hr����p��W�{P�7���["��H�e3eu��6�A���&:�I�$?`����Z$�)z�}�j����01ӋD��ZA��k�d1�� 2?�O�DY@X�['��n��r���o������Q�Ӥ.͂&��PE�1
��+Mhq�%���Λdߞ-���:� O=�L�_9|�v]�^��U��%}�l߶Yn��~�4�IuA�}�Gr��E�a|�����!��u���5�x�垶Ll��'�Ԧ������y��M�W�;梋kyB���n����o�{�_}EJ��?w��-��˜�N�����@�$�XR/3 Aˡ���uIu�=�9
�'�`Zͪ&�i>/�b( ��"J(5P>Q��ۑDÞ�ق��1~qs������	Y�(��,T��G���[��W8��Q��+"#Э�7�� �M�@F>��#2؛��ZCn;4$/���������_��$��'��1�ֽ{�#�b����Ӓ_\�n�E	} U*6<=aq8f�g5�ݻ�H�0�a���˼�<x?�?t_��+�Zx��F��i?��Z�j[+r��#r۽wʟ>�MY��Z�lxw�tl��|01gNVWO8�X�^i�Im�&*Q/� Ɂ��?F��r�1�l�e6VDB���n4�5�	H�O1�aI����p"�`+�wx)	&�m�0~|�i̻���`��;��At��ݻ$�Y��Ȏ�R+MK|}]ҝMS+��Ҝ��1�i�&M��evf��`h�F}k��ڇ�Mݲw�V�<�'�R��3��5H��{�e|l�%:u_Vt�._��x�Q��O}��k����3���,��W^����jG������'�^++�ړ�����_[�#�c�E�ߊϭ���@�eM�V�F<Z(����q��-�k��/���zV��61!�d�u,�����q߈��2�0s���'"�_�f��qv~H>�Ѣ�6��!q��A{�z#�1��Z��Gؾ���P ����4��Ө6���k k��xL�Y��v4*��~W#�	
�����S�:�Ab�F5�� �V�)5��h���Z�Kf�7,����ڹC�卵:y�y�ᣇ��G��#��Q6�uL,� R��Rdc��E\�M����([����!�ӭa(^I}��8<M���ox� �?�#�T�8�����`!��Q��Y0`�A��gL�����uC!�M�ƀ�^~-�։G��h�ȭӰ"���R�˙��
e$	ut���0W4PXԀ�^�I.��߻u|�lߺCN�R��sVguK�[__;�O}���Qy���� ���
!��*4W9;�N�Y�j0�Z��m$�Z��bU������qt�vkY)��������6:�g��a�u�\�,l0֘%�ݳOB�p�(vS#�Sw��y1gЈZ�x�{�a��3;��F�z�N��~<�Ԋ�ނ�`�*�L�7o�!��z�/]�U��&~:ETpY�v�@Oo�̽0-���y��5iD��K���ʮm;���>˄IE$j]�����41�4<,�=��N�{\f�f�;��s|��y��[�@����Q�t�\�]�>Hz����Hԭs��,m��-B\҄SWju�E���`u�uC�
i��4��e�x���Z�LxNh���n�����4��
���(`k5(T4�h�9B��G�7:���?��6є�����n���4�MbvM�N����RU�$��o�Y���̳;���2&�O'�9��ϝ!Dj��f=�uv�bjK5�z�W	E<����� a�1M� ƌ`�v���?�����w�M������3P߽o�ė���d��ώ9��.�2茡Q1�9�Ǡ��@ImU�Ƣ[��i��~��?�dj�&ɣP\AG��6�3�FFF�Ї���ɟcF�!�:���&]x6��t����u� ��o�#:A,��KAv�>O�]����;��Ytk���9�ֵ������rx��禼r��|�O�!�Ϝ�N]�@��X_���E�z̗@F�[�?tǲ��&Y%9q��<���c�.J3 *�w�MR�wPm+:�o;.33k�ӻ�{�.vd1�v��Y�>'���?#?|�G�ҳZG$�!ё1��4n"�,�3ѿ���l�Q�$Ý��-����Xh!��$ݗNZ��08ߠ�F}o����r#n�F�~Ey�X7FB���#i0�S� �\mRc3F�i����Ǒ�݇�,���.M,��tmZ�l�����|�{rp�f�����r^�.��=��j���@S�Weth���?.��Y�t��$�:X�CB��Cgȏ��"g����K�}h�����{L�G6���Y���}�����I!�ʀ�S����nr�N�]���-�g>�9��?���RB1Qm2�]݆�$Y��3 򾾾&)�AvZD����t�N6b�0<�q�6�t�QH�ȴ�=8^aE�ͽ-	CB�8���) ���7�A $D�w�KƷ���s�K5�p	xs��¥U������{�%y����G�{��+W�Jʯ�zH*ڢ61��ý=��5��رQ쭧����(�K�.�8����m;�ay����Mr�w1FJ��I����֖�7׭qJ�gkthDW��ڵ[ƷOH��g���g]�MS��t���5�� ���c�V�Aש�26l�����-���A?�)���a!!�fѵ�R�"����k6DC��3C}aH������_[01;��L��bHUk�xZ[Z��~^v��)��"�j�?<��x꓀|H�-׹>�F~��>4J��4�0�������+=��RۂYj	���zzrn�g�͘<�A[0ѤS�=D�z�' a�_��T������I�4��k^-W�Oז󔊋P;����_ ���2�ɴ���0ǎ��5m(c��̂�s�a�".9�f����������9��ϒ�7B�Aΐ@��ሖ("�B��8�r�`���P��KC��z��@���#a���	�<��]P%?���n?��9|[� ���7�iP��6���l�.,.�s?|���m��¡m�?%�	�5Y(��R2	��^:G��A�^/z�3+[�l��^{E^��	��{j��C��؄��i���l۲M6��*�������ś�l�$�J:l�Y�@g����Y w�\�	���@3�p	C�,`����4�%m}��7n�æ��~A.���I獊sӺ��c ���*|� 6��ލiz(/�Ǵ9��:0��u��r��v҉����	y����k��l��'ޑ�����q�&Mۊ���uWf礢7ǎ��
t��S���?���wj�7Fj�ѱ���4�>sZ.M^�G?�(h�q�:tN�ط���9������]�Y8�
0���u�uD�
�7/�&II��I�Zy�Nq=}:�o�bg�l�.d�i�f�Xp\�=��2�dDD���nQ���"84+��vt�0$q E~�M��� �Z��5p��Ba������_[��w�/��#2;�@�ą���g���&6���,�C�z��r��<�NmJ���t���H��+�33�ȦH@�RÝQgܫ	F�{��^�ot�Q%3���g倞�O�Q�4��ù0T��~�Y��͚l|����o����C^]�Y�dw��4��G��h\�ȋ�x��kZA�	��a�� �T�؇X�̝GZltI4�B�777�a,o��H.���p� �����:-2�ʺ_q�3� C�SR��⦤J�����Mp�z�"����yu�<���r˾~���I�}�����i ��&�Y!��G�ֳr�؛�!�[�e������oej梞�8���C����"����i�[� ��O��;���#G�UN�,��rUZ�t���Y�~O_?��[5��>��C�x�Y)��V0w�Amzӄtvw��
��(r�ا]�d

e�2E�Y
��2 $�DVRz?3�j�Q([6B��뚢��!�C|Z޷����Ђ!h��ާ��<K���I�Rz�M��c�潅$6���L�*SH
��QhB�/ޖ�[�H@�ǿ+����]����>9�{P����Y�����E>r�]��=#ٔ������ࡃz����~ s&CCÒՀr��K|� ��O�i�Nٱkg��G�YTLM�e��&C�}29}Q׾��)��3���'Mݟq\�����rU
��e�epkU�}��?;v@�@2"��Bh��d�O�ޠ�T�����R�p%3u�w�I�8t�0g�������#�l\6���-���>Ix�L���<�1D �*! �����Ä�������v��^�o���(~����/~V^}����w�S�!�⨮ao�<����E���G�s_����q&[(���W�	�)�i�]yhp@�Q�$/8S��s]j���F��Kܝ��!�"�N���h*��)��6�Mб"�H���I�F��C�ȉ�Z��<��V��U��-#�CIxO��t��B;���l(mP����19$
&J��j�D>|�)�p���4cOc1�6�Z�Ϫg#�z�������ܞ��R�̑� �B)p��"m����ʫ�?-�v���}{4~X��������ҟK�=Y�����޴��Pmt����;|;���S�q�6���-�>� ��Λ�W����������f���~oV��y�פ~�i"��C��&G��=k,dy:r9"^�-�F���w#4F�:�̲C
&��Z�=�,'��o��1�gGip��
6������k��Z�od:F��C�-i��w	�'��Ar	��T���A�1��%�L���V.��=9 ;�o����Ԭ�W��F�y&8#7}eN��%�v��C���˲�����I�Kh*�|��p����i�޹N�pL�%���&s�RR���K����ԤA�{9���
���j]�t�>��O�r~겼��+2�8�[��<�����>{$�6�h��s���l,,Kd8!9�`��M�m�z��F�R���nd���AY�:�r��X{#�`�f�|��B	!b3�hD���P.�%C[��@��Q\M\���]A^�Ghn�{�z	���Ʒ����߸�qn�?���E����0���Y6��V)B���5+/����"�5Ѹ|�IG�x�>)�F��tE>��Q9w���4c6������L�j��Ғ�tG�.g�Z��-�����G���`⒂�sqyE��i���z�,=z`ǆG�|ŵ���ڛ��'�G>�Y2�}��o�jYB�yQ�ތ�f�vSJ0*,K:5�xml�&w�HxPn���ê<���ǒ@#3�u�Y�LE��x��JU�T����y@H���Z�y�I��چ��8��e�?��m�K6ے�_9&[&���zP&?<-��e@�co�-�����zH/༼��ffӐ��A	U��������I5�R���ȭG��4&�F�߂�s��`k���ib!i���>T�أ�_������_>!�O��95��t�g�^�
�����Ei{��9�j)�0B�30H(8�r�í4�$��j���s:��Qw;Z~v�a�Š���!;���~-������T���'��"YA�B��0�p�������p�����+2�u�|��h�_�w�y[V����_�y=���AH͟������^/6ei~���uc��	G��j,����=��Cr�w�;�����y��Z2O
%T�ҧ��܂|x��$t/y���/|I�f�������t/���dt�.ҟc��Y_�;z�i��@�M�s��� �`�C�u:�0Ę�,N:l� IS�U
��FR��ة2���`���g4��d9�3b�"$e��(��1�5C����p�H���`C�:�k�10"g�>/����Eٽw���o�k9�o��|����}�ݯ��!I�:���h �i��H�1��N���7�ٹo��9��X�Qg��:�N\	��s]]^fu:��?��D6�e2������Y���Aؓ�QM��b��2FX,٠�Ea*Ya�zT!�6+�(��aN��8`�I
�F��)��e�=lh���7D~��K�ȳh�¦�5@�:!e� ��i��j��N}����0�唖�,��hjR�B@][j# M��4-���J6��-w���|�0�8 -�N����¨|b,��d��P|٤A���-$�A��A#�Ж�k���ӭ�.��h�Q�AG�Ɉ&��������-$�X�6��5��%�#���&���U�q�0�%��:��V���3J�o�z�>GV_AOE��*�ݬ�Gx?��N���9��Ś�ϥ�~ې4q3���I�:�~�U&���~_:����R��
��JK�~�/�DI�+�g���j�ѳ�/=]�Dx�U�� S~e����D�b�	��ރ��Զ�kr�{�n�Q��eس�٫�q@D�r./.���G������!�  E�>j�GGF)������*�$�7 7	�nz�7v(+�k�K/��a��+Ñ����HFra����$8���e� �Wjۼ;�|�Ԋ[7��|s���4
}ﺜ�:^Ш�mA��#�lZ�1��[��:B\�B|�V�ކN���́�s�=2ԗ�Ç���������~�@�G q���(�},�4�������6�)��z+�LSW��(�� ̨����2� ��hC��*��y���}�/-�ΉQ�
83�$�top_��9�N�|�!�E�W����iꚼ�L&|�K���3Be��f�i햓�i��ӯA�ɇ�c���=�=#y �M6���q��(�1,JѷQڵ�M�GȼJ}���Y��!�%���Qۑ�d��'&������d�T���i�'�9B�4F��o��[���}����iy��t=���ߣ1v��<cF8łc�HMANZ�[4f��z{�T�tJ�#'�u�ϩ�C�C}{�])�} �l\��ո� G4և��ӯ�(?x�G�E؞>}-����#�D&�B*¨����Pл����}O��nFS�P@Ʌ11�5|$�~���"FR�����5�8+�_�8}@7�"(ZbS�2���!g	�S�\��e�ߝ��l�g?�i�fJ!��s#y7 @���܍�0;"��h�'>�������a 1 ��7����7����/�ɯ��ߔ��sH�9�Dtc'Fz���5���a�3Kc�a�	b��:���a�Q��UN@9��.v�z�`C ��������nx���a����=?�Isr�w�K�7��YY-2p���EU� .(�Na> ���7�f��j(��� ha�An�n�}(6}}I���&>"�+���@5��Q�`�ߜa�1���Nc8車�F�〪�e�Qn�2�֫'������#��~��C��ɩ�����^���'?�+�";wn�Ύ.2���+�ȰJ��9��َ�t���h��m��a$5p*Ml0ԟ��f'�T����b��J�C������_�FF��_���k�9�O���2�F\^\f8�H:� m}@M�� ������!�S�I(*g����ʴ��@f��<V���M�q� S?���<a:�&3��hQ��G����@2�8�΍ �@%\�P�5����v���9�Z��mnjM^{�Y97|J��>ٵm���_~[���HU�}����s�N1����)�S�����{�,V���
Ht���Ȁ
:RYTC��ժ�u_�؁�&:e��&9 �<p�m�rU�Q��Q[���(�ȱ�n���hg)�.O4�c�Հ���Iԣ��W�.uv����w�j$�8#���ID����+j����J�A(Q҈�B����'��%���f2j� z�z����%��ۮ�َL���|A���w�R�ݠz�������#ٖ����u�rA���HOgu�}vi�|�4����a�苍�������&%٥	�����������H�&v�mѻ�tԒz7n9p���ꨏ�'#�Y��ӯ�.�A��;��3�nj�`��.��hю���3��=��BQ�{��p �B���Od��lP&Ε�@���}�]��38"`���:�?�|�?��B��cI��.q���Xw=佖&HxqV��ԖO�b_6������/���!B+������_�~���;�F��u��������yǣz��Ȁ(�������s3�-Ξ�j��B&uT�x�Q��S��o��#hߪ��/��/���q9}���2>8(�%De�X� �X\���)IA�c�D_h�D.�����K�N��,�u�u3hA����Z^:1ߋ�N��Z���"��"�"PG'����ݠ���͎���5���pƦ�BK�  �ʂRY&f$6ѽ �0��b�F}E$^���'��GdlS��?=+?��	�f�PLiP��Z҄����(#��늒Hk����hW0��]wݩ�N/G.]�"]�`�@Ąy��ꝇÂ�k�}+�%)T�evaVW�9�=�y�(@o?Ea��My���HN_���[�u�fdin���ym�S;N@9ESq����Y�4J�dӺ��Ms�&b���c(H3Os�9�<v����F��n��Q�ۋ�O�蠴�I���!�I�P�R*��O2���L�
K��k�lu��vH�`�tu&��瞓��U٭�3���E=w�N�SY)�|����[	]kpd&���q��q}�$���Ϟ�w�}OVWV�͉9uS�m�*g?<+�>�g���~cH����)�Xi��Sr��E������;�b~M�|�%Y�tY��Hݜ���ɫR�(�6#*z�t-Щ�iB��;�������(��"�K�{�v�t�MG����F�Zc��Zqوa����Q`M�AJ !�LC	2�d�~�S�L[7,L���irծ����sf�(s��,���0�L����C}��>��m��Ёa��F(��=0n�FB4�Py��eb˸�Ol�;}��ZQ��1��	Fя�~��o�=d"	$�>�ψ��ʓW�|[^��kԧ���m�
��g;�L�$6��4�Q����I�*��<�qT����v�Q��L�y��+2=yY��ɑQ���b���aT���>I0��^D��_�U��캷L�t�m�$�F� �Pt9�Z�����[g7(7F� �����:����\"�F����7T��'	`�?~�k7&�χG퍍��'��>!�=�S@2�A��j��{��j�;3z���r���l��\*�*	
@˶Q�I= �������HYz�0��9����A�0lh���_�8��Ny|ˈ��I
��W/��X�t&��k����u����	�`��AB|q,f��uC��Ƽ�u�����>��を��D�uP������:v��UýF�D�=�\狉����C�^כ�����@4�ئ��'dlxHF5؄ 54��~x���#�C�ʩ.�Y5jZ����O��ň�̭���M]�$�G�D�όي��9&���ftϩ}���AU�B��پE��t���ZI����L^��rVR`�D���ɞ	�� ��ʎg��W�W�M��c��ʎiDv�6&)t��NL��?"�ݨh�묳�d���\�	���/X?�k�?��#$�5�����:�Qa#�OV��o@܀�� �V#Y.�rih˨��/�2g7�M�A[�5L�Sr���s_��&-�2}�P$� (�W6���7��y��m|_+��vB԰ALz�	v�/L^�nu�H�Qh���E9
V�jҋy�G��ڬA9���L�,���|F�#�M}�h2�Af~a���b���v��,�ڃ����~W�UJYxф�7���bš�Q����wc:S;�*#�5i@��ګ�(�p$I2`~�sՌ��0��q��ltN�>�k�)T�#np{Јꮾ��̜��g���v˿�(C}����ՙv��w�ĺ,{o�-��;���Q�ɫ�  ��IDAT"�r��߹[&&�x��}�=Mf���+�,Ȳ�O<��<������"1u2#z��4����{����<�i�R�����CN������g�e�y���s��y�gzrB�HD"(
�dK+q�������֖]��lYv�ZU��k˪�XiٔH�@�L��3����s<�>�wnπ�\*�1���{������<?����jvS�(�֚֋��\Ѥa���A`zMs�]�a�l����q̕�.�Y���P���G�MM�~7�"ס׳��k���/f��%�z����AU���\�G�C���P.�j4mq�7�����M�E!t (̨-�;����'�)S;�O�1����䍟�)�����������k9|�Q�G� @��?����W�0:q�7��#(?p`��5C�s����ޜ���>BB�Z����wޕw�{_��W��?d��^�c�ܨ�y��Ѹ��]$�y������?�$�*�瞗���^�(�ץ��c
�ͤ��R�[���ŇY%}^d��5Q	���2�RR�!p�x���{b�&��$�¬�&�*��~E�%c��!���1��ڒ�b
2 f��M��)���Ttn���8A6Y��D(��H�;�^� �%�Qc�H�0s�)D�##��21�O������B��e.vT�R�رS�M_�?<��S�M`?b�`�3�˫$$����`Zx�Qٱ{JV5���ؐ�g��t��w���<�wѢ|�S#d��HI�����g�v�xX��{1FP�J�:x@�k�$U��ss7eeu�~��5ڿ�f���!&�>v�q":�팪X􉘵u;A��������+�#� �E㵵��m�p��5@���Y�HZ�/��§g����O=(���òk�!j����+s�U	DS2��`l�+�;���KKz�#~���N&4���{�gϒ�x���&����.y��g�S���F�g^�~{=W*�ǟ��k37���+2�cR^��,�&:�S�E� _�8�o�s�d.��\��j�#;�fP��]2��	���̪��P��1:�]M��AB��N�Vg16>�	Hː�b^c����E|b�����3d�@Dz��R��L�=�6�na�?�Ͼ1��{l��|;V�$�w4*�tJ2�&���tZ�[y$���Q���	��h�7/[�c7��+M2WONMh���p�:�*����*���(湃�н�������6�u��M�8����zβr��<����=r�|H6�
�A;�K�16����d`�������6)�?,V$!E��'O��C��<0��&��sùNĈ�p�r[ۤ|@��O�#�Qf=�DC�%�5�_T;�M���s����sb�S4 	=�w�i���LӍ��N�L������#���KM��u��۳m�T����W$������5���<���r�P*R�����4� �̀���o���i����m�Z�ݶE�D�� �WL���P�x$@Bd�0v�0�RΩ���2��L���j�b{���%$qp0��K@�W����M�������4*�a��� �9��A���g�3�2�����dvP\��6L���%f�O2�c7���߽3�i������2I'��P��f�M1`��5�̹�t��ڤwup�!��7�Y5J�HH|�>I�Ր%���M9���Z?���_PG8/o�����)0Jè�U-�Hi���]�ը��/ym��ԐT��\�&����J2�=��ց�m�Y��>�	M ��%R�ט,.��k�=9y�=5N����*�&���-��v�<�3�6�r��!p�g�C%�]�$G��AJ���5L�p�����,'�a7�k
^�1 �����g�v�L�Aa�d�ڮ�X��xm�0@ �� �9衴��� j6M�֣A&;���@p����/</������[oI\����df~A����R����Ȏ�)�kp�eW�K�nE�N����$��7�t���l$Ҁ�-�k�)F��֭[��q{P&�G��i[�͕eMrA�f����(�B�|�vT��	��Eɯ�K-�A�"t�mG
�����VcRR�	�]v����@�� �̇=SAu�<�C�����scT��BA+��u��'C7�YI���&	����$���Z�vN���Y�63 �!�GL�A�-������[�ڤ�T\����\��ɹ�W�&�ZGǋ����wW�������|����F3_�Mw�S�����N�	���]��t����]��"��k�	�����{c��y�Ï����������i���o���Y>*�&a��ղk�/��IS-��	��0_�jvWƆ�zo)�����(�ݣ����3��|q~tv;.'�w���ze.P��)���;�b����k�*�&
~$MI��ڵw�����-�V�h�S�N\fn��tD�x�� �e�«{$��G�������瞖��aw0.��7����=$���79ׇ���.�:j�EX�h��[0��O씲�2��\�t�R���D:rT���(d��{��?��~?,W�\�W����y���k�|M��������V�)V��,{Qz�;��d��c�
$��9M�
�u��_{��`�~��Hmz6C�z���.�ϙ��kj�C���\�0tX��{���2:|>"<N�m
�n��ۆ dm�H�H�i�������0�wxN�����>P?��D4-+�X|v�S9��g����5I쐣�<,{��5�˃�#��� 7�W5�ݔǞzX�4�J��^�,Ʌ��I�`]��.>������ko��sg%40@Ҋ��)����??d �W��1����h�ǟ]�u�$�?;Ţ��FAb�Qٿg��w\b�q�~MZh,��?�1?pr;Pæۙ�Z������[&��rkn�ڵ˷V$����P0޲���I��^w���.�El�ޙ��!�C���Aˉs���$)M��2}}A�庮q�h+�;8��'Ѳ�N�����,�f�������\��각#��uQY]miP?��pS�dX62g��D� B�8�8�oɦ>��L�K�9.�ǂ���Ȃ�cfs���M ��@�|dt��۟`6Z��-M���<{�����(��Fܪ�BhM�%���F�)YH�w�*�)�A���x��5	x�R��@����3a�_F�!��%�M�?!�q������u�sbB��1�n�zAւn!��3>�=��[�&=��$u�a�]>7���Rp\�K�HU}�g�g�ݪ�-�/e%P0��j�.�gxݙ�^�;,7n�$����qK��!=Cv�QFQ�B�y�(����!kO@G�󭍬���q��M����o�p�6#BM�P2&��r�> Np=O�>+�51����=;nv�1O=4�K��jg�	�yƨ����z���U����U��U�P��2��q����q����� ��(r��-"0{�=�vX�[M��0l������D������&�Јf�g�����C?�h��&�o�n�I�w��h��{P�oY_l��c�F,��p�H�y�~"��r��e��ʬ�h�0��k�Äj>��4Ӻ���>�j[��S't���c	un��bb>�0*��.}�>�������ݲ�^%�0�S+zp�ÄMx��y���C\0�I���� v	����,��X&vNɖ&}g�A8J����m,���v�<CgΌX����]�ڙ�0s*&6�C���L�@(U״��i�L?��ᬟ�U�8�#��HAx��Q�;��'��aLiP24��u5"�	��o(@"���n�}G���Ļ�e�e��lYҠ;[�e_|H�K�d%[�c��/_��������ū�%*� ـ��f�Hj(%��'$����+5yX"T4��-�蠮[��ׄ�! 0x��HZ�1Y^^�C�zA|������[���d2���	�<R��8P�����f�{��0n>w@*�L�;��[U���F�C���!��:�����nz�BC�cVS�$�0����3t���{v���A	�Ä~5;5IF�1b.V��7�N�&�V0dh2�D$��y�01����Rջ8w}]^���|���R�+G�yP^��K��[��{F��k̀4�(���9x� ����Euڷ�� lb ����%�b^s,�J�Da���x�%_��v��e��k?����W_������3�c�R2��P�X�
!���o�V4�~z-L�v5��q�ȅ�l�S��S���1�!��&Pjo<Nu<�Љ�>b��M���\�ř���:�h�t-���g��y��tL����	V0�E��؆�[��I��Օ��z��W���W���巾��rH���zI.^��³
DG8w���:5jVM�Q� кcߢH2wcV^{�'bi����a�J��`�#�<J{(���ef�
��&��#�yw��q��A���0a9����a���x1CZ�Mr�S�:�A�s�&�v�tB�7��bhp@�z.ke�^��i64�ɳ��W#`�Cw\MH�L2��^+�m�kG�NG׉�^�PDN�_RG?W�dyj�A��*;�B�P����-�PˮeVL��ё",�sH�Q�ꀡD�[��l�#�������*-���|E��EYXZ�'����ٿ�l�-�~r]~��2:>� 1(���N�c�L\�|Y����]G��VeayY�}�Yy�4YHI!_bB�	�7;�_���*?��5�� gΜ���$@���٧g4�s
�/n9��k
8R����,��o�Ȼ�+{��A]37���I�W��p4eݻ�s��"�Rn7�,�"� \���rD���Ƥ��v��,��2 ���Y��ݻ�����O/ɵk����Y�#��Ǣ��в�3���^���rC�x��o���dptHJM��������4���R?� ���;r��N<~�|��i�ʔd'f/��A& e-��U�59�qĵ�i��P���e��W$ú��74x��g���}S� N���c\���E�X ���O_� �-G���e��1�{������T���z�N��
�S��m�Èb�g@A�������DZ,D�G,h��2Ce�K	���f��鴺��%�f�9&�B�p�fI�!���]�ɰי��p���d�{���i�	��BU}�U���D�5�[�D}S}vK�2����U�)F�������G쒴�$H@�l�8�e����[|��JIc?�Y}&�X�*V*R�ՖX@mwL�*��R��-��%��c�������	HI�%�32����O��!)M�1��d��� d��0S:*-�����R<����~z�Ѱڹ�#?�rQ�DcT�	6��V7��)��)JT��Ĭ����pl�q���?�%���%�w��-S��|�A\nos\�ii�����$ĕH��~�P��뷊5	����!	[��{�mq�ki�$�h���(�`OC�#�v�7'L��K��uOp|�G�Ϛ��3�/�y����� m�5�1'�#��^B��T*Źx�#訃���SPmb�0��PJ��gA|�$��Z��\#A�l����@��E���c��toшr��'C�9W��Мbi閬ʺ�(�f�mfq�Ь	�yV��`*)���y�����v�adM�Qu�	�%	�(�K�n�?����G��r�q�$����ێ�=�8�L����e4����o��/v	��0�~g��f[��+�&Hr���
%Ҳ�U�������_��<.�Ԉ�׀�cc���� ��n
Bbj�; C�]���ʺ�M�9���;�/���C=��N�ï�n�&M`C,W�r��grR��׮q��Sg��W~I=t��4Θ!r�AO�+ٗL�v;k�L
��Ǉ�v�Z�l$�ݡW�UtqZ��n3��"����8��?�g���(p��nT}��%���{�e0Ѕ�Z�zX֯LS� mh�R����Ŀ�6&�B�������˳+��0'��7�^|Iv�&eh��:tTң#��m��/=GH�;�/��;-�}E�^���0Wuee�L���zTe����7��y���{���#�%Ց�)
��������U��refZ��g�4��対b��?̹ɖ��dH�����ǹGv�6]B�țJ��2"�MfUGO������cC2��IL���c,�����gj$��A��6�C\d#��x�[F#A������%���E�n����u�߱S�lT��)9��
Xt|�� �JKB��z�)��!��A����죓2���+��y������&���]�j|O��"�w�T}�����4�Rc�sɖ>��Ҋ\�6-��Ѡdf��8�jď�w�稽]en�+���ډӟRx���u�Yv���k��L=%G�� �i�х�i����>�4Z��ި�W煯!ͨ�axs�Ltq1�U��	-3$���nC�A� �H�Z��ޠ;{���4�*1=����h��g:�pr�z[&��gp�
H!LL�b��o]��\_(�UN�CC�$G�3�mK6oX+��돧���󽟝T�\���%����[	q�'u{��n{ī6�G�� q�ǟ�׆�Y��!�04���Y[N�?I=���:;uN�xRϛ_�i���������Y�e[-Cc>�?����$W���ʲ�G���8'�ق��C���G��W�JE�т���_��Т�
v6�X�nn0|l�M#��w��\c�g��N�ىR6��:�y@��#�@�G�Rv����krZ+�\��t�%��s��{⊄��ILzx\�������YRqm~E�;���J�ޡ�	�x��,�X^3׆�j����:8��a�;�Nn�4���_n�����O�	(�	W�]ͮI�����5{�|��	Ba�>H���[oɩ���@�V�Ht�y�@��jeh8��]N�c͙�4�L�M,����+��W{���#�-j�R���wTm�^]���@�&QK@��6P�M���7��l�d0xX� ��H�
h�����i��ne��q���%��m�3���j�]B��/�H�,�-[�����duyKֶޕLY�yL�j��*9i�-�@dL/d��%%2�b�"�M�5�=umI>�p��_����e�����/2��~wX����9p��q��ܼzY��u�)�`�uE��͵U3���\0�,��� "0�s�_�}_�|�oH&Q*����[r�������HJ:ޮ��2�o�DL�M���F4�P{�\_�[���`^D��G1��wq��ʈ�A?�9���$�
H|1?;{�o4p�.Y���&�i����Ȏ�ڤ�ڋ�l�dl���"��{z�9��#��a�ܶ�ٰ�(�;]��dЫg����%~;D�{��H$��uU���{�g�ym�r�#q�u#;�慳��X#ARW}��mt[gfob����嚸4��� ]�}a�s�(����i5X�o����~;�IB����G���Y��=jVi��%^pD�2�	kY�jVc#�C�qv���=K�nD�"4
�W��d�z]��˺7>�Ȁ������AR�mﾽ�g`6�vM/iQ��L����ճȦ�p�K�{�د@��J�H�sG�H>[�bYdf��k���J\����� :�;��>$Q"^�G�<��ӏ��6�IQ��!0��Z�g����~fN�}m+��5D����w�Ovh
�3���]�����3�x���L�H�j�F�y�PL=��p�5��y��5���fʒ���Xէv�? ���%X��{�^�g��3OȾ��8�[�55=/'O��b�0ϣh�v��a�[��zUy���䞻�d*�IwW��_��Zv�Wz4Yvj'�e,�X��C���kb}>Usjl&	���Jѻ�{(�����K?]���v������~�Rn���g0�͌"�Ht����-�H�\��[���у��L]�U+ ���JSt#D�5Gl=�m�B�p���$�r��y8�����Cj�]ۤ�B%�8�~����%)�1�ͱ͋�p�����h�S^,Lo(�LY�r��Z��n�J���6r	�4˰��\<��z�ҧ�%z�ɧ	cs[��#g�0�!���J>"���3�J_YX���3�p5��V���L/�K]�h��ͮa�܆����|�!tA%��R�鍷?� ���|�S�12��4$���%�ݷy��dX�u���?fd�-c�
��ey�7���+��B�033#95��U"�EgpY�Z���&�@'N�l�%��� �2�;{�s`��9N���Ы�Ghp��%P#p��}}_$w[���|Ց�;j�1��k9"�]�_�aAA���&����vjk�%S+P7w�F:�8`B�&Q��Q���EMh���HV���IB���=݁V (zOn�]jm&!��I`���8�,� :�/����E�U2<�O6-����S;ds-��o�����	>/O$G�A-�i��4�I�������������u_�Y�_C�9X͐d��A�ѫ�Pv5�;,�FɅm��tE��5M8�W5������Z��
��32E�,��(K@K3�j�;�`A�8j1�E:|H�\t�1��~��4j���R�!i�K���q��p\�>9�ϧ�9=;�W�IB�֮���ݜ�������j��Z} Ň%�X�!z/�Ǳ�ۿ� `M� �� ��I@?�2��:�?������Y�Y�-���[��CgM�N�!�� )�����My�]��%��X���济t�v���rE����{�amJ���|fS�U9t��yC�	�0:�������J�ʼ�E*M�x#��y@�#㬠�����!�pw]��O�2岞q�	�8��7u��qX=/5)��4�>�AzD_���A�vDq����htc����Y��!D����kX��լaf9��ђOO���s�5QJ��b�s=bB]�Ov;��Y܎�t��Ffu�o��m�l��	�%D٭�׏�Z�Y]Z��~�{�ge2ub���Uuu=��
��j`��0�P��е/˭�Eݯ�@}8�=�E�V��&Y�\�21��_�'C����K��=
<���NC|=���'���� D���"�즙�w�Q+-#��X1�+�7!Q��u��j�k�}��w���n���A@<G�G���%t��f���%��<(ެ�nʀ���`�̗v�HZ"�	���P0�Lw�$r~ii����8����ֆ�J>& =oD
�:�?���76C�y�PDC�M�**5��,�n<�o�lmal}����Dm6tA�f�b	������ {k�9r6u4�l�s���c�20> eM�=q=�	�w�Y����8h�9=���m���4�QZ�<c��ċ4$��2��H\���MQy���HЦ����}�P|�k�Cd�GȬ�3g�C$�63�����cA"L�`yT�n�,�X��ѩ0��2s,��ײ�A��xf��k`��[��|�޷`�м���x �s9���7��?ˬƁ`YEWR�c�DFZ��0�֪�G'�ɉ1I�U�����/��G���U���4�@Q�':��jU�n�5��;94Jd�f��q�ڴ�O��fѷ��Y��%B��@��I��/����%��q������}816&�|�5��k���&@�U��bl�����祇��q���0Q$�/~���v�;�`��[�ͥ�x)��+5,>�OT�Y��LntPY�t���D,�s1�@�4�k�E��/l'��`�$2 l��|�?��z�C�`��O��@Py�y��'9�^0�O�@����R�"�|���.\&�Ч�g��!y���I��yMfؽ���2G �2�ƣ%�-
zMz��Aၦ2X���Dt�M���K��ذ���A�5|j�Q�q"b0#�޻w���o���g1����>����'>c�24:*�������1��?����������X�^w@~�J�b�(�xL�5��D�;���|�mg]F�a�w�,�̿o7�����V3a��9w��zGt������h9���O���3��5og���8�M"�̘\����.ؼ��3�4���ec���GO���Ø��'*0�bF�?���:���LW�� �3H@��m�;>Y6 F�V���"��/����4a�J5��p2I���.p �h��An8::�@�/h-�6ͼ~8R&wz�A�/��$�Q���Jv���-����ݭ�-�TP�Z����	h �k��p�Z�s����4ys'�<���]�� ��	�b��b��_�;$E�&���c���VW2j�ݒ'K���@W��̹�L��.C��'4�MX0��v����M0��.��!�����f����z��\-4+�������wT�t`����pm�lS�#!db�b�oNh�/:@� K�b\*�;Ơ��_�OB��%u5�81�1jpI�T:'/5,kl���O.:�8C,d�B��ga�C>(��n��t���ա�m�ȥk�r�Ƃ�4k�1�����	�'!������x��K��>[� �Ju	��� ]��|Q�8�;	��F��V��tPv����g�ͩV{$ع1{���V�@�
�0li�
h7��L���Џ�
��g�Š���<�����U�(�ACD1��^=C~M����B�Q�N:Z���J��~tn[Uik�Z̮I>�a�Hjn����`?���`��;&����
fN���t-C����I�X�x�쏴&?Ǹ�Kti����e�:f�i����5����zB�;��âI5�*�u{�sc��ꀭu@??f$i��bр:�6�b$����1
���j%����h����k؄䇞K�;vKi}Y�px���S���R3��ޞ�9�u z�\^��&H��[Σ&�~�5���J�b ����Pܭ�jD��qV2��4��!��W����uii�[��)�g���p���D��l$���1�?���΢�lI:�qț@����N ; HO⑖Io�ϙnGMt��Kr�ݏ�"��7:�Cn��A��2.��"�p�$��ꙙ����oϱ�=�	'}"3�;_��4AmT���M.��i�\��އ�=�� #�yx$���A���s�^[aT�˚�^��A`$!&=�ם�:"�$�aU�	�C!H�y-H߸1v���@zP��~МIG����R��k��l�W#=h���7A����9"��_$�
�]X?[�*���<��S288ș$~)]���ܸ���.@d�b4���Sr��r��ɰ�F�V�V���NȲ���lY�gI�����!I�$��Dm�ilG�۬�a�u�eF\0Smf~]�A��pS��M�_�����Q�����q$Ö}{����!��-
�{\x~�|���d_�:�z�6�*����^�1g�b��A��G�矐�(X�1;�9t�M�j`�1/
��C���ؐ|xn��5j��m��ܘSA��e{\(����0O�	7��!���{��G� �v��̨F�������hR�����Q��� },�=���O�c�>J�V�Ӭv"�W򆜿2#^��ф�^M�]^3a�;���wv_w�2�}�t�t��D�p��6�qd��Ե�U�!���z�(c���s����],FC~�ߢ���B$�k��l�|�A<����������OH�l��� ����$��=�Л+U��+rK�FH�CHAg� ���D7��'�9X=�S{�䞣���ų������T;�����ˣ�<&#��2�0G�x&&��?}]VVV��b9Y`5ΰ�߻��y��{	~j�/�J0�+ח	�:M��/��{�E��-�9�0]\�a�'w��kg�;�mdW��h5_d��}�m�o��z�,�^�.�q��9ƃ�n��S�]�cc�߯��_��	�u��߸2�l��xC<@� �����*|�������.3`�9=w5 A�hy�m�h��H�"I�GnMdu��K��ƨL~�X�j�Dt@B�d<z��+��C�!���=('>�L���5=������Lf]�,�7g��73[҂t�~�Ω}2����k� ��5�W�M��۷��V�g�r�P�,�G�S���3����~���w���:�a���������_�,�;�4�m�Lt�>���S�p+p�hW&�jV��'�
Ґ�Q)#>U� g�J��u�'�ֆ�G�CgDh�!j�
��}j(9˦!
|v8��l���Z�I
i�)�� ���ã��OM��{��`�1����"��Vh��!�%o���Ar�P�����Ag��w�%�=5��\!	E���Z�ty��DQ݈KL:�j�P��|G.[�n\����غ��W"�%��m����c*b�:``���!$1Z6t`�j�"���Y�vU�đd�F���<�`���$�~9H[>6>ιN��=Fo���#�R�{�����$d�ձ������\N��1 ���4�-;�w>$�Y�ߐ�W�_���f���ge{�jp�Q4T��*�z۳]s�LACQקA�-�}�x���3�'+�Jj��!��#���!Q^���4�KkےM� �[u5p�1X�UZL܀��l�$�ii��NQ�C]-��oq#B�c��o���*;��]�¬�XR�$�&��F�f�s�<��]���Wc��M�c��#��S��u��V�\1�utM�h:wQ�X�ˍ+פT,�Kn$fezr|L��:8#a�9�������u&bЖ{Dy`o3�W�� M�&����������:l�&��4�+أC#ܳ��@
��7� �G.��l�gķ�Iٻw/��i���@���s��y��Is��d�C�*�Z[�Q��|��95.�g��9Sz��3@�d���<43��i�����$v�5*-�<�	�B�����_�ͯ˃<L��B�H��� �f��4
jjj�^����5Y��#'������ȗ^xZvO�S���/h���$ka�M* 5j
҇����!AF=����;���p�Z��@F¯a]3���&Eu�E��,j���-x��ge��]$� �����i�����\�x�6�,�nӡÙCm߁r��dlx�3� �����������Pm~S֖V��G�ȞC��u�8mS-�c�8̿=��%��s�DN�ab? �ӥ.�m6>�Vie�^o| �YCb�9z�����=)`Gw����f�:��]��6��o�;�ɉ3zI^!��S����?�=���Mhn[�T1��d�h�a_����JY�=�Wz~ڶa�E�?��:v\�����ڦH�z��1BF��54������Gf*x8��t�l������\�J\G�@�k�I�s�^y��g�(����؟�䠮U�I�'F��b-�)�m�+�1�$&�p䫜r�)���LҮ~�BM6���C瑄b�/|�*��l|�-v[�������4,p��BHj)�>=��r�"�I3��C#2u(/���8�������!_+L6�U�k���ם ,�������4�rnnI�_[&�4J������1���rB��S@���,�F��\X�΃>$�Ԁ�jЙ��[�g��)��!��):���_��ܦ҇&ԮA[��#w�%���\��H�������<m�7$�	W@�#�s�����|�چ>�?���:�D��2�<��A��C��>����y��U9��p�/a�U�j�}�ո�Ǝ�����sY��	��><�k4jrsyC���^����@T��#�j�q'
�y�w}_��Av���W�C�.㸮��"|�j�0�bvb`@�?vLba�,,.���:?�$AW+�U���"eб�%�$���s��!�j3�9����R�wmqE:C]N|�-�H&��5�c,$_S{��=��?$1�Orjw�m{[Ĝ	ۉ��>����v\o�.-cW?#qȅ,#} {B~�o��i��>�(כy��X��Q����-6��	]Z�x�)MT�~����*3���o�daz�0� :��K�P��\P	�K ��J�C1}Q9{�G�Z�;���x���z0��h�V��Ɩ=�qAI����!#����$���0�\9�T[�q��V;9��	
�N}&.�������?��ܼ9/�|I�j�b�<�����#������L��5�l���mxk;��W8��3H5۾yX�	�A�l'����~R��!9�����]G�T;[�w[�Yl�h�s�M�;��Q� ,�9`��t��6��`��=��Ú\�K}p5V0��gD��Y{���*7u�^�m���5h@Uv��}����Ȏ�Ԛ�S0�"�A��&�h:↭���>xXJz��m�N��0+��f`�5+�dPP�G2*�`TÌ!�6�v���b@ʥ2zXf�;����r��5GʠCȅ�g��mC<82.;&wi�d �����L�w���L��
�nnl��3��弛M�����	��>�}���g���]'��l1�:��[H@���e���@�@������;\L~-j�7��[�Y��9���n]sI26QT2W���(���� Y�6���@��%"�	�h")��&օ��&�5u�Qo���qI���|���A��漜��@�s"�젪j��@r��"�(���ĸ9tP�G��<k�K��z�������T��uu��An�y�iu1v�Ͷ�ҽ��������s����k�0;�	a[�n@�~W��;�@_�]�Ebg𬰶��Թ��r�w,��PH_��ƞ��m��V����u���v8�~��$ �oȳ_|^����d���V@���8Й	�<~Ϝ�)����r���� g�Ԥ����jKԧ�2H$
Ilr�?au��n�lP��C��>�ja�	���ǜS�X�FG/�$�p�=��dxx��θ�ݻwS$���dh3"�M3���m�� j@��cr���߿o�>�a�?򸌌��dƒ��gd�֊��ǆՁ�X��Äb���2Sc�I�!��H�)`���7,��"o�9߄�Kꈢ�B�7&eM�2Ś��@r��nś� �l#X��g�`i���٦\��)ã#��=�O��+�&Ã���z��d��p1���!a�� ��?�Px}]y��,��k�6H���V��{j{�bk ���Ez�X\���C����^y��_�x<!��^�|�������,�ʵ3|>����>6:�4���Ok21 U����!QX�l�����_���{�����ecyQ�����w;���nC�t���Ȣ\ŝѫ����^����-��:�Y�A�9D�������l^�Q)݁n���*���� aRkV؁�ۗum���d[�wT�Gx(�}�o�u�%�����&XFQ��7eT�/h��jP���ɲ�I��Jh`�4#��h,/��.)w��<��ܨ&�ò��>&#`F�Z�d��~+�q]��,��z�Em1H^!	�����`,�ι�g��`��)�ܓ�L�"'/]g ITɶ 3;��߷]��=�� o,s�`�e�Ν��\)| �V�(֕����m�[����ټ�{���`p \�lf� m`��V�X,,I����?,�#�&9���[��W��R*���h�:�[�A�F[�"�#  ��{ǥ�+��M�3=0A�<�~J��M��>��o$J((�l��Or_��Zc����e��BG	�ݹ�����Ht��711���$����g�P�[�K,�Sd�$j*����d�n�/��NMZn7>��������GX�O��e����̷Yy=�kA@�ش�6��m�p��h �>Oﱡ�	�,M��M�M3)o;�U��7g�M���H�&����ޚ�y҄�E�*'��e
I,����|�T
�n�Tp^j67�&�L�i��*=�O<�$%���P.U�����G4��$�����_\�\,���<���r��U9��F�V�%��ZכUvjQ��1�G�:,��ޔ��5���%��9N���b�3�@�z��-�=Fsg9��2�v?!/�E(�a`oҮ�;
[ﱼ�g�hGvuAJ9�gE0&pb l�I��@��nK��0��8@K{��[�S��� I��yW@V�IP?>�1wrdLυiD4���h�fL�eq�4�����Z��~�7�k����̗���]��L"ѝ	X�AS(�YXM�hlӒ�1p=��97��y�S2}�!�YV�VeaqYl���Q	@W��J<9.���X8�iԃS
��������tG~{����wc�/������yn\�YEYY�>/3�_�e�љPL�[Ɓ�Y�A�~
��c5�>&�v@C��B7 F�,�nښyk����g�%�׌zp��*�� xl���2د�I��P�j��2�sYFM�Fb��8�_��!��3
|�m��?m� $VM<T�zY+T��̼�4 @�p�<��D蠼n��jz���vY�hK�	T�W��a*�L˽��##RР�������r��c������9�b!�#+�!�	���w��:r�G���޷[�ˤ�.���fR���ӋԢA���OD�%�~eՠC��.F�@g9��������`��PRd�&l��Es�HI�ӓO.�K���n�ȐzH�6�F�L���8����Р�ɥ	�������Qϫ�����Dz\|C  �S�PӬ�����\�1��:d z����#�+ ���1�d����>���IQ���E�[��g��ݲw�~�䓓LI%�k��s2.?�#��0l�C�K����Hˣ?DF�U�W����Y5���9�p�Hvl��E! ����^��]�ab>7�5�BB�\��40��Q��01�XG �"��cA�-K����w_����$�I���ԯ߇�/Uˤ�_���W򹒮ݨ}(ɽ�� ��7?�@���Q9�q������A�:�_Գ��U��|E�ъ:���L[��u���{��� �2���5I����L횒�������L��F%��![[9&�]��� �����z_���lX��Z�"���W���?�6i��p��.�d�u�%bO�.S�4m�ԞckAh���͹�&�����ք�n�������يr��$(�Ϟ;'��Kb5�R� ��H(�χm�h�81X��y��±�&J���;�л+[[�o���9�X�`>��IZ�)�Ԋ�"� �k%����Ұ}zձ�^c>
]ڊ 4`�AoP��&�S�JK(��fx�z����ր�X,��ZRۈ��E®�۲�$ �}�9n�gɻ%&*�TZ�w��r�ړ������]_orD���8:������n{C��Mnwy��>�sn��mbo��AZ9�ͱ����Sg����3^]��:�i~�ǀ���u�OQpC���I\�kdxRFF���!�.v�
H��g}>�{�c���T4)i0���)%Dֳ�C��vHO��am��y9H!<8�z~a[�����buqx,S?��7��EM�!7����F��,k�y�b���5��]���рt���kk����h��|.�Yjz!��~=#���`�-��X��#7p@(���玿2I�϶��=�.�_�4�%&�!�t�dRz�a=�DR}wV�2�Ҭ�mF���jP��P��w�����nmH(��K�����,�6��[g"�LI�@[�DE�=�32[y�J�1h�~�~Mi����A6
�����0Lw��M$��h����݄o�Z���2&c�1��9s�����0�q��y&HQ�Kk,��O��¢\�rEnܜ���=��6Y ��_��_yE���?��E��ӹs�H��D,Ō��N�g;��&����0��2㨅�P��`��9,��'���M̙��b~S ā��\�=��R-g��� O�H �/ ���X ��ev�Lq�srHu�$�G�-��i�����yNl�F� �D��[����\�ʥ�W�V�Ⱦ�{�˿�"�A�33$�:{���������چ,��HA�'�qHjǤ�SM0��\�0��4�+�����7m�����r�cr�Cw��g�����zƽ��@�Y{�c��2̤��q;	���os"Fqbƞ�GR����(�Pb�����C^#^W�r;iOC�����`*U����&U�}���U�M�%[n����,..��m�S��k:�=3�Dxd��_�E�2�x-m�d��`l��PcN/��(��A�j�(���D.4:!&F���)i���ϩ�\�}����<�ܳ,��ާ���Oe�$���P: �^K�:�g�E=S��OOɥ��51��xjP���Wd���������}_�]��i��b���u��\N�n�w��6Q�mm��8��gf�y�����~�ן!����m�h����_L.q����y���Ӱt�K&�_��W���eBG�Kݓ��`��fhi3+�����*���So[���KA��>��36~W ��e|�]�#�V�z�%��iB�P�]�Eq�6�ཫ�+�w��T1� �M��N��hG�,���E� H�[7wK���]:�dzX��ը�ХP��r�瀹���Zh{;�βS�N~pdL���4Ȫr60i�ہ/��T:`<�)HH=��U��k�L�6����W~no�;+v����5��4��h WO���&FC�β�Z�)���H�Z59~�:����9�K� �^s]�̎Eu=d��Ȟ��Ch���g�vn)+7�PC�`���;@*�(u���P��BQJz�U\{$Ι)��\@�����:����#�X3G}�-0��ϗ8�����g����H�P���Q>�Z�ͺX�2l� ���+hP���X���]RG�=ը���JF9�_��+�2��m�a.Тc���Q����n��1��k�.;B0�H�=�+�$p�&�8znv0]n?�/�$���+��ON�V�_b��1�p�g]6TF�Ő8�(��a�!I�GE�}MB*R���{?}��]��&�s��#��i�Ð5(�mz�I	��� E!�;��x�W�� u�(��`,�]���j���zcFbuq�s�9]�����Dw��g�M'8�)Sc�-=��FU�M�5H�`�ʥ+����G}�N����h\�$�7�:����C��\ԔD�`�u�#�I�2�O����"��KfS�w�J�x 'Z$-�D��v�t��khhX���ll,i2X��: �(�m6lŲ(� H��,��JP����>�L.�5��}.��	%I�F�?�"
hnɗ�h��5����d=_�{0������t���zZ�PܰY-�� �c���é�D�/�9��PP�)M_�!���>g$��@�{`���ڈ�Bt�ϟ�ȢF`676���#���/Pgl,�1a4lC6�u��2A��3C���_�mVȲ���@�>����yRe~����
?����P���(h >�AQ��kY#2��s�m�z-�k2׭��@��0���[0ς�t�����5v�p&1oY�f��a�1o�<h�P�`rXo?l�4� ���vx]7�V��"f찞(<4�>3�5�\�;,������DF�Yu{������OYΟ�ƌ����OO�G7��t�����W��r���4y�	��pn�eTe�u���Xز�[{�a�KN��ϖ��̲��E��x��d�:�5$g=�u��i��YX���kR�Z���	�Iݧ a!s(8
�3�A?�0-�#.~*�T��`�ĩq�M� Ao5%<�"#4��'d������ī<�]�z��G�D�>�@�1 v��۲�Ϣ+!�m8Z��h��xky�>�ч!3�������k����ax]�[���%�� ��,	�t/B�nxd\n,,kB8-�z�h��P�djOS�Ӏ�?xD�Hn�$���z�V�r:��S[N����9�/�?�3h ;�2<�xX�iӇ��1I{'�[�$��Z���`�Y?EG�b�>c�]����S�Ok��8khx�z�{'�dr!z	$�B1�k�gXw"�k;�KrenU2�^�,a����,`n�Uz���v�x��x�������4y۔'OJ  taq�dG�&w���v��t�P8�z�G&w2	]L� �i��[Z]�h���)��'5��,'�\���7SBqv��o�0��,��tʱΞ�C�����=Cgƶ�!�7�M��6.�9���+�:������`�~q鵇����=�Q_y8�xږ�Ѱ���,���O?�v7t^��k|��_~I���^r:�d���ߣ�!�I�B�����!&5�ֲ(��,�&�&�j�_����k۷g��گ������eY�z�MYX��p<D���/>K��խ����9�|,>#F���4�n��W�<���A��>��r������|I��\|㤼��'�O��C��'�3�LѸ���֡8��?������򲝻�����a����6�rO�y>Vd�?������۝?�+nnB ;�9g#<�y,&���2t�d1C�H3���lz8�MЫ[�$�(4:�Щ��Lc�{�p����a&P�@t�����ں�U����a�t�ո�4`N��#H,��+H-?@�ܖ���H��)Zl�#�����E*��u�$!YEU	�{�Nȵ��8��j�SE�X��%�-��l�7gg�0h�i�S���9�\a���� )�{\s�':r�]�F~�g���ǐ�t�?eSt�	��h)�@�m�NDp�ǐ`����sz��Ŝ���4�ΉnYP�*L�V�YH;_XsZ�z�A�R��P�\�A@���aM����Vǡ�n-V4�q"��)�{�1p�m 浺V�M�e3�G-�T�HN�+@�0�@ ���ƍ9��Ď]|���v����"����7�f�0�֑-�U>��1M����A�Qq«@�ԫsF,��HX�`H�J$>��q$����i0�Inlq��c�;�s��������Ǻ���ĕ�9�3գ�pD7�l���,,tjeI�"$"���o�K��n��,mq^��d��C��c%v���m�q�zC[���ًj8����uLpM�0������}��t�73!�s�^�@�����n���͛��@��~O�9�D$�z��9�������;2;�$;w���"Ã#����3/�ǀ�wz	�P��T�)Y�]n��+���� m�[[���͘:�v�A�
���XaEE0Pt!jj[��l����.nj2蒊�;�rC��b0�{k���4��c��4�NϚ�.���z�D*E�=��Y���	���a��bn:6<�"Q�ͮ頡�f����6^���/.�jB�S�р9��[2����Q&�37feC�b<����tɡ����T��|�ϙy�y �
�7nܤ���}�����{D~����8uE�g�M �yܠ5���ř5]1�=bEM�	���?L��nΟ],���}Gq�b��'����	�Mܢg�^�j~M��zo��7��X��!�G���E���u�?{��]�8����'�A�R����XX��W5�hɮ�Iv�P�H�Gexǔ��4�MV�ShT�ϐ�u͜3:%A���!M����9t���3��RMxL��g'?�,.ٺ�m2Ѕ����<e���3�BA�T������?��q	�>�Z%��}Z
����ڛr���|ԇ"�@!�q bt�	����CYwY�b
�&�&�X'$�.�H�-Nq�����B=�!�{@�~�!I�^����j�M��#r�ƚ�b�P{�P������3�ɷ��?I��������~�k����i�ݒ����0���d#S� Xt��B������	�ś9q���oYmd��$"�o�P�j�m�#�Z ��
��Z������y����yD��npӚ$���Y�����]�D�����å�5���م�E�$6i���?������=#�x\��t:zwv.�� v��^1�1��ƞ;�x�u��عwD�	�p��qC�Z'T�ޣG侽K����5 �@���r���;��>�622�����Y�%rhbH�}�a��~6M�	MB�J�$epxT��"و!I����y�P�F-�Y�����Z�IQ �mj(�?Ӗ�N]��[��oڊF�C8iP��s�?'%=O��o�Y�l����@,)u�(�ϟ�|6�M8'Y=G��]�]��N��|tF�\�.]_Lݧ�K��M�sl�)�0��L���!|����tu�cf����L���X����k�19&����;:���ƶu�x�U�˳�i�5+d7uC�q0�1�������x5�K%	�r��<��Ii3lk�Pa�: X�>������'HR��3ɮ����5)h��A\qK���Pat�d���`��Uti�8/f���윚�W~�k���O0�׳a�D8�h�C�gImlM?���M��������}�>����o�H�5I]���{J�N����]��W�3�0�H<�ukxV�Xj���(?�}9KA���<�m#m{;D�����c����o����>�1f�m�ݦ��s�+�� `�a��Po�/F0���=�S!�m��!��A^u�v���Q��H7��^��"y�n:wt%4#)����a�#1E�h�5���~&��|�)40��d�?��ؖ;H�B2�����Nan~!�ٵg��3���ZH�*m�!��~���Nyꩧdsm�.�H�54�X��,葍����꯾Bqᅅ%�X��F���~��t��B��I�	ސ��!����p @c�v m��%1����GB�q�{T��.�p�C���W��C�ш�� ��!['�{����*4��&"l� �����-�X(��1�����.j����&Wu���_�sO���Af�9DM�C��dKM���po�:j01gv��]F'�ot%��Ñ��29�K��n�V6�g��4`��W��u=13r��Y:��s�LbA����R]*8F$Fã��_��U������_���P$@J�:j�A�|��6����qN,����rj��9gN������C��r�,g�X�w��3�S���`������%5ԛ��=W��ni`��(��CL��\���dr@J�*���n�Z�����wk���q�̣�%t�� ��\Xkܶ�Iu��IU��r�ř��^�� �9shB� �bm�n	
�R���5}�빜d6�$4����aT����c��tDm����5��DP�d0�v�+�G6W7䮣���_��N��\����������	�.�"�7�&\*e�njU"���lS��m&�.$��"��9C�4����f����1q5���/<��muFyMb39M��9g�mUI�SI�u��D~��)�y�:8M:��2v�|����PJ�[)lmh"��`8Ȯ6P1jֵeU[,="��ȅ�[dlrHr�X 	�d�լ�yέ�,���-g��	KQﱺ�$�>���\��ф/64��I�&8��: �v�#Y��P�@6�z[FF&9;����LN�9��<�kuJ��5�r}Z>9u֐��P��~�C[ѡ]A,C���FȢ�:�謠�E��j�>3g���ѳY����a}΀c�H	�������4��ozSi����nz��X��``�J�DR�!�j�ܕv��~ll�XIԊ2��C `f0��N��.�mf���{�y_V�0��bU�FuOwe��}��wϽ�C��H[������Z_{ݖf�l�ˎnבH��7��D*���J���[O�X�����;th����#.Q�@�;���	�\GD>|��v������$�k�z��^��:g�J6�����)�̸!H��@|%���Nҟ.kO<���Z�v��=&����y����G��>�ڒ���_��D���-c��S笣gU��.�I1���em8�{�%$�K6>��.;b�t�(��d���Q�k��Z��;]<�I��0i�L�?	�5��9r^Y�2�-�,!A1EfB>%ׅ��u����q��=��ĵ��X{[8z%�����uR���n�=ø�4�5؏k ��Hf�m�ZVŭH b	 �%��*b ��R�a�y���PO�]��[{���?s�:�:43�Y�jƛ{��9�ű���~9�=p��(�Ǐ�fM\��?�x�M��F\Q�g����v�_��h�,����S'�VRg�_�v�2���VX��[w'hM�e��5���+�~��v��i�0I�O����Z�x�k�37}�p,cpE.�=�<".P��I)/A?>��[�*�#��ST�����LG��H��^��򔹙E�������+ʇ��!�K��c�`����YW[R���F�,�����¶V���1?�Yߦs��I�K�'���/��/���N{�/���q��Q�Xo�&�|P��s澥��2��v�IШ[nkՖW���1��'�'����܇��(�,�FBT٧G �AoX2vU�f�f�w}ȩJv��e�Z\F�Y��ײ�֖���O9�
�⁆��A�����s��iOb��̝oMOЧ��|�"~�Q@}�P�
gk�W�)���ە�U���]8o'�|]��	\���c���Q�>��>\���&��Za�fW�mqqVq&Ց�*�ί��m)h7�o�F�Gmce�f&���-#�<�n�r�XV�-�^�-͙�[����yKE8�����^�=��u{�o��"�(�-�8��&��AĹW/^���e�6A�����쳗Μ�o|�g��ĔY,em��x����D�7��\����P�s��	�o��v1]�릵D��.0�N����D�_�rb%<�/הP3)w^]�'%VY9��K3V&K�r48 psn��� v+j�-�1��{���s�Ve�O�DfaE.jj���>,�;��;u�-[[[���z�=�M���w$K�JĔ|�R��j����<�̓6���7O_�Rm[�z�p �$�%4ă���k�	l�!�'���l�-�V��3���a�q���q� �
i`�@�M(�.���މ2-�<�<RO����HV�U�����UWc�#&Z�O ��>)�8�+�d�����NU��UR5��`>�L>�צֳ��V�����5��j�d5|�[n?b������Մ�{i�&)輌�HU!��������?k�-�H0����'>j��Y1��=Z�NL�(�"_�3%}n|XJ9<�S�/!�\�H<e�d�T�De��g����h�=RN4G�@Zt��8Ĝ��L������<$�(�C����\�8h�֮�܇��E��o|㛖Τ4@f����f�X���c�-��O���|�̠��ތ���\�<ld>�+A 0�@���Y�`�y�M�Z���'U��%��U;4���}�I���ׁlsu5缠�@�κMV�5�~�K��*ٟ����?����-��ew�~���w� "�-�&�7��<7X��%գeWp�|a#g��ɋv���������bn���@1�q-"�iv�e��|l�ƴ:�t���N���u{���k�H\V�6I�[V�H������{L��l�\���H�����oe%A�XZU�g�< ���݁��T�8"~�8�S>L�/�romm� ��e�CG��j�;!V��G� &��m#�Vs� �����',�Y�Q\�Ie��hP���[L�(v�|f�� U�ިc�&K�A{ꣿ�=WGLB4�����U���"^s*���b�f_����oY����(�|\A� ��?�0��X�*F��H���7g�ا���q{�3���˗���(�,�V�F�27<^i�K��;��n��9z�ݢ���z���Xc;6��hkx^M<"k�L�f�92��(wUT/�ל�5����'�P��j[[��X@�����xa"[�)j�%�4r�!( bRg�!��ʛ��oG�W�~x̊�����ß �oXw?�K]�ҫ��L&c�X�~�7>-?��g���������J~~�l6�X=11.�e>7_������ᮌ͵-"�J���SE2��HL�ݫ<�6
1��~�tX fvfIRF�}� J�=ÞH�:m������ᾦ.X���g��a���z�tZ$�.�D6��(�U��8�S�`�fO�����(�$Zu�)�]�3�V@��`��D� R�b8���4�K��,��L��d0�nˎ&����g7�Z۱�����H����e��~��QuPϜ<#
�&�a@��.�GG���vĭ=�^��v�X���a�<�����S'qov�w�}c��l��^����WoZ���;d��{�k�U7��IG�eT\NՐ���Ӷ+�	Pt�G�.#v`���<@C�V�d�˺�����k�3Np�0�XF��=i���{�����Y��w�g�o=.������ٶ��m��,�� 	0H�SN�*�c��EٲH\�/q�*}�<��b�����Ѥ�����i�)�`���uGmn��ϕ5N��"W�NO�.�?g�i/gC=}֝�P�ܢfY�'F��Ygw���<��(a�E�|��~ܧE���p�So����2 k���_}�.�,h��O<�����^�~k;k9�G�e՗�ă8�X���3���!���?�Ӓ�ZU�)$ˡ<΍����� ��.�>��+��{	w��'��e�x�!������n����=��Ӷ2�	�0J��[��ǵR�+;�J춲,���"�?���(��g��"W�f~�p����KM��=Z�޶H3�|�92��`��+8@+m5͟�ݻ׆���{ou]I�+^g�/_�js����&�|�4~~��;q�<Y8o�%J��쉩��|q{?n �i�wv��o�Z��WKU>4b�4�,�!�Eq!Wٶs�v���a�7�3JÂ�����1��ͼe:����p��Hxl[��b�*��/޺`k;~5�^{������\��=c!`�d{�����Y��7�I�����Zh�5��U]��h���HHN<_�����h�y����;;�������Au=e!�Nx4CV_L���S��̂d^j9K2�~@,S<6+n�z�?�P�,������)+�.���צ�-�@��H�]��R:'�r+W�ɋ;��-���M�Ml_ ˿+ ��BnS���ڞ�v�;�q����=4j7�l�Ɣ-!	�@�+^�ϩ9���f��{������;ﴎLV4�i B��H���=P��K�/����Tָ�X�!�X��F}��a����v;s��}��߶W_}E��u��*��I=�����ЅTD8O0�GAdu��R͛�=E@E���Lr���w]�p��N��� � ����OB&�G{;�G�BPZŵ�4�p��9ˤ�\;���%E�U{}�ڙBbY�p6d[�-�����k��6,��&I�9m!Q�[�;)��� G��l�R3dw��k��`3HX� B)lpzǴq���
$�++k��m�?�t�Oo�������AϮ��2���g	�d��3����w�P�j&��oкم�����q���W�u��}�ON!a]����j){LHZc��6�ڮ� ���{��v! %E� u��"J���a�M�Ū��L~�'�P�a�D[��s�1k��cݓ&s��i�V���ݍ�a��E�,��t�q��'ɭODCF�Q�Ȱ�H:$��7�ƽì��<hGO�7Of��m�Nw��xT^r�}n��i�^�����llO[_�0�C�3Gb9<<���jq$f�)���@O�� �I�E���$�T@� �dL�X2'��[�Ϫ�N��V� �C#�n �(�++��ssu�4�%bd��z2�K�C�B>)$�Q��+�!)n���b71���t��Uz`�0���T(#	��{�^?w�b&C��?�*�Ӫ��;i������v�:O���%kO�I���׹x��}i�_ٙ�޴��Y˴Q�mG���#cFc��^yE��=}}��������ڨ�����@�C
�;2=gw���O�����$�����B����伥8+�g17�f�Ϝ�k�&����)$i���,�.����O ��N,�P����J����{P�镗^�Z1����a׽��s��@Z]�% <{�)!��^}��|s@��Q%�] =��]Rѥ�N9K�\Q<?���f,�'��k����̬���M���~����OZ�R�s�x��T����H؏��6[__��}��V�ܴ=8'������oSSS�؇���2������gS����-gW-j���߲O�}����6?q��s���Y���CLԛLґ$�+R�����5��3?�ӧO[Wg�Ψ|&+� 7��˶��$�2�4��T��֫�3�8�����G?����r�^{�Wv��<gο7%4���h"#*dMĳ���i��X\�|?��� hf!���E2t�)m��B�Z�vr����j8�cv��3~�iK��o}]]��E;�0Q��v���q{��{���ƍ	��:;Ҷg��x��_xͮ�;cQ�< DO����v�����Դ,u�1�uá#���'_����>kx����s�V��q� ��D�ygC��d󼭺�Vɭ;�$��+��O��<�ˆ:��]�P���}�r��2Z�p6�G%���S������7 x�=��CJ~/\���w��φ�E،[(م?���l#M��;����9�����X��&����z�̭Jh��A�t#���T_El���x�5ba�j�Y�/�kb�
��#������{�[o�'��[λ��{��8�FblX�$�S.���;h��r���ͣǣLn�`|z�2�)h'�s�3�*�!���s-�+pf�x�߼�*������̐�p�?��WR��+��D�[ ��4�̯^ǚ=�_,���K�q��J��r]��P:am�����slurɖ(E�`\���������L��=��J��� S��B���ɾI�-��w�@K" "�d2�����g.O
z"��M��ke��Q��q�{�q܏�si#og�8��[�O>�1{�#��XO�z�a�v @{�=��s<���qK�����e#{��̣P���Ky�XYSў 1!���yK�j#�eۭĦ�/�\Х�^���X��d��єr%�|�
,"�DB����^E�Q�����V^�.�X!���dE��;4"��'߶��K�X_ec񦣷 =a�c~5<��U����h�f���w��r��/������;��_��o�jh���憎]ռ��Ԥh��gC��w}nFc7��6n$v x#�o�����B;>~�fǯ؞=#���}ݦ&&e�Й��,��#�v���+jХs�����ıS]�<�s����f�u�X�[��>ۻo��虳�5w�=��~������}��"Hj1]����iO�b�Ͱ9 S LeS�o�а聃HXY�a�z`pP	���v���ͤXp�J� [5�/b�,[o�
��v�}�MEtN�����
�� �6�6`7��a��@ge`K�|v���� ��PS�R���1lp��I���7�wv՚g|��ks��|�׷��?y�n=~�Ξ9c_��7T��琐����w}������޿�� ��M$tU���V�:=q����h͆�{��'���W^���%���;��'����w[�U�:gN�~ �jC��ERX�����+�u#QkM9p��s%�)|��L�k��jMP��F��%|��51=o��ع����x�--."P��<9�Oԃ���8�p[JrյfP�v�/.�i����l������\R�y�Ƃ���&�*�쨑S��S~dŶ)������W�}��p/�����@R�Tl�cO���A8����k��M��~QI�3 �Ã�6y�]�t��K�J��M�^��^�������?��p �CK��,V���C�^k�^���D�*q� �6d�N�A���9\F�H�( ց��1�<���ҙ�:�RE3��aa7d;��dm��6��H�u����l��reU�	J�m��2�%��'KW@!ݶ�tT	�5�Q6͚�S�2���T�6���ݗ���(��a���I� +�����\U���Ho���W >	Ē��[#��O�^}�ā%�b=v섽����2����=w�ڳYۻw�}���ۡ}{�����������;�g��CG���K�������I[X\����>|���V����[���1a� ��X�(nM��f�$�������]����;=��f��^	,j�m����,��ߪ���R8����WoXdj^Tё�I{߸v�._�a�[ۢ��*��{$vC J1
Fi~���kIXIdd1|5ǈ{�j���XXiTU��`��7���3��:�d[ |������v�^���>KG�� ��r����v��3O}Z�.ϫ��~Uu�	�՝X\xٔG�nK�62�c���'��#+:E���KQ�o_������Ͻ����am���mL\����-�B���>/"��R�>�3q�'�m����籉�q��_�`�����צf���$�F_YΩ��K�1A|��G����,b���^�����׷mrf1�6�i����f"me<���u�y��A�ER��؏�q*���b�6���t`l������ҩ�@<�4�>@��V@I~��6�&b��Vvꭥ���4]�(۵�W��c�l����Ú)�=�,tU�,��m�Z��9�8������=dx��b>w�GH��6=��.&i�G��R	=ب��ǽ�8��,4ۗMI�����6q�$�Դ��e[{�%)�� D�;E��B�Fbp��]�T��@�O�9��pT���q֑Mz s�t~iݞ�����ܬ��m�ܫ@ɲ�}�¾�gqV�~Yc�^q,��`̣�R�jw�sԎ����!�5m����_�p�gw�y���u�r �o_X��.���ĭ#*����^�S�.��ڒEڂ�w׼�$���3'��=xd�z���W��ԉͭ[X�����!�Q��X��B�U>�xK�$	j�+�DO��s��RoY�pOK
Ϧ�$m3�*�Du�F����xUJ�x=��"&^���$;�~g+�Y��/"[1���!�[�py�oo�����@��z�m��>[�Yx��s�Ú3�X"��[���2 #U\kE�h�|-�#	��y����|�f�� bGH̉����_���Q�C���Δ%R![����'��=k��w@Bw�*��Җ]���f�y811.�% �WF�X���ą����k�:�lK�S���<<Y��()�!u�9�]ƺ.:�2!��b��w��\o^�����Pך��ĺ���?Q��o��*\�5=�ʆ���b,�\�@�i�A�}ұ�8�.�C0\�LU��~KD�� �vt�v*�,�V���JTonjF����=}V�ޣ�;�eZv9�j1=[vU�~�������7��]0��4��^1v��j�}_jU�ץ\7�x(��`VҨ�(�jU����]��)h`��<���*%���g���m&Ƨ��s���tᒔ����n����58<lG��u$�@����ZTTw��h�=#�H���'�:�����J�zT���3O˺�mj	�	�3�C5g+W-�\SR�J�8������w64̯&-@B��Sg��Č---Y �
�VR)�b�l�5w#ʩ��U����0�ٻ�ߒJ�w��:$�䥋���-ί!(Ġ� ���4� S3I��A_ʊ�.�N U�؉lV�tI�sr�C i�O��R�)!��7k�,��I{�96@<�4	\����& ��o����`$`]��v���+�om�r���C�� c~v�~����@w�!��t��*�]@�_+o��=���������F��W�fׯNY_'6�Fl��po��e+�m�&���9Gln͟V�V�PB�e%�s9/���<���$�&��3��!���a�xV�TܔG�����k��������嫶�gD�84J:�^*����3򌤶O �n�l��<�hO"**$�GK�[�
\MT&dt��h{<��.�.���WUe���T�YQ�w��+j��&5���B: 5���qP/p�Ϭ��a �=�я>��	�fE�DU����!�a�߶��q����у����>`��s���F/���N$�S��+����f3*8x!ă��-�Cj�U�h�FE��DM$[�Q�5JRp-m �����L.�c��뒕D$*b!85�D�-QuVQ��B+Q�bƶ��� c�";M<�[CBD��搄ǳH�ۘ���Ķ��×)5�{UWB>�>䨨xf�m���Ɏ���5��SѨ�RI$�ͳ�NĀ�����Q�c�5��Hte���Nu���ﶧ>�!Qy�IUdW�󲯾A�x!�n�&&���A��Q�Ϳ�IܷOZE,���LX�^CB���q ✞��Ż��K�G|d�B/��-������j�1���m�mnbɦ��ڇ,|Ip�LM΅T}u{	��?�\ t;aA'�C�;�{x�	,x�ڐ�mڏ�y����O�jm @翓���c� �mH��,.�ú7�Ӽz��M�]��D~m}@oN���&��(�B*������33�A�b����.���p�X<��Z"ۚ�.-/Xue��[�/""=���'������0Π'�������e�v�lv�{T,��oȇ���J�4=n�6��c�YIl���i¢������e�%ZѪd�.��"���l�`��j*.�D��E!B�ާB��2*�@�&���o�x!�KT^f�=M ��A5�vTi��Ȥ,��cY����8����lϭjSq4�D�g���w[9�&`��e�3R�)%j���q6|5���~1 �#��z~Z�.ī=8w�!\\X��p{kmi�r�����R��-,,HM9�N���?��m�yo�9��p�G^p�=�`?��굫��7 GH��{�=0��`�Q��ZH͉�B%�:~�c��m ��g�*F��Q�Xi����|qP�Ws���s�}�h�����d��u�'
�bN�������A��Y��R��ln��.JcC��=��#��Ia�/���鳶27/z��Vf�Ma�W�*֙_�����
��I�7E_oy��k,"����!;q�Ӯ^���޴���T�YY�y�~�8>��0c���g��E�Ԃm���-�-'����a�|麞 1Y����IF-��7leuU9���
j��ܰ���H�dw���A�#v���SY4C��� ��9`K[E۠�a�͚�Q��.��w �Z8����BE��㓣X�lR8FdN�Ev��������7�HR�M̑�7&%�E�����A|�$�Y��)��뵵�5[�Zf����s�b1�M���Y �
�8)^攱lh:�FK(����X9���;~x�V7D�C`����[n�k׮O ���0�`���{����	�$�6��,�>w�r "���A"ڰ<r�x��,.�����V��8׺���ZD`P�ͪ�- ��<�j<[8QN��d�}�Afz4�θH�P��=���1��$ۭ�(G#�;?��j����ʭ�J"虾��x������e.FϨ�NI�d[<!�J� �}��5L{*�]�l�flpl��{�$dX�i���X��K�9�{ ͷ�� �׊�����`�4h�
6���_��W!ērT��D$< r�ۀ�)���\,����k�i[V��ba�u`�	�6���qy
F�4-C�!�o��~�؇?b��rgY^4�t&+J�嫓v�-�DC��Wex�I�ݷ#�tuwZ76y�L"��PP8A�$	�@>����r���@t�-�qc��f�C�$��R͞�}^V��pi��Vr���2AY�7��!<i��l�;S�p��jV~D�&�LLjv*�}BDc�P��"�~O^����NP���FY�
�J#�zu[��e��`-)Z�[!�f��6��֦�)#9�8	�5�LGe	�%)t�^B�����'����o����Sv�f�W7l��[���<��sz); ~�m�ه>�~&MwK��RG]C��ԓD�@�_��}k �y������m����4��.LJrUO����*p/�?�R�@M��D��N><+ä�_J�A�a�&��Xe�oι�um/�@�����J� I��G�weX`�:����#� 7��=�"��a vZm��Ie!H���֒�a��TváC�c*}u�%���J��d�s���qI�!z���q��U����A ��v쥔���_Eͳ��d�8~X
���K��/��$�T���]�����<=E1x�X������HS���@kYb���17<P���汮�_66�X'�z�Qs���A��O�4�
	-Kj�	;fҭ�Q0;�a�P�i��J-�MN"Z��:g� "8'K[ 8�ޅ7���f�m��6E���ikd����� ��ڳm�i��V�� �uut�T�^]��a�X{�:SK+��œ�;��j�:'�݉TF*�o�:e?��O�#� �bV]����Wdu��8e��}�S��N��+Wq[�v���S5;�o�%XH���pR�����ʪ� h��m��޲��%�|L��"G�Ԧ�Zf��;57T+Vd��.ń4�tv7xe�B����yS�S�n��IM�'��G�02�׆�Ա�|ײ0=c�u�� �evx�:�F.z����j�h�~��R���s��DR����G�w7�A��?��=����6�;�/~�#H�b7���Ӭ���_��E�@��W_�?��M\�j��G'�R�����o�Z+���쬕p��f�ljz\�&�d�J�N(�*Z&�ё�>���i�N&���-�;�ۍ�)�o�t�K��u��m|.�/2N1�Y4=�9J��w�z���u���r�҃�hS$v�jx��e�8I��}��cI�q v�8�h\?h#C8SۤnY.���/o�\"�n�ڳ��T�
��֋8X�|��ʳ�B�R��
�T"���=ԡ\ ڱW_I�~�#�/|�),��D&ְ���͟���uň��>��G5R���l||YB�,�R�vm~ή\�����į��z��Y�p�m;|p/���[;{T��<�@>�Wi{[����3���TZl�b����͂�m�-�m��j���;l �u���V: R��ِ�B/�:v��3QA3��^��:i�>L���X0��Ǣ*ȴ%�o���w!�qn�����<r���ɼ� �#�-�5`��3[���KF��3黚��YcN�0�wJ�,EƱ����?��?�N�������}�Qy��e�����mjnڲ�YQ��W���7m����əU���%�擐Y���*syP4�r+挤��s`��O�\Si�Mv�8��BU�Z���<|Bqj�M����x(i?y�5�ſ���wx]X��c��}� �|�t*���6d;�9/v�����'�ܹNF�3�� k\dq��W	&5�|@b��r���Y�>Y���<�o�������0&����98j�XT�*��O�4ț�f%�pB���� F�G_y�5�H%�����^�cC�U��9ƫIۣ��H��+x�׬����;,ۅ��!v���"�a���M�]�#��m-��x��n���Ws(�� ��;�W�'�b��� �\���y��^<�ޞ�M�9j>�2io�S�I�<��>[77���/%����c[����B�U��f�5[�9���g�� Zq^�\{� F޿�1�-�Jd9K9>Gv*�#:{��y"bq�y�SD�wt[��wA�nkQH�8������t��98���A����6,�o���tSw�:o1� �*��L�m��$))+��I��o���� �[ե�����e$��Ф��9�9�*�*�d9?�
q��/�OWX�kJtbu��_S�U��h�7�<���s�=�d�� >}?���cqʻWk���p���_Z�ZZ�\>x!�&y(q'�Z:��'L�DH���HX��z�Q5d���k����p����]�J"�q�_Vſ)/���}�`R^|y�h+k˚%��@�ER拓��A��A2�	�ߛ�_���f�Ա�;�M�i�`�m���n9r!�`�͜d�'&nH��=w����:a�/�� � �|׭���SO��E�\�t2�9��������g ,f�r �y<#V�7�� �p�x�������K��F����3m��̾�����2��V� ��.LB��C�$� H��F�@�Z_��WbЩ�!��w��	i3@Kb��U	��	�/$1E�<�H!��H��T>� �X_�lZ֓�s:xҒ�Ú�
 \��q�gz�����"Y9���Y&Q��@s`>���}w�n�Ɉ�Y6V7����5;p��q��7 <��[V*�;O�-GG5�:5�h��uA����_�
��+x;�"ӓ�6<�*j�sZI���n!��?�Y�W�>;=5�dk�"�R� �h����,0H�e�������p�ܻB�q�)*�%��8@Ef�&�����-�n�		i��ֲ���ƄV*��T�U�h�O~:M�շ Rh���vwX��&="�۲ h��:��a$~H��VD8�9"�TQ�k:p��b{*��%�:<���{o��������������/��_��������<��8���<z	َ�<yN3i���5�E�>��gT�GEg��^�ى9<;�W���6������c����@ZVǐE+��U�[;�L�Sh���cw��N�S*�� �p11��X����8$�t��waW�`g��VV)B�G�R��E4qV<�)�J�$Ź�PI+��H,hBQ��>1�E=�A<��5Gl�yIkY0�9�(��sd��LU���&x�`�����ި����z�߉��v��!��S��VS��C{NXn���������H1�"L�pږ����%{�Q�_�Ʌi�2=m�>�s�Y�@ �1 �8�-�����l�n��$Q�rcA�9�x�N�q��\�Yc7(����u8ü���U�BV�r6���Y�6<���=��G?no�>�R�t/�p8`m]�6t���=p 9QTj�u���G��m����.3�ف��q]�<�:�[�L�v�ѧ�R�y�D�����xV�k�j��S��$G> ��И�=h��+a�WZ	����H��m1�[��XP��>��<0�ϻn�'_�{o?b�w�%��h��������{�c��`w�V��=t���n[�߲���9�~mں�{5wہd�"!��=��¹t�����,��fY3��D�RYD­��J� ��h�H��-��"��VhK�v�8���:��O��r��}�,�H���Y��C��*ۃX鬅�RU�ڦ�Bç'�gU8@�ar��R�(�f�ߍ�TP<�J���Պ�,v��RZ�5z7W9r�l��*�;�ʴez��g`�qV�Nu%�~׻$�]A�7���⭳�q]M��aY[��Hu���ξu�z:���~ĮMްKW�ٍ�)�%ۿ�}�#��5���_��!c���M���ݎ%A���p�6V�P���������%��2�$�%Z�K._R'(�NK͖{.��ٔ(����tG���2۱&�Ʉ�09��b+����ؑ��eg�¢��d�Up�G��c�_�-�p%`�4�25��-���bl��k�c�ņL��;|\'��x/*�Ar>8�Xl.]m8򖧠�!���Z�����ޏk{vn@����ߟU!�����ӕ�с;�֣�5FBn�[��XP,ż�� �y��d�Y�,0�qMS���� ����%Q�i��Q���la��K��R�h=|;���v���6�܅���'���\^���N�ȅ3W,־���LuX�j8}1-�C�k ���L�yٲk����Vg� ]�
'�(�(qj\וs<�%�Ȕ1�D�ǧM	G�E��Ik6�\��{ku �
 �s6m%���/}�%c��lu
w�I�"����(��4N��x����S��FHQ���5�;`��H��Ny[���x6`/���}�#���������_{[`�S������?��5�1�ۮ���g	e���(QXX��Q� bH�����hP�B�x�C-j�BwO����,\�[�F���÷ܪ�� @E3U%����pE��_��r]�t��i:M�u�+����J�Pk4v����d��V5	8��K�;EV&N��h4����9cR��\w�F�Y �p�K��&[֤)�����[�N�ٯ{�@�3����n���=x����	Hf &~�Â@�O>��ip��oōE��ﶏ~�}��%�ϽHp��������TRUJb⠔��2�8@B����d�/_���Y���F"4��f�ǏX�RĜk@�c�j^�8oҶ:�%�e�Ç�axl���o�<k$��o�IK��� ;4��:[���`ԝ�-;�J�E���9P�\���F�CQu*�l���̥T�Z� I�T�+��{*p�ڑ1AmkX�)�ݍ(�@!�"ꂛ1���b��~���c��O|��^�RP��Z3�i3sa��g��9x�H/��"_�G~IP�6WV
@2��_���� )��@�cj~�F��SG�~tLzVV�TU�"���ݣjeL�uXp�ګ{E�aOg���8sG�E3�����i|��v��U$��"5�	�w�Y���*������@6�#YQ�9�LV��|J�UR)�A�Au��p@p��� d�!RBB� t1��RX�͢��A��������n�4�A�:�D�#A�g�[dr� ������l��9����=4���a��,�w���!{��Q���"р�{b�}��?�M������p���� p#��_�n�}�~���g�4h�J�u0�� ��}��'<�����,�C���Q{���L�k����2R����*���F�h�t�����G�te�ŗ_�� ���%���9d{�q���F���P���q
T�2�J<�Z��$�o81�7vmH�֊��y��'��'_s�m��L��"�����֠�Ut��X�����Yg�7�eӼH\ �<�,w* 3I�9 �أ ���?�xȿ�7��~��N�m�������%���}�Ɇ�ĉV\�ۥSo(.�?��]<�&��v�f����Nɤe���9ľ���87p���z��^�}{F��
۶�^V"ę�0�ac�S�����#H4�\P�c������U���*E]���<���?<f��ߎ�������^�^B�l��2hH�pAÍuPn�ϓJ����b��s������f�ˢ�S9Q1���;��MN�*���@�G����c���>���i����y�k�4��P�l�n��8Ϊ0�evz�^{�9+ .>x�m֓M���a3Н���u����fW���^������w_�������,{=���O�.EYX��vX'�*��8�	|A�r\�>i}�[�i[�6u�Ζ�HS�M��8��q�߆DU�x�Iu�)��`Y�RI�Q)�D	|�k���R��  ;�K�(��T�P���l��b�C���X�Q��:�%�F��:-��^�k�R^5�^�8��~�����fԱ���8s��M�L���L#����9˫������G�~;s札n,��X�8�ߎ|¾����V퓟����W��ve|ƒ����弮��I*Hǘ�~���y�F�����蒕	g��V7��k�Rs��ꘛ�S�NA���"Ф��k�O���}�.^�a�<�U:�9� ���¬��� U��0�=�!A ���/�s]��y��57�&��3��&�A���8�C�p�޼� :�R9���s�5��6���� .8n=ȍB ��Wl�R|N��5�T��\���:dĒ�m�wu$�0 ���Tl�v��ML^�_���β���Ƥ�seq���w�{����l����۰�2�z8"���;5~��Wmnq����F�W�$(dѓ��n6dR�,�X��.9>����bGϜ=�k�b��1��������<j�V�"wV.�T8}pqs�u�����xC}�;�q�gW����&@���,��A#{�+�H��ﺸ�bV���ۍ|:��yP���H(2�=�3�5���l�5o�C��	����;|V����d׀н��yAo����-�����W�Zors�u`W�����Ï]�L*f/>�@�����k��{dr}`��^{��v�`��AK�3֙I��{m	R�UUrۑd'��������������Cp�N$���mUu�3��?8��M�ި��>�|N�R\�HpWVWd�ܞIkyp��y�]ؔ����8X]���hC�o-�`�(��D�n�E�|�Bս[V��<Zn((� h�c~9�*����AAs �U��~���ƺRK���dXٖ�([%�a%��g��S]�o'��y�Z��eh�=]���f_�O_���!��'��<� 6w�e�����5��ОakOE��+mW޶_<���/��/���a�t����~��#O X��,��J��vNB������6�_<T�Ed璉>O�:�%���L�yذ�R��6�D�>��OX#��o}�{� 5���1 ��RR�g9ghd*�֎�nxӇ{Ca&��M���f�[�	�j+���$�͝��~��	�fo.s�l˶7 �}�3���MZ�~[w6>�RM�҈��TJz���Ŝ׎*U���nj����l%������ey��v
Apt c_�ʷ��_���X<�)���f�_}�6�n���_����=��Iѳ�A'=2�D���k�����6���/�	�\���=c680����@.+��b%���:5qC�.;z�B�J�:�hrO�|v-�C���e �i��0��Cidh����j$�C,��KץPϣ�s��t&��Um8�0�[M�:��Z���EaPa����*�����sH��
�b�P5���S7�/�'	$�Z+�T�=3s^+V�|@��D7�zc־����ؖ������6��=�rv�����]�p�6� �G�w~��v��}J�z�֕hZ��$��b.�$�g�p�RH�(�N ńh1�>kk+v��A���Gf����n�}�3��\(t�ѕ��c�Yu7|ָ����dݑų�
]����1����H~#���~,T��=�;�-	 �2�%�tB`|��g��Ws�~q�S��>���%v��7�QI�����Til�*��o-я�y�5p_6ʔlH�;��E���~gj��c��&�(�b���E��v��C�g�����/�CݍDg�:��?����&�O���e?��,
���HV#>�睴O}�}��ߺ���?�'�6�&���ގd�bK��R���z*U�-�L�܍Y)�Qle�ڸ�@F�i+�7 J�`H�#�n�*}��K[6�幆�Ɉ��U��Wmc�(��(�9���83y�|2)�ì�m��k��f�
�������uG��^�V�^�k�Ǧ��<�(�!���k4\�~b�#έ,�?��64b= �>\C9U�Y��,X�<)u&h��c���3��g�>!il�r�P�s��Cx�����G?�O���[���._�o����ZWW�&'����~�}�{�(�mo���9k�a�'���[�������ܼ�Xٟ��a�O���ѕkW����F�O棡���U�K�c 4�O
���g/�����}K�ze ,.�<��[$ݭ��z���YϠρզ
%A%�N����ħ6��1�W�v�X�i:x�W�
�*j8֐JM7C�p0�n={�Zvp��#Q�=ꡖB�_�N	������/�Fgx^9�5�d{kb^U�yۻm�'k���C1;~��8�����l�R�O?�Y��{��3�����?��^����HỴ���)V��G?/��6>?/�ؽ���!�G�xv��U7:��FY�oJ�~reA�U�D����_��|�snt�N�0_b��͐Gij�v�ټ^�V�5�Ws��8�\^�tE�@ı�T��}ǝ@i��T;��=�\^�{+��E��GǬcd����p O�n��ϗ�Ll���3�qT��l�0u"R����벧#+m��|Q��de��nZ:�������sȒ�u�4mm����!������N0�$�H�A5�p��;kDĤ+��0;m]ٰ�� �,��Ū���6��*��(tE�y�)S�3���>��ƞ�L�c��m!	M��,�͘���y���ͳ�7���KMc9"!˞��y�Όgz�����JԩԳȉ��8쐳�CZiU�]D]�d�Q5���\`#��"��y�|Pw�v�oҸ}�����7�y��w�:yMM��WEp�1l���@n��.���6��4�x��]��<��yn�[Y�`eK�q=��9�LjΝ~�^~�Y���'?�M�nޖuuvJ��¹� xU+����608d�7�y)/�*�T�"=��$������|������M�KC�Z���_�3z�2��eӖC�[]\���>���҆� ��`�]���8�@`[�)*���
� �����E�U�������r �|�|>��(uH����x]!�	�H�L3U�\ߴm�Td�bF2��э��i>�
�~G�Ӷo���7��sG�c4�''��U�����z���L٣=��Nz&�\�f�0���[o�J��[� ��m��0W� qʚ�p���*�����������vcjJ�z�3����u�$:��P���
vCs����ЃG�H����gӐx�\P��i-�-�i$�A0+�z����>g�Θ���� �>h4��7(JbE��{��k�<}iȾ�nk� n9��HX(�D��7%�Cz�`��U��bA� �����
�8
	��m�m���ꚍO\�B���Wl��Q���?`i$�o�����I^�ϝ�$�O}�7llt�~���6??k��C�y��6 V�wH��!X�.5$��k���-�6�&]K�E�!�
���.�ҡX�����q+�s�gߘ��H�m�kvq�^낭����g�Z��V�6q-��;���,��V����֟�^���^B���FMs������΢Uӣɻ�]�UC$k�+� d�I��0�N*�vs�;�N���ѿ�Dߚ��� Mk1�$�\X���
�gȆ�z : ��w��������~�w~����S��1{��7��~���_�62�o�sڃ��c{����/���T<��2�R�Aެ��]�r	�p��]�q�:{�l?������v�^R{9k��Te���vв�� ;3���������<�M!�����XxVSׯ� ̗���J`��t�(���л��b��]�d��E��}-�	;�;J�����q��t8���S��>cqH3���c���z�c`ȚєX ;N�г �lU�%FMonP̈��H�4/n��b}4d�j�zz�4?��?�3;������7lv���m�����g�����~���@��?���wX��K<����+n�^��ރ����C��li~Ѻ��cG�<����}ppP �1���1���|4�`vvV�y{�u����?�3�>1�k,��D⸹�`jB��N�J��cU���g������Q����o%M�|����>�V��(��Ê�oE�1Y�����32"�ǆ��o&5nv��}�n2�4�j[]]v ��bQ�
vp��k�G\���~�� uѾ�g߲������7�Jۿf{F�����ؗ��Gv��c�������{�4Vk9���S������Ç��s�|I>{,������J�?��s��-t�u���L�#��JH���uK����gmfvJ��kˊ�u�25$����j~�>�Ob��������d�Ν�d1�n�G���ků�������#Q�I��2Ö�2��l�������+YMG�g��+���s"(����]��kL�ч������,Dl�P���e���=��#6vlL���ղ�oT����ҥ;}v�c�"�NW�u���DQ��>����|6�xޙJ���G��&h�5Nq����b��Q����9A�+W��uF��c�Z_:kWnL	�D�lJ(��@�h\T��A��7�����փ_��ka{��:;��㈡Mu%t���wB��C,��s�gų)��X��ãV �i�:_M/��O�Vu)sMg�9$�?Z!�Қ�fc��G�R���8�=��v�}��*�s,l�[5�� !g�����zPE�s����im��^3���Ƴ����3������635c��[���e��ld�! Ա�B�P�	0�P���'Z1��i�t}z���+v��QKuv#wA���a=�:l�q ?�38��~�}n�����e?��r�bYk�Ëm�&i6Z����(�`V���Q�s��)�r�-�E��L[����9E�[������^��ܥ�\�w%�Zͦ+���%���:���~�o������֎���;:��/=^�����wz�#�������!�G��ʶ�q����ig�\	`b�^{��]�:ax�	{�㟴�܆���9��K/a�MZ�S}��#�e;�D��k��cUv�����U�8 
�+�Ե �%��nER6pA	$���U��;��:/�֛%�" +W�[��~��6?�Κ�a��3�VB�n�O #,siuH�hU�<���{�q�%�a�m�VǕ]A��� �.`xB%W5�1�"E � E��d�'� ��[һ�Ս�Du	�Rq�����i� $�v*�f�4H�n?�����'?h���>��p�1n�x�E$�WԺ�3��}۳�x�Ν;o�d���8_��*�l&����%��YXB�����yjr^0���`N�������S*��qEs)~Ql�{�y{�{ߑ�k
�5�@�g�_]���m�my���Q��Pk�V�~���������+:L}�y��S��Y6FUR�EG�dBN�����❔��E@�j8�WM��W\K1�"nZ���E$�R����8Z'*�/y8��\�u�m�\����v��^{��O x�����%ĒI�p2pl#�OH���L ʅ��rG���g�lvle�`e<��Ҷm��	X��e� �T�6��e�B����~ї�m�~|�(�c��])���m�Ƭ}���C[Y��el��M������}�U�Z�N8Mw+����-����J��oz�$���<`��)�SGeB�Ay�u9�I[IHG���5�dy۪�.}��oMgY�x��O��$�����L���а�����Sg���?���v{�����x�]Z����i�G_��چ}򓟰ξv�]޴M΄ L�Y\�4DI��S
�ò�1 �E�{��#�ÿ�1���o�$-A��xR��7����������k�����msH ���3�ۤz.N߰6�v�V���Yܮ\�w�s�w��zS��Z'�nFK~��o�8h�<a�b�쾆��x����)�u����E;{�kh�ڑ���Q�ĉ���/Y�8�u��6���v&А��õR��U���۴ޮ���A���V7�7>���9r��ſ���=6j��C�-����u�;,��.��^$6پ�a�-�� ;��m��VD�s�R-���q+n��}Y��nKQk�G;��eK���fT��Bhiq�o�"m��{Q����SV,�5��17�D�gqO0+ږ�EG�X�u5hE�AM��s��G�v3e���;� ����`��.�m�@*�����ָ��}{mh�~��h�Z�t�/It��^��	 i������A���ż�)�>��>���؞�.K'bxv%�����b�N��=����m$��Ё}��}�z���+�ˢ���C�\�f+k�d����N��uv��f�nL�J���{n�> ����M����J�ٱ|�0QVq��%�az�Ulay�BՆ���w����H&�o�Z��b������z]Vo��vʵ�\^�(������_�V]�]_^n�i��CaQŹ~3��mK���ɟ�Y�81�kB��g�$J|^ǲ��� d�y���������U��+�����X2C��?�MSCb5b�y�T��N��*�"��% R�;��;6���Vlf↭-$�����:Cqv��=�H����N�d�. ��H��ޜ]ž���4�b1m����ڹ����(�:�Vc�v��Lg�7ҖF�k�se��j�b���Y`u�m�yݪI;bvDb�3Hfg�	�Ԥ	���� �_��~��â8����M������$A�.�W����w9$m[H��g�u�L�H�D�)����4���$��$b�w��,?���,lb|B죋�gp޸�����nK>�B����4�a.2<�!5�W��4��@|Ȧ�lgnYœ���օ}��b;�%檑�Fn�f &���<}}j�ַZ��<UP�2�����70dCe�I�>�#�P�S
����y����kpꪭ�&���kx�����=�f�[KR��KY�]ϚW�$�(���vw��������(vS�E��f;�4�~^?�o}�'��eG�{��7[j�޼����C��3�j���Q�*|�����
'M�xU5����LsI��K�Vp��nA8ʡY$�3K����H~s��G�x  �����,�^܎6E�*�UW�U��D��D6�M�~ ��n,�mW�=.tv������I?�W!���){����:l�s�nݚ_�������D6E��D�%��%Q�d�lYH`	[�� ?��$�	`F۰ ["$ђHJ��dw���f���s�sݺ�pN�Z��ν�IJN��Wu�s��}{���k�J�`mM������ѝG�/}��KI���ζ:U��j̛k���,s����s|���H���ܽ:��&�Ǧ�f���8�U�+�N��,�X�� ML!��='>�aP�Ns~ဟ2��\cW
~:�sgN�+)h��0}�o+m�O���~�SrK��g�� ��~^>�ߐ?���IU�5���Q�2�Ȍ�!�_�Be�(�B���H��` ����X�����}�h ��Wp.���?ɽ�w�p��!婊�x�]y�[ߖ� ��12k�jj�|ԕT�ɪ�� �,>�=2�-�ч_?�-��J\0�3ՁZG�`5�5g>��`�� L��:��̂�Q��Ì��g�| �7���hV�̓�TZts��R����A��ҹs2�A���/��Z����ȅ��￰��h��{����?����*5Y��s{{[
ټ,��
�c
zn��_(Cy+�W�zUZ;�ܥsR�I�4zx�/��t��}�3��#R,�K%�@�v�ƽ;T�|��q�3�oȢ�����w6�g{���{{[6��s��_4N�N�k�����{�� 䏑)��7��ٚ���x����uD3�K��a�f��#pp�X��m$>�;�!) ���{@��~�C2���8�
�����Tk}����߿*�ħ��?�·����Ȣ��~�*�6������`�(��e�pVl����DK85侞����>9u��_Rz?g������eϣN�=D�g��{���_�E�E>��?)��� M=����kR(�x3��6V"t�P�]k���e'	(BK��F����[�-`JQ<�Ѹ��q�
*���g$U����i�^<�gkI"������1�D0-z�2�{�ND��(0�=:�'?,����R�bi~F������'����`����S����	{����;���T rL�_|�	��R��S��AWO�h a.�ā�r��mܒ�SKr��)����렁Ѕ3Rяa'�V-P�nF�2Ũ\�f����u��,.��3s�o7$�~	�}`�xj��<���<U�  �� L~�v�����$�Ď9avϷ�x6D cƄU
G2�G�D	:��A'��P��K�͏��5�ێ�l�Q�����y�ڀ&���$zm� ��I�l��u�|�c��^��ҷސ���?��x�ʳ���3��ߒo}�5�IVVVd����#�)��w�����E&-�ѡl���5��~���˓�����ɝ�ems�����e���E��djz�=�9��h\@�!c�����Sz�w䥗_Q�y(���HN�Z�:�C�ǎ�SU}�|%�����΀�����X�����p����*�_��3Z���O��ϲ��O �
��^{k1�1q�hgb"\~�Į���N!t}���	��.Ĳ��׾���~@?m���
h�|�c3}�x�(W��H�)����^��(�t�x��g��bsRʕe�X���|����)T�Sr��m'���S����c?���L���i���#����u��\�~�����}��)��T|Sv�s3r��So*�}e;
���Ue�MOƹ��3Ĥf�lc�Ԣ�O{v-f����C����B���᳡b�{��ݷ�>^��%��6O���ځ�?|$#}/0�Bgo#�#�% ޗ�~s,{�~hr �A���k����O[�	��P��{���PF�NTZ��M��_�^�z>��C�cݑ�w�S�aNm���xK޸����O]~R�j��p�Q�-G�M^���{7�R�q��L�[w�m4G9CU�t���[��ę�y�5����ؓ�>���!d��>X0*�d��V� :�&�1�`[�r5N��c�M�c�쒓�����\ ����L4�`�j��&��y��+��ޫI�NAʃAC��xr�9�/#�d�$���K�"&;Q:WP @�p�@u��J>����5y��+r�ަ|��T����G\��ơ�9ulg�>�U��$��*_��/�A��S�`!�@���5���mV0�]��ƥN)?_}a��:���
$���ل�F
����P���;R�ܑ���	4��v;z#P�cNj�$�({�j������`8��'�?�BG�?��_��A��I�v��IQ�Umn�4�Ĥ*�#;�v� p��3�2)+�GT��2#��8\x�)��'������ߖ����?�ay��̮f�9}\[ַw��g��O��R(�����ln6�tS
*��Dź ���;3sK���o�Qm�R���Ԝ:Ģ�^�K�&Աz]
[,���ta�	���C���ߑw߽.���_�K
ޑ-�녅H��f���	*\�p�t&��gk��	� ���c��z�<G�@X��kI����!]'�G�ӳ25�@  E�����kV#�Le�%,#3�,��P%N�����FO?[Q~��I�/W�>)/}�U�
�����?'�s^��F*͇?�Sr��~Unݼ�FqN���7es�P0����z gz�
R��8���X^|�I���/��Ҽ=e�wA$��L�@:�����]��Y�_��b%/G��ܾ{M6��T�J����JV:�=f�%���:/��襹gɤ�M��Ib�����WВ����*�n}��;ΰm���:b�V�/Hun��;z������9�h�ʒa!A<�������E6����ʏ���?���r{u]>��_�8W�_��ߐ�fῒ�^ �
���/_��Ԓ�ϝ!����}�"<U/K�h���\>�9�\ ���776x-Ν�e�,8Oy��������j6�t����_3
:+�
�H�# ^:yV����e�MW��>>�����6�'CRB5�Ȇ&�%�bdA"�C0�4� �i��&�>�(r�1��f�2�Z���2�|BN?yEr�i���!M�s͌�y�ƪ6d"(����il=��4Cljv���ɅS��q�|���K�Ȯ���'~�y�W����|E��&ǫ�r|0��������"{q_zC}�>fo�Hn���̥��)���[���\~J^���dgԑ4����}VܽE�˟j���*���ڥ@Xy�	� ��vKvv�I�GO�w^y
 �}p$'O(H�3�����o���49 {q}�Ld�_� ^B��]��h�#�Ӓ̴wmc�(n 4{�R6$���&����/�߽!����M��Q4˱%2��H7��A���A)�q��t�d������pEff�|��ߕ��u
���m�
1�G����Ύܽ�@��{�".�
������1�>�\Zm]��@�P���t�����<s�J��}S�ݼ)��3�̕'��:��"8\��H}�F㑬��ɻ7��׾�uάͦʺ�]
�'�H%q(��d��%��y�֗5l�h��f ���c6�%�V������&2�,�Um'Y^�	�J���q��7�n̮R�S���m�0�G� 9fB�(�V)L�r��BM�=2�0���XE�����I�p�`�ƀ�{@��g���Nӏ�9𙐀��Β޿��P�}�U�R_2_J�_{K^z�`��uF�u�\b(�L���8>�nCW�"�}�grcc��}�]��3qC��!��Y#��F!	P�xUwT�1�&�\g���Jzݑ��L�T�G���� Jc,S��!O?�-�i��2
��z�8rD���}ĽaL�gE�&��)℄������hs�`C�E��'�mN�T�-Uhˁ�6�YQ-�!�3�DKI}N�Z��UQ����Q�!f�]�	��h�rX���h�Siy�ʊ���I}����ܿsC�[��n��^E�X��^Y�������yK������"q���
��ܒj�*��Y��X����`�a����
�/�a���Q�}�_�m��/��'�,��
-UL�6�\58v��t�=��׃b�bw-c H�H|>#cI3V6��ȯ����#����@���	(��j�Q�� +O�l&4�ҠGjH��N���W��A���?�s���]��_|[��]���O�ŧ��\I���G�·_Q�V����!Bnc�@��=�O��� ������B]���.�fO,q�jO7=U�(������.��3����7_�@�HV��y���������ecs]��<��a����h0]�;Ių�Ȍc42:V�����8����Ll�� ��)[k�.r�mdq2�g!}�+���H��ƌ��~��|��=��%��l"�����R-?!��J)����}�Ʒ^W;-W�}^>�3��@�X�����[��=�`q�Tٕ3WdqyE��>���%�0�9a8 P���J���[�d�᪜�uJk��,Ͼ�4!���A�P��V@s��Z��!˕j��F���-�<ͪ!��Gj�AK���byV�z�J�P�9 �{�H�{�C�Q���.�G�{��c'��V��NY�*��U.c�c�ƹL}uV]�Eן�꼣�#�pc*2��� �Drr������}Y�.��}�ߓ��]��ڒ������<''N�7^��|�{�k@z���2����t��|��w��A����4���΁��:�L��vP��}�x�[[��'�-��~���R��6;+si��A�����4ff$PW��ũy����_��l���姟��z�"B��"�\��gXu�<�rc��
$Y�1��B��K�.�g,Tm���L���}J�p⺩�k+��@���B$�IuP��8���l�$���!��+����t~��~�;os�Z]7o_�-��ҙ��?�7r�(Yy�����:����LM���|��/�]�3��v0��X){O�-�����-W�y[Ś���礮k���&m=G3j�5̏H߇M�_�'XBvʍ�{��P���W�ߖm��~�9���q� �"���*v�oNM�ӨG�wj�����D�\�5v�{���oR9 �>>$�F��ޅ� F��_�B�VP[>��l��b�4�	.$@vHɏ8k�Y�}50c}���-P���\��@n���r�7�L,�\���H��6�+_I�AS�ޔX�f��(���,�ٯ�Oɩ˗5 )��n����w��) ��T�Z����5i������|�PD�ɟ��@�p��u�`t��h㨚����2��@7;-�����\<w����?봏9v���1E_�Ȃ�	)��(��S�RQ9f"k#�N��z�����] @3�{H�����l}M�^u�rX�a����b�bk1������Ro4;�wc�w�9r�f� C�,� ���������;&Π��Q��so��A�bIʵi4��gB��M�����'˧Nʭ;��^�O<!�ۛ����zW�;z^g�K���˗����v�/�������=����g�7/����J�Z/z��g==_���ٞ�Q�	�1R�����gLB��{��� �%-��FI��'�'[L0�60�#K ��zq!�S,N��l�X^��zd*� h�]�bN�����*dC��E\Ɔ)@�!����!���k�$&Һ���{H�R�sg.P�����
2.4\�x^�זf�A�( ���ޕ�^��ё%�c�XT{X��Z��Og�_6��QDM���8�.(u^y��}����qj�J~�
\�H�2F�>�Y_,ԕ9�C���@|�1���Y�H�ӰihaAB%D7L��Q!��(�z�z
��w���qڍ#i��^I�b����ǈ<$�b}J��T�s#)�G��������~�B=��^�O�����TY׵ϳ��r>S�Q�+M}�]�S�Oh���]׸�o�͏ʕg.��/���?���ζl�R4q��)�{���Ӯ�=��f��ӗ�?�S�<?#�(,*N��LVPC��aɐ.���υ�
�{Ϗ����q����h�ş#'9A��\Ix �k+��[��%B�+ʎ��.c�6&t�A_�Ne���ge��7\b�@�%�8�0�j3=ل#��H$��x��d/F����>�{qƯ�?��9�3<�@�Ȩc<��ﳟ����Z����{k��}�oɵ�T�0ў"��_��7�11�
�PN�tz�Ԇ:(��]H�olu��`[N�^�k��ʛWoȕ�乧��b&͡�i�,���!;;������ە7�~[�t��)S
�����JF�Y�Hf*5)-�Ҡ��)��	�C8�E��S|%C\����6��>��� <`��*l�y�I~x�Q�aD'aB\*H!ռ�|M?�'Y�:�7hD���3�W��߽-�
�,����Hʝ���|�� �~�_���%Iu�����-���w-(t�.�9���wﮬ>�uW#:��*�jn߼�~����������"���P��v�&+�zo+���5Y�ؐ��_�k�b5��0���l�ȡ���g$d��yVw@7�BV���A��nal'˔]&(
�8��Ї���*�)롈����rh��h"�f��DF�B6�-�Ȅ9 �7Bpj����
5U{���ڜE�ʖ�R?}E^�@��W^%jt�Đ,9#��qG��q�s"{�~)8�Ϯ�5DT�C,�2��F�h�l˝��4��K^A,�����l<ڔ���==���Kz����J@Z_7�繩��/����'���zސ�_{Sn�]�ߠ�2"�ca�_Z��EY:�����c���L��t�(��y��'rTk|a��K0�#`��?Pp35Pːr�\h
�H��Y���C�����ݎ���wdA��ȇ^+���{�_�ȅ�A��^nܾ)��)������"�[�݀�	� ØEҪ��g=�;8�d7 ����` zOa��D���Ʀ��f���s�Γ�V�h���Z�da������偞E� [�����W�+W�_grj�6N(X�{��,B(�	��1g,���47���4qv0H%MC����|�A�
M��[�'MBқ��n$��-Yo�\;���i�M��>�zŔ��t��Κ��<�8l7g�Fi2Lή,r�
�3'1�f��K�C9�pZZ[r�ݷ$OI�)]ڳ�N*�/�ʥ����)|ҝwoJcgKA}]J������r|�';
�۲��-Aa���n����^3f��c�_�P�f�rV"�E0.�b�#�|Vjz61j��՛�u��5��c��ݢ~�׋Y�A��@��T�ܸy����d)��'���2BwN|X�DE�5b�̐B:	_�%PI溧]�,���A������E\f^��$mA�p�^��x*�~9 ��Iΐ=��`�J�{�)�,Y�\I
���q[��!�d��M��_�%W)��?�1�?sjQ~���y�f8���8�陌4��w޽s[��}��~Α�&3�N��/�������u�Oˣ��:��o��Oj�݀R%�[06��
�oI,�����ф/s��`�=���`-��|�W�tH���L��y�^Vc��2��e�u-���i{� �s�B� `�B6Q�NR�GDB�֔��3�K$�2��,V��]	�����;�ߝ�'Ο�ř�|��?#g.�H�Z�j���j �fS�z_[jw;j��޸'_����fn���)J��O~BΟ����<ƛ��c㞕�i8��זkS����w��$e�/�ҹ�%pd���^�,F`�r`��}�V��"K^�E�A�lgf�)J��T؍9٨�ٴS����z�R<�!D<�ѸikKU���>�h�JUc��Gs�)�%��YT���$�'20�[� �̑�*�K�A��\���A������t�>��}i+X��B���˂��]��ƕ�<��,��y�i)(�=,����3�Q�W�����	ɟ>+�\�qnW����J�,���l[\O[��ݻ��ߗG���f���b�������]R�CCL�8�/�y�9�Z!�Z^t��^�e\�᧽vbE���u`�&b?w50��8� ��y_i�y�Dn���J����V�ǯ)v3�Dd,6#c$���. Kٰs��2(�b����$]�*�;j�mq�#��y�n�23Z����D�N�A�60oGoF�M�vekcUFj�Z�Pm�������gŒi!��
2�zH�m�G��C�o=�40�V*�;@�q�+���Ü�+rs}_BTt�I�'e���Ҥ���Ml(��㱆B:22q67��� 7k�����p�al��7FhYK	l��@Կo��ɞA*�Ƹ�Н�2T���v ����U�u�\G.?�F '�"�R�v6)�RU3����Č�-.HQkF���}��
�����zGv�7dm󡜿x����-)��x��g4xz��>��ѷ����wPA����]���o��PP���A�+�/[4�p:Z�+�C��22�Ί�[�x\%�5�0_��Y�kN9t��!A:�2�)��ܷ�fs8g@E���Q%{>AА�AlJ(PkG�@��(ՙ23a���XA�F����$1P�g��?8:&='��R�2�,k��^D�Ċ��\AAgN��74Ȭ�=� �?}�On�?���\�Co���<���ղ������P@��}�gB`F_��*��!�_�����A����p�	������x����a�C�h��e3΢Ů�,v����� f�s�Ȧ��\U���*�C�Kh3�# I�ð 7?�dTb ��xʏ�cJ���fdv�b=~���2C:�XA�t��;�R��Ҟ�a��f�yD:d���	�_��������/,���8�S�N��|�C�Q�z��M���F�a�T�!]-q8/�F�a����~��G�̝;+���\9�!���k��G��vAwH5=Tl�bj�`L$�����	_��
)����'��$;s�n$-�H��Fܻ��������1�nlQVuC���*̀JT#�'�!��0�� ���s���̬��Mq��������.ݦ���<���H�^W���]9X�d�:����.����ߑ����4�_������1bW�� �
�o%_���YW��͗�#�^�Ef@F}��K���Y���3���C��c����Eb���rz�����̉SR�R����@2��c�;��r�wI�S�P{CG}��?\��F�� �q�󤙥I�c`����q�	�}��d>��O�`Lz���Ɠd��m�4�*c`�&��`ݤ�̪�������
���S��Db�"i�̈����T�&��ž�r)+�������1��g 9@���������_������
�Kzާ�S����?�!��)�GםϥI#E��mA��9�T���*��U��d���L@"	<��C���%��%������~�����?c)��L-z�`���!�8�ĸ��j�	L��oΓ��Llq2Q	�e����5v�Y�C�1H�pτg0�su�{�C&pY�r�сƍF��m��o=�o�eSz�[�Q*��Hj�u���έ�Y�%[�q
�F��Y����K��Ֆ�8U��[-���R���R����:�Ɔ =��u#�Q�r�ўD�d�S�����}����/��K�K�W�8rIK�fe=0��^���f� ��I�׀ �-�r6"��K�!vՎ�J�m��֫O���'d^�F*��T`�e���)*8.>���̲>�q��� �7��UAц�A�\6���oʻ��[�b����1��'>˱���Ɨ��x����)	�3`���f�#^�A��|��h�8zP@㍰�{p`Xd
"jP�q܉��-*��c�n�X��^�Ηd���<2�{�\��%��?ǒ`,���8$���I�1�J(�����2��E"">�Կ�뱡��o��k܋��<�ω����_�7qA�`d�nd��^,i���*���g����"~4SJ�wx�nҳ�N��}�o���'>�3l����z�/���c�ho_m$�r��MfQry(j,.���K�,�u�]i�  ���C��+�ٺ^KJ.?��t���#3j��n�X����'�F8�eqYWW;��QI�[<�$���(O���꣉>v���0Q����g��b�m����و�,�,�l��a�g�k8�[�Lٮ�%��@�j�dk��A� L[�d�Z��}��27W�+O]�_�/�����t�
�T�YGK�8>���z�t��oݒ�Q��5P\�t���+P�C�A�ӿ�Ψv4�(�257�F?��fԊ�w�kZ`5)����'3H�����s�GA����"�v�eLAW�\U�*Ib��F���].� S��,k5�3(!�R�b*��4�I�`FR�=�Pu�k<{"<i�^��fb6�ĪR�Z���W��4?���"GFD�邑�6����~^>�s������������'y��ט9���a�oukK�A,����շ4���X�^�!���3z�g?!5]o`��+Kq � P+�H1�N���x�~ܲ���%P�t3�����p���7p��q=��i'l�G�ф"�����V�(�3A�|@���U?RS#�{�Mڿ���S�J�B9E�s����-l�4 ~>ȱ�/ |��Y��B@��o7Y!-�1��~�buJ�a���o��_��m�G�ſ�����9�������V���e_��� ~�����/K�X��>v��Y�ǿ�[��O�4a�b�-+̂�������HAн�]9u�9�ʺ�	.b�C$%�1V��}W6��Iȡ�+!�a�!e���g )�L�*�DA�Ά�H@<�1���}��ސ�����8xx���t�.���6�t��t�t=�0�3!E���9��.ŚRCF%��u��~�Uٹy��I�8��y9��e���sz�Kr�ڻ���7u5�E]���i������#�(5�9}�/~�L�4��@v�CҶ�뵾��@F��S�nʁ���%���̧8�u�l�����gH�o�Y�h@XJ� �`�P~��/��=����HyjV�E��4����E��mtG���h���1�O���O���/���{z��*d�b����*�������-Y��Uy$����pPڒ<q�3�.�=��ؓ��Pn&��l�8�mF1:OK��占`:{�����?��g�$ِ�<$% ���`{�Z���;�����s󺯆rt(�p�I�	�ܽ���us�>���j��l���|��[���������^�����ԣ��i3��!�z�$���@�$��l>���_�F0���*�J��y����W:���&M�ɒt�Kb[2��A��id���s읳����4{�O8�["���� ��Ե�I�ېͻ7���Iu�*s�s����q���U�pW��c#�@�{nIj���VNK��#��Wp��kw8Jv~0���6��:-�V��D���Ttg��+ԥ#y�o��������>��$�Ęd��0K��,
̈���]�2ek�X��@~F(�K�Tc�����~O?W�63�~��%�As3d�o�i@M�r?1�Ԕ}1f��_�Jdl�7�\��ΥU\�F,����1�{L������1D�:�.Y��v�l�t�Ѫ2��R�s�䨎���s����CCd�Z����z�j���`��b0X4&��:��5}� q|�% ��M��Vb��\b�����e��g�Y���4_��k,�Zr�#n8��=���(a�$X���9�w%�c�Q��+��&�ȸ(�}��E�U�=6"y�_ܤ"���3s��h��S��L)��zC!V�4p����i�u*U)?��:���Ѩ�u� �}����|@~lzA�
��o��ޜ_c���]Nz�!�:u�_��wd]�d����?,���?/�N-HQ�W =@�:�T�(��R�5xE(
��`}W�m�R�Ҳ\�~/������0s�¤���X`�7�O��������H��ȥ⩡�'@���9
ס�����R;�).�vF�=
m������v2b�<1�k��	��{2�xN�@.<Y����ef��D�
< ���^6�����}y��
�m�.�'?��O��O�
g��0r�6dLQa�1�:j�Zr��:�L)�1�W]s��$�a�Ƀu&B}��sp�����hK��?:�����@�g��' ��pܡ��w��9b&7tN� ��}��h!Cܓ����@�oI�/Dg
i��0�=$34���$&��IZC����X<��>7��pȞ�5�,������u�\^�(H	��O�O.^~^�jH��-�A������/C����r��A��n�������jc�K:mPip��j�������Օ�_�&wo?�*�=!m,t 0v�����$��ߏF�*r�{��2���1_�!K�R�ҺF)�U��L��ť-+����*��!5D���)U�[p}}��X�ׁ�RJ)�$Pm��5�E����c�q�0��C=�ߢp������
��H��^�U�I��}�>�'qГ��mҢзz��%y�G�r�N�>3˫)U�����W���[M�߷�� },��83vccG�4X����k��ʴ�:h@|(nX�(���`H�T���FnV$@=R��VO��R�I7T�������U�G��O�J�QI6=������d��@�Bx�P���X��d
z����;�w��V`tmT��etφ��#0>�L�M?X�/��΃[f�ї��ʕ˲r��ҷ�ޒko}_��;�٠�T��^y�u���]�ӊ�;��v_jSSr��)��L��sR ����zx�>áߨ�v՟����_J�`_���K����ʜ����.�(?[Z��k
�gN1!��͡��Ť�ѧ}�U$t�Y������!�8��tx�q&�T{��x����+aPC��{�wm>���F��>`��M?�B>�]bHl܋���jGaR��l��g�&����Ů/'�s��v���
T�����\�ln��^��Y��&{M�
+�(B��7�	w�b�`��OUw,�MeE�o��c f��9���%L�Qb��> ('��~�~�Y����	�\\3I��}���j�T��[�o䭯$�I,����(��7�����?�t�+��e-�T���̟`z}sO��ې��#�Uu�.�3g��|VB]�nX {`0p=b��GY����O�/�x�{��y!����a}�D�/�BŴ����
���?�{Y�vp����c9Ley����
���z�P5%Tl��g�L���p�5�m�#G[��j4��T-��9s\X�F�H��u���?��Հ�����/�{Ù�z&���s �Q��=��n�LϮ`���t���8Sm����7=+%��Z>�wM��da咤U��vԎ!FBE3�1�ȪM�@A��|N�}Yz���y����Y��¶����4��l�l����O�����!%��˸��!طQ��%�l�n��.�x_��HG��:f��d� r�Ր��]�khl,��B�t�ZL8Ê �%�-b���} ����K[�~�6��PzI(!�5'A�{�/sO��YOO���0���'ѥ����y���Z��>jl'�e]x-�I_��w9����fO*�)n�G��q&]�^e� �rgg�R�U�	�_�-HO�������{T��笩������>_���Ng�������JT=9���-��S$`���~����Q��ְ�P��`2rk��@�Ud��/����X�0q��@(|�������9� J.�?q����F�q�6f�n�ݗ�^�{�L��b!�lZAz��L� �~(!��pCB�P��e�,Js_�G$/���l6Y�C#>�"����T�ј��X_{$�r��� �l�9�U�i���:
�.���` V��ߠqt�~���&�jQE�h���HC����x�٘<�@>��;�Hw�Z*( ��ơ5 �C�0�TeZ��
�<eQUGR�94Uˈg�QX���rg��S�T��*�%�I� �\�KQ_�s�!���(9�%��a`���
TYձ�=���W��lU��O/����]���i�9���[;��������P�[� >W,�������L:�{�p�Z�홲�՘��D$�X�b?\�b�̻9N��y3>O� A������0���4�>Y
4X�����[3E1��{C?��8�Ltr3S7����\3����p��"�{.�!E5Pi@o)�iPc=�_�7_���ۦt�A��[Hf�]�N�q��t���Y������JP�����}�w�r�n�z���$�(���8����y���_Q�P�
,Fj������.� :��+�Mf9"�C̬(_�	(�n���V�I��*T�^�Z�,�>��k�Y�Ia�"�hV:����mW�7e���2<Ֆ��/K�������/ѩ<�}Ž~����tSX�ڋ�G$����)������]ٹ�@��O�[Z��ܙ�r��Y2X��We��u��lH��l���c^��l������@o| ��3(�Da��cЎ�<��7�ԁ��ꔂ�E��� a C(��~,d���^��>P{�Dz�P�t�f6�3�!�"�]�^uC)���KZ��d��q�����sL&3�O�q���!Jq���äd�֋��A�vH�P����zc�� 	g��S�Ս�ng7��^%��fa��+�9��6@���? :�$-m=z�TLv5 �[���,��m��8�ʸ��� �ċ���,���ɡ�c.��b7 �$���Q�Я�zO�xy�56j�J>�N��ϽFj�%&�5��������8��7y�8p�����e�<t��Vrs����gg���r��
+��y[����`G�9�w��/�ҙ��G�)4�A�W���"�Jn�0A1��qb9�����]?�c�N�=�E����a���2���)M�2�S|M&�S����)����K{;�K�/PmK��b��������xQί�a������4FJk|E�R\G:M�>ӱ�%��
�n�,�yJz#����,�<㛏��nwd�q9�����Q!4D��6�V��U��0�Ku�����'%[��6�H�_I�HA�� ��i�*f��պȑڮ�Q����n(��{�7?�X�����}��9���~�P}q>���$�4�SF�D�L�V���T�xO؛I�x�g̢0�#v�K�]@�u�{,�#��7�-|�bX0: <W��IE����Ǖ��W�g�<L.yz���@����保��bǗu9�H�s��f�^��j	Z|�꽰5�a}��g�,�Q>�ɣ�#����8��ב�+8P�z�eq�9>>f����32�CS^\V�[�,��7�k ��L��g���䨅��>i�؉ ���>/W��(;��(��@AR�g��6?�G�A��v�1|���w�g,��	�쀘o��N���O_�����Y��%پ@�>�X6/H\X,�����;�w5�B�n�FSv߸#=t�y*�
zo���IggK���!,S�����)צ�43#s+E��
�6��xI���dP<����R�,o�S�B3�P���Ԃ4e ��)����<:�g�#�5Q���kz�ފ0��'A@k��QJ:{��o�4R�7��b:���Z�,�ܼBfuØ}[0�C��}�ԡ=���},��+
����y�4a'�0�滙LH%��X�����M%���|�.k{����9��Yȁ�g�hcW?�RC	
����ҹ�2�xZ�>1�@dC6�?�ݽM�ټ�x5$���n�i2��h�*E�-)�IB%h4�*"G:�q�-Y�ؒ�&w�3���ʻdb�!G2�P%��>��?]/I�D.p�	�!�<�M�&�H �OG���?�$P��O��ȾYY�g@�y"�ϥA*j�.�e����0�*���+R�9e��d�0�3�mU��o8Hˣ[��~@�b<���3AsnPb��Ye2D8�#�~��e���f�)LA+C�����k�A�4)V#�.2т�R(�3�L�����JD��ϙF�=�x^�kK��ӽwR��-S�liyI��@�wl��~�*;U�WZZ>#�BF�d�]~~�[��!!�g�v�v���OF¬��
*��{�y��lݻ-�����̼,_�$瞺B��G�ȝ�W�����In�l����/�)"3�������R?uR/��ܩER�w�9a��V���rU��%�6���@���A�K�O Y,D��}�]ߴ`�|�2�c�it��.tA��/*K���y2[��<��u\ϱ��_�:�%��y�#K��i�����jc�Ry��GX�����)L?~�ă�/?c/6 �C�I �(�c(fX��{HSAJ�K8R��(��/�Z	�W-e�|ʄ��|1{�ٕ��O�Zg���!|о|MӃfWp�#6Ñ�*E��P���.�\��|��*�o��ʛS
N'%���ћ���Tg�U�|�������"K��Rﱓ2�|%��9Ť��s�l\��Fd�#H^��ˬ��~,������G�����V�ק���ɳ��<F��^����ZH2��z���Q,&`S�ž�����Ƌ�r^�/��Z�eI{!@�ԴU�=�'p�>c}�zk�ƾ4@�*Y6�0�=��:nI��n��R�_�3u9�@�ԉe�67�IW�b)�1Q1k1*h�J?�5`���C�*�+	�
�њ}��w�R(��>3���"��y�]_��	�@=���~�6%e�;�#�����@�H��r]�Պ������}����T[UɆR��C���cK���xosU��u�mK��
��Ih� շ:]g��k�5��HI����;z�4�"��L�0%�|�u �jh�B˓� �x܍y���Kɱ�&���|3�p�a�D,��S�:Dr�}�1 ��#��T#QIZPG�~c������oNs.�%�S\˿F�_����?��џ_����of��]p�!�0Ni��q��;D�UCg|���s�0#�w�JVl�U,2��QN:�gq��f��wq�n�M��~���P���ޡ�2�j�ei�dB���	E���}��%=�э�AmzV�2L@��3J��/hp�BcqX��g�Z0���y�J��O�?��$�O�nSM�:� /r��1��Ɔ&y|���wC�o�f\)�j�۸����9�wpf�<0L&��,z
3��Q��``h26��b,�#:�����a��P�PE3��d6S�|%�nZ
#*�	��\?��p��g� ����%��=��:�BZ��=�Lnp�Aeb�0�� TzPs�N���CG���a�U��ňLI�ΐ p�hF�K�ؤmV�;��eeJ�a��w��uؔ��'��w��<H�3�8E9�j���T���d���u䡴�y͗u]�ق�~Q��� p���3
�n���]�~�'������L�u9r��l������-:�-��\�2�E�Dij�Q@�-���Z]Iʘ?�*�'-V,�)��df:g?H��]3p#��^��OΈ3�c(.I2��@����8�"4J<'��l��'�$��q��i��AƂ����󘋄d쇃��[����Ś�oq��`G�Y�`��?�=@�2  �IDAT2��tiƩ����>��֧芴:2
;v�lN�r�n@0ȩ��ev��. ^hHd[S_:Ͷ>~��Z ���d��ΐ� ������@�v�IogE.=}Y�,*�R[q#�!��4���dU��t�j���t�$M��
�3�N�:��H�&f�\��"y�U@s�#���h���d����rZ��r�ʞ���ץ���l\��`�Ձ�PTYߑ!� `�G�>�`pY�Ν��*'�����)���ޞ�A� ^q�A'���MAB�(JSML������G_�#����0D�TAh�)I+���6
�}0!%a�WH۳"f5��� +�*��99@��s�C�]�� ��Bu�W���`&eJ=	63F�%B�l���1��q֒��)ܽ^9ӵ5��`�^H͎0ġ�I�`�hSc�oc	x��f��N��<cZ��)��@� @����@���0�(������B����rظ��F^	�)B�1e�dl�Ǒ{<^<f��� ���D�fQ��V�qe�CS�w�ŁA�@�=OQ�ġ��XLe`���복���v���@�`�:�Q�f��֋_���ڻ�{�������ݖ���tmFj�N���		K%����h������c����b�S)�ţD ,L�*+T�R��y���LS4Ib6H��O:@�e���sl 1���B�ӎ�sϡ���؎��Pm�@�z���_�����r�&���,+g�H�q,k�Hcg߄e`k���筨�9�]�
����a�l�K�T��Ԧ�jc�
d2�1|O�Rd�
������}뙴�!�]׭Z��9(�`�(��JjKC���Ig4`B���I�`_�h�������\<}BN��S6�;�Y����O�>�.Y��P���j͆�\���hJ� 2;(�\�"O�?��3�^ő���[G����1�c�X*�^r$��)��'a�;�#H\�5�.1)�۫g�}�ݬ_�?�e��Q[�ㆆM�zo�����tl���C�;Ctփ�9R�q��E���1���ǧH%�Dl?�����?<#��q�ON2MA@it?{��A�����o���X�����L�,�!	]��5��\�s-!�
zȀ�K�.ץ;��ɑ�9U�cٿu�@Qw��� �ݍ-}lE��d�����HR�����Z�052�T���H�2MǊ�aO�����w4[J�[��yp�#�؈�oy�b�D����Ǿ<9t�������=��l��z�h0����D�s�^)ә}�������SR�QKH6�σ�5@��C�B���3��(���节���$}i��!ۼw��_Gf�XJ�)�;Q�(�-����� �fd�5� ����q�e+̤��T�ք5B0�B�*&��:�ތiP`�S09d2���,����<�"<���P�цt���o t�zb3pM� ����`(+.[C8�fg�90�V)�:���-wn?`���/���d�rt
�{����������[��Ձ��.�σV�>Y�F��Cu�P%���Tg�4ۖ�qK����d�s�s�N^P�W�I}n^����0��$���.�����,w2�� ?$e��������O���
56�3hC �����$k�m�͇�Lk��_�0�e�x�;W������<vCu&�`�%?}@S�Q�Bo�a@F|2�"U?�6O54���}̃bN$m4f�ȕ�����p6�P9���g}�{�DLn@�(v��猐��ǒ2�?����^�IKļSȑ����2 #�H��L���%��̘�}�Ů%
�p��;n��榄���$�q�	��J#��w[r�𶬪���c�j�k'���;ܕ�Q�l��ѥ�ˉ��R+� �e̡s�����`��Hr����Y�#~� o�:��5�
��Ο<I{���7���28�����gFTY}}͎� �T��"�hrr��9�Ԋr�8��;�v���;�$�s��B��	3�
&T�a�l���kMP�Ϛ(z|Q��l6T�4�(d��B��1PG����Ȥ-@L![��B�� �2NE�m6L�����F��f5��5 �"]�{�$�;�)��X��jmV�Ūޯ���¾L�a�����8Q6g`�
�N���!� !�kdR."%~Vr²�]�]��<�dx�}����dBG�:�r���!�X襶ĭ�/��WD��}ʸE.��:�ؓ��Q0�E�A�N8�c۰�(v�s�L�2��b��������=_�p4�$*0.���x�e<�6�v:V����p0��mL� k�O�!2Y1�m3���⓲������ d�-.�-[� z���on������ޤL����Y=�b�������ۈ"
yD2n3,��}����scU�m����<�\|��a���/� ��$<�9��N�����}v}�uRl�R&<��(��:jcL(�k����w�2=%�zJN������G���TE��s'�d�䲔�g$Ι�o
��7� kz/��_�����3��s�?�c��vZ]�}놼��Ǹ��.H�z{YoM�FfuՆ�k]XX�z�$�J��>)V���7ޔ��GR�U�P)�hG:ko˔^߅�ȳg���MȔ�dj�*��9i���������۲w��z�S�G향����j�1�F���IY9�('��j��1�lIbAd���T�ZCa��S�g�� ���D��I��  ����9�6�{�+-����vk��ܗ�\ZΝ�W�!��j<x���~��S p���A�%G�C]�geviYφK�����&*���K'�y�c�iŲkވ��pc��`@��* x��;:{��A�=�P�8��(���챞z��T��A)7Sdf��)����z���œT,m�m㷠�%�����˙峲��o����Po4�ɻl؟YJIy&���=P��n�!�g<�0��d��H�n�g���H&�L��l��o�{]>�gNǈQƕ?Oݰ���[�k���(�ћ� :�K�1�ݨ�n@�� ��)O��M=R@Q�@��;����C�^_�{�һ��s�4?/K')!�r>���z�0f�|F��2�h�����(c��[F}�k`� ?<��8�^�4��k�23�{�����ZUV�5Τb��Hst�]H�Cwo�zv�)Ì���B�u��
Yi7����_����ؘ��Xo����'�􆱅@�4��m�Xy�⌏�A��E�"MF�%��*�x �0�X�[pгG:��aynY��u6u�w���o�N����"KgsrbiAf԰"��B�ݤ3�d�
�����!%t�z1T 
(bA��%U����]
\RȂ׳'��T�R3�v7b����*�p=�>/8�z���xQ
�	�}���m�S�l��Cw�Fc����4��y�Y%#&-%�*r=f�ȫ��n���J��si*�Y��:>�}�V�S��gC����d�1eu��8���r���N������v�UJ�s�UH� JZ��	� &��J����|*��f�g�J����5.Pa`�Qu�<8�FY)Um�2���J����"����ߤZ/�-�#�8�'v1[��7��-�/=-)��bE�-�J!G�t����Q�ޗbE�8t�0Gp���ٻ`�ꭵ;���68>�AkGR��U����9V�A-ںS�nK�K���`�H�3+�u�*�^�hK咉��]�x��������n�H�9���Ԕ!V�ے��=K����I���1�E/ �G��g��zs:Q�еݷH@2�S��DuZ�JY�s�TX(n����v������FCm~�=�V_�Jb��fV_�B���T�}7��O �<�7� X�`/V{�eeqg�X[I͞`�UcV����9v"��;-9�� a�%����*�a�8?�(e��8M@(NQ{��>��6C֪�c8	�����)�����2�^[�dLuV0U�,eQ���{: �<����`��ϻL�5�'����``��"G���$El߁R�~H0��=G���hO��.�v��u�/t���͢���~��G�Zܷ�vlZ�������!c��X����%�C7���1��#�����]C=������̜=K&XqzF�X��b��`���8� _a|9fU1��-���E&��J(Nq#Тd������/�$�� .qn�c�(���C4���k��F`z����4;�Q���ٕ�޾�H�<��ڟ�'���
�sݻ{O����M���^Z^fUQA#�J�ʁ+00�Z��0�諾9���u)�Z<��y�ҽ��5Y��PVޗ믽&�j������MY�>�Rb�� ���RJ*Ռ��9ɨ� �e�V�����k���9��Y��+�Ş��K�LA}��P�	��RL��^~А�������ץr��9�e{G�[�WK�t�4���˝S~�͝���S�ge��HP���nds���d��C� 殍}K�����'��/�¿�j��A�X������P�ؑ�rN�N���K�y���3u�	e�]tO?������O)�7�e����|$���rU}�_�%ʯ4�Ӗ��Г7Y��x��%�A8� �Jz�Ԑ{-E�nQ'�l�z��v�ˠ����܈>�BY\yZ��kĮ,��!ѵ����ݬ�Z5ad��ѻ���)�k�*)j����X�3U)�̫K����`���w�5ߒ���VѠ��w{wWFݾ47�Yi��(���k�"�G̖0���A&^�H̤�^�t��������\&�`�wIe��	�8C��K�]��D���8��:���e*�G��i%��Ow�5�����)E>0
)�`�g �q��2Y��S�^(���d�\{$k�F��./,��,#g����BI*�1��3�Я�1�u�A�;�`R�9C�1�JeV!��쨑z������\�"�N�U0S�C��ѯ4��UAr��1PvtC�#W�d0�G�c^7ޞ���b�e~�L<o�Ȇ�G�8���w�WR��nz�xs5	b|O�"�:A�(@��"���qJ3
�1D6LG�K��F�d�,�,lm�^���#kw�P��x�sj��n�v���b!Gzd�9;�	�[��UH���}�3w�b�a}v*��=8)t7y\�9�4u���܆�}��(��+��fqU��V.pOA�ÌNf�]B%�j�=M�|ݑO9pɷz,��)lv��"��l8����@y؜�z�C��
0��"_}зF���!������A�����6�f�;233ˀo9U����sn'�=�\�}�+��83��L;�:�L���	ۋ���cD�Y�/319u�0�=�kv��6���3<Ϙ04��kg}Mr��PkK_�*��z>��ZO�8C��k{
���'���V�@.��՟����+��X��������e��k���2=3M����)��R+�emK*
/��T`�#wt#�m��������XAj��/3�h���]W��Ta^��GjPV�����{x� 0��s��hqǔ��RN�c�O��t�3F������u�m��z�.^~�4���-ΰ�ju}���O={Y����{@o\1K�0���>gK��=T�Zՠ��3�dskG6�J]���0�m�Z���*�U�s�F2�����&hi �r��]n��(BU�ԙZ�������S���^� �Rdu����Ԭ9E;&�8�]�D���ȱ�$�zB�!p���!]������i> �H���L+�X<���au��䧂�Y��b�
�+�]N�:sb@7����x	���)�d}���
O��}��A�赁�o8��W|%��`lc3j��cn�}�:�鍩C��-�cbDm������o����c>�	��%��mm�(b;��2�΁	�z�+˧e��%)�fX1G������ӽ��2V�&�.AP���^�c/r�7r6~�x����*FH�M���������q��[�aߤT�U�"&�B��@;d1@�=�jO�n����Ɩ�N��A����l�(��V����ٻ7oˮ�}�H��&c�>� �ϝW@Ve|R����jl���z�S���:D{�>��ve���|�_�wnJ,�fK�`B��>m�5g�U$����i�j\~$�TO�xc��fg�F����.�s�
�f�m4OfI��s2�^kOc��ښPr��J�e.ˇ/�}9�n���!���Î��P��80��z�S��50�zS�n�+��).�Ha������aD���Q�e�dI���V=s��u�/���2���u(R��W��?ޗ쨭1���3OȳV���S��4���Y�%�uv"��S���ʬ�����h��@"�%����eI�>��/[˟�з?����aڒM.ڄ		0	�4 14��sw͕���)"|�9�ވ�S�x@ud�{/�ƍ{�9��@>f��X[�}��[4Q�җ�����{،
)S����:=d=���T��)Wj�	k� Xpe">B 	 �}~0�TF»-��S�h����8�!��Y���Ɣ~(�e����V��?Whj�
���r�H�*��Ist��l�)�zVjr_M"�4"D�C��A�,��U v!K���J���f_��ݢ��128\�jx|r�J��)���h�B�Q��~&���,UX� �iP(�L�P��a��1iq��j.y�E�c*�z0�<upM�S�琛�pSwb9$���KkU���Grol|����ɐ҆f�B�iD�����ȅ>u�v���M�������lS�4�����i��-��Oj�p��ġKiv�.5��e�-7)�u�VA_lRC�85��I��u�Qc��GD*�"Q�u���,ӈǴ�t���.��}%qN�cdk\��z����1�Q>���Fh�|iq�V�)����Y���1̖H�VI_�x$�3%�<�IGl�٧�%n\R�&4���D���"��C@+x��C�j�{6���"����k��e!G
Rx���Ɵ9\�Q�ZU{*��I+�gNU8{�n��M��ɳ�g�{މ�'/=��@�}k�8�w���y�sh9DM���� ��1ܘbrc��hSt��!�ޒ��:P� #@u=�g0f(��!J:T-��|}����-�������H�pkk��l �%��M�x���4;7%��d�J��%j�����}��C�vu�����R�W�J�� �F�G-�w,5 ��<E�o-HJ��11��m6����E#o0�5�9��cCN�CD�x>�����iZX��b)���م�/����#z��wi4h�j�j$ͭ��"�i{�/N�۷o��������`  X������ۥ��Ǵ���T�RQ a�(�Ro��Z`��������|)b@��T��r��l8���oA ���4j�`c�ʠ��ͳ�5z��]�~�*�bŽĆW�耞����hnz�����7�Mb,U~6r�hU�r�� ւ��s���������7�<F�����O�ǯ�&�<���p�8ѹ6�*DWWV.���O
�\�� �����gRʁ,�����^�ɛ]�sy=����sj�� ��ν�wx�L�n)�<>�?���M�5��ޠw�y��ݡ��bIw�}i31U���D�������ݻw�~�s�������@�XCf�D���@�bg�h�g��c���4|Ǭ���BKӂ�^G�O����z.ER��LͰ���q���J���>��z_�`���4��Ң'�}��R ��n�(2����ݠ��yp�+�R�sr�|kd����xU��7}{ܾ������Ƞ�P����{vrB��B�z���A�l�"�ޅ�Y��~���4��9*M�oP��ZȲ!}#�W��"�}���XF���Nb3W6��f��F���H1��Eκ31P�h�,�<~�}"�8��8��<i(��n�ep��K��=!�}>l5��4K��ޤK�G��7Wש	����p^�D�oߤ��$y��1�G�J�	�y��ֈh��.�z�{#�"@��
N�í�g;h�8;��� ߀/E���#�'��#�?G�=��=��)���7��Te���R������; �gC�e"534����`@X�н�ti��s�^� �S�n8�Z�C!`������&����g=ೞD6[�G�&��#:��t��;p�����l�`���/r^���QF�O02�?�f�%Sj4���5�w������k+�������Y�|��mj�=���	������+����������A����w�i�P�\�,��bkE$��(���ٜqF�;��Fd��N�j��l��o�R�p�B���Cʢ)v�B�P�b�.�+������;�X�v��6�i�I�ڇ4y����ƈ=���[#MMAz�ZS�H�@��`��LHT�e�2Aӗ�a�+6,�A���X���+�I
�e���}p(��+?�c��sT@ߧ����Md5�n�?T(�F%y�i���=[?�5��Ix�֘���Q�q���������~֗o":��:�15&�����=�Mψx�O��u�w�i�I9�"�HE = ��#=7I�c������ �Y�\R�C��v���������/�@/�y�*�V��Ӄ���A?���B�N+;Y�O�>�sbkF]K^��r��qL�ߺB/��2=��C��kPl������W��b�5W
%L���q[$qQ�|y�I���F]�*N�$ut�g�49E�� q�ߗhd���:����k[s.��!L�#�z��F�G�b;�)��^�~ <��j`���sz:k�8���L���!E����a~��N�:��6@k�����4˟���y~��?�Do0H�)�`���<Ԙ ҎH������$0�j�Ғ���qCj3�����3M5Bj+��#�p�j5y~�k;���g��e�3�� lHT���8`����d^��o@�BURm{8�BЂq,�����?v9��V'ԭ>[�F�!%m6(${��/���J���ivv��l�mmmI΁V3R��8b`v��Ew�-+hk��eI���'%::5=K-x�Q��K{��#:�Z�H�2 �㣆�����=�ˬ��!�<��mF�`�#�`gX6<�Cj�˼�a\����F�<�o�؊�	�����$�3f��$��6�P�{���3��H#m��-��o~���+_(Jy�`��L���,����)%��M��QZs��X}�m��w��)�h���K;\�����=��b��%�<�+�4?�mc����8Q��~��˿�9ZY�c��F���M2�X��f�@H��'W�n����>�#�������^u{�
_#l�|/��ח�%�%�DRF���)`4���W��1g�Y/Ӹ:c
 9^��R:v��������r�AZ��1��!kOy䝅&Mx�f��x���T�k�ja���d����q2{�61��z3'��`QoÂ�N�r�F��E�iiU�	��@sK�3����gΣd����g�Oٙi;#9�N6�|��x�Ix�?�^�}���V��̟<�@{�"�/�i}?�P����m�3�:�Vgjt��-Z\Y�2�ͧkt��O1z��:r���Z�v�B�3}��`.x��> �Q�| �j� 5����#l���҈����M��C����daeY��YG�� ��L,��kӰ�^�McG�j#����W*�,t�t��>5�,fB�Ê�.�,RubF�7�vx� �C��p��.U��/d��t��9��1d��m��^��ￃ^����_gY���>�U�y��]ꅨ�f=9��Q�M(A��v��-�T�j�&)Y�4�zx^�&�;�v�����e7�Ę�ken�~�ӟ�O����Y�3�(���fh���}d��跾�y�M���D�>ۤ���g�������9�P�N���=uUǚK� ���%�ڱwŚ��"��>�٠�ߢB6��V�s�3��;��S/}�^|�--LK��N/�m6�?|�Io�����oГG�q�_/_����5y�X� ���6'L�c?��E^��6�HkBJ�iI��!{��!̕��}����p~~��֒0�򷏶w%�-l�P��9x���օ��O��"��n��iO	g�x�dD(zV�p��ǘ�q����9sr���3|?M���}��r�9�@�X-��>r`�eV��1  Lj�v���!�k=���H�t�;'��D9���Y`P<��o�|a�z0 {��E�A�s�l���:u��I�T2H������x�S7�>ZcE�ۑҳ���d��~�Iǻ��d�F{��PA�G�\�z�s��8���qh�|R�E��pl���霷H�utb���+��!z�hbfN����D� �w������m�5�R�猗d)`=��آ=����S�M�v7x���Z����yr5��,�N�~Ƥ��� �>K��$)eZH��'�q�IEy<%��ڥo���;o��
�8H���5@1P�q��TA����"'�0 [�����LF�����ߗ�rժȪ~�+�P����s���T�B��f4P�Xe �Z��Q��5����N��k#�?��h��C����bL;��e��:�w���*�T;�:j��@,Γ�T�ԛ������4v�\+�NB��"J �5җ��+F�6���4�ttxH������L��g�R-�$�/�@#
�)�����3m=����=e��{��$Qw#T�u|O"l�Y��a��=������#"|�o�ǈ�W>��z���P��g��5�l\1(-Պ��A\�l@��d9��@Z2�B����:P���K�5}�66�,ڡ��:QfC&+i�(� ��G�|����ݥ�{���w?�g�;T]\�� L�a��+2,�Xh����|m�}E�l'>_F��ش�	+�W�M�c-��}$��F�}+��K��,�	�ᙣ��طP0z30Xց[���(�M0=~�@�,4Gg�q�R`0�r��������$]1�"w]�W�_3��%u��-mi�uO~F�-q;7^l,
D�L����)v�ݧ���w��$6�=�\���T� o�=�TwIPqt%#�%�'���R֒g&6r�i��j���wCx���B2"�`��Q-d��pn�S���1�ʰ����]���m:>>���M�c;rm�
���e�r�����0�"�i-(�)5�r�X�K#�1�nOX�6��v�E��G��Cˎ�>�z�>@&Haʕ<�*�� ��rj(��:��4%ϊ��1J��*�c��ɱ΁C-��)�@W�x��b��8�f�Ӥ���jГ5���c�	�s$���TG�;T8b��:�s�fGT�NI�@�umv�H=�s4��V�z����"� �@�,��~L�v����=Z�9&*���T���1`�L��A�R��a~��-Z���O�9�w�A.�aq�9�G��Q pV��ox���]�_��������H%��ڼv����x�|���sK{J��L�2��,�X�bb����hw�@'^-gy��M!��\�/~��o~�t��U���M}�H���7�/w���}�w�_�+z��G���]��v��s�EB�a�=cHK��e���_��h�Z������{[���b(J���
�ˀp}��3�++l��0��'x�h
#Rc{�"���{'g�����)et�
��
^V�:zyTv��ou,*v���|߷�����/6=�T�X�/z͜�g�lDtX�/]uf�*�<��iwO�I�!�M#p/k�B7Vcd{.}�7hƣ�x}LЧ݄�)���%�l�u����Z�ږ�Rx��b��<H�q�F��}�E����`�{�]��\��e����y��T�[���L�ڔ�� mP�'���{�����{�1�ր�~���DQ%�Xh�+e��p$x�����N���k����s��8匲׷N2,3B-���4Fґ��sO{u]�ଗ��.bo�9�����Zָr@W�Qm���9S��d"�ghϥRD�a�R�IR����j�����U	��H 
�j���oMթ�ZHOGԤ���W����y_�T&+T�Z�j��n019���ZI�o���5�&f��G԰R���e�s%c����с�?Qx����n�1S���s�0
N�%���LK0�^ X�(�.� �Ck_j�G�j7�� J	��_{iaNj���I����c�\��ד�V�5v6��/u��HwA��zU>G�^��
�(C���
z�m��;��9��M룾:1�� �9_,�9��tԁD=T � �X- �#~���eD`��J��O�<�߱7��&��'H} ؛2��������?/=�<�O�d���<�X�k�P(Rmb��ݞ-q.+~��C=d�U�in?
k���1Ⱥ�o��O��5*N���O}�fn���ǂ�eQj�B��S�M�'*��H�,�=~r�tm+��@)��7Ԓ#l 8����2�|Q\���'�މ~��#6��~W�,l�.K�dZgz���D��q;���E�����ܿIywF�:�Hx\mb�}�L:�G鏋l3�$�!���M�ǳ��ll#7O�v�BYqr$6�ߑx8���lJ����9�/y�Jϐ̐=^p��1 �Ɲ�)��|���m�)�~g4��� ���Q�{tH��S��x�Az�eJE�t�-]]���M�{�؎�5%kii�
]�y�ʼ�;ҟ4�TX[� V#Z�t��ȺP�G i rH����u3���n6�	i��ԋ���2�:���AuqI�5������J�l��~TVa8K,�o:�t;"C�S�5<x�J��r�k�`+�x<�9�D�����D���`�7`C�fG�������CBF�U�gwo���K?l��HO�PRM}_���|?��	ֻuj�-����Dq_tm���>�9�p�ڣ��i�y�a�������R�<W~�˂�-=kڦlӹG~ a���4}���X��ܭ.LQ��NA8� �i��;�!�`P�=?I� ��M+$.�,;�#:f$>�6X��c�/����_�+z��������BT��/;�NMV
T���W./�������wo�ѳ��d�bԅ�F70H����E�ƌ;�!�_��ɜ#F��AHyS�2A������@3�uc�����M�͊����<�!/���&EN�1R����(
���F���ؤ�Yq�3ce��|e���Y�X�G�s�����N�s���+�Z5��>$��P�Q�]<�{8��)�1�LΈ��F%X�$� ��\�k��Z�K�h���nfɽ���[��X���G;��?��B�b�"�J�2h5LQ���<��bb*yDi㗰=��Y�#��ؠ�����K��NQk�Ӡ���"��c�2����S�r�]��23���f�Ā��F���Pi6O��4㗞��ȋ�Ec���LO�4;����3�r���m�����暞���{cx����޳�2Ғ�o��񬓽?c�ڵ�I_I�
l���=25�B���v.PǠ�Jt����>ڡ�|�{��i��jE� 
�8�3�ԏ���#��"�3P�H�ii{�00����h4Rg@F��w�� ���F5�u
k�����25C�?�n����Ov�L�#�ǀ�.(g������٨���d. N4�K��0S�ߑ�Y�U�h�~l��c��ie�*,��ӅiiA!�5��C�k`�.�����;	�/Z9��/�:͌C6�p-�@%� 0�ўz����X�I(�(7$ek( �F�k �3cyN�/��Y�?���!�655%2`smM���l�@> ET���r�j�*��c�?{���5o߹����O���<?:H-���L�	��G3ӳ2/0��̌q���	���7�ӟy����ߦ���`���ݕv4���R�*�[��fc����
���8�p�Q��|����mdZFi[��X���F�ɲ��d�{��#|4�(�'�x|�F�)o�>��s����9&:��sG
j���>����Jش|2rl��YP�AҔ>;�}K�c�e��:��.,�NG�����V>�~��$	��Mik12�ۨ=`�`��F���Y)[��J:�~@�M-_d���:�͙������/|Dۡ�����֨'S��iK������`�3�Fa{7�5ww(f�6h6���P)��s�����?�O�[;�a0���KKt��&gȲ�#R���۹U�X�a�3��;0�b̈́8�o�ڮ�
�P9��.���P Ye�Fu�X�cI�t5��:{��noH�ր��&p!ؑCH7�֏ho�1-^�L�>�<��)��)#� _��ȇ��=������=h��ߣ:�AHV��)*
�N��H��G}cs7��a�X2
�
C!��q ���z!?�e8�8'#L�=4&��®�@а�y��0t?۲u�M�]]�KsU��(�Ƥ+CF�Ƒ�ll�O���ț�����m��!�� ]�H�2W`3��:����ҥ��@n�Ƣ4���:����=�Z������_����_�
�ͅw(@�se}m�
o��H��3�"}᳟���#��ݧ����xw�*Se�yY @����0�c�(8s�KAa,;E�B�|y���X���u����8��U^�<���<�f�$m�ѯP��F:[�p�Pf�1P���VZ��ZwG!�b��5�h�Ƽ�XO�]�����^��)>��u����gL��P�/6^�|F=�H9վ��ţ4�Lo�b�NŘ\�]��5&N�3i
�4�>-@6�Է�y�o�vM��2V6��v[Ml�#���؊��0��B�n=�i �Կa�� �-�t�8��3�7����	f[���{#��	A�f3�>vi�=1X~�dJڽ$�'2���4��1?D�����Y�U*K#`)�N���xrI�wJ�5	aO*GZH� �؁A����G��X{�}w�Ax�w�=�h��H��Lld�=
��=����I�M�y�z��/��	�i��x�X�����T>V��;���,a����(<�% ^�0g��(�%���B�VVV�Y�Gt�חZ����$���M֥6o�����=V(��[.�iqqQ��;�--U��20C?Ca�˲` �(��7!��}&�3���t��uz��똖�y�[//m�&�Ӓ�	P��'�����q��u -zߗ�Q�����4+42��"��t�P)�h0�g`8??+�J�w|�>�z�s����%�/��8 $۝������� ȡqq����y�~k)�D/]�$Ú�9 �E���r�*�����9"���"��y7;3K��+r?ƻ��#B8W��$y2������L1�E�	i1��'�	���dqO�s3��Q�g/ƨ�:��HHJ��r)⠡0)+�smD�����b���Y��CvX�3��F� ���>`g���b����S}�|*&�qk6p��g0�cJ@�5��9	m��u�9g��o\�.#�v��?��O�S��8�Kq��q�p��������y�O
 �-�I���F�ŊC���i����&�6�Ṑ�Ώ��V�Kr\���I8�im>�[2)��o(v�Cog����b��)�s_���k�al�;�;��]q��7��#�<� �؎�����KEd��x�z�9�y�9YW�=���ui<?hu%ز�r��޼A���y�u��x
ٻ�+�gb���M�{��������Z�����xƗ��R�B�| �飑�l�n_d)RY�G�R
P�OIF W��@.#�u�/l���t��k�T�l>C�өCۇ���qL���=jS{�i���*yR �}�-��_�ӥ��|@��Պ%��4�>��;,�3p��MTEG�Y'J�9O��HB�#l�ѠK#O{֢͞%6�K�X�Fc�.�D.��9����5�zi��y��ҡ ��K��T����5K�����ݻK�{�] J~FZ� 9!���~�l'��Y:��۞^�v�"
�f�����&eJ�,�>���]���BI͈J�j�u�W�7����@M��XXS���/�(5���HB��ʤ�Y��4������=wҘ�g�z�n*,|��C������k7�`kM�9����ne)�1L�L���e���$�<,�-WW��؋lxLM� �@ڒ�/Y� 3�QJ�|~����)��n�1u�/JJO_��G�^ԋ��J:�K���[5�����P���I��<G
�6�6�=���ʈ�Ƥ��q��,0�?���}	��I�9c"\�26!�@%�3'���*Mz��	c���ٶX`*��9��SF��'�<g�ڨ�X2��%6�cm���ՠ/G�94;�ӆ� m��՜.��3G��ON��^�aq�3��+��������QG�3�,<)�VB"�L����@�D{:�e?�`���[�|C)��Ɯ=�M�:��E���aY���9	���Ƞ�!	|*@���H%.�3�#��O�Y�V<�A[���N�ASO��H錣,�	��6e��`�|Y@b-y�$dE�MONK
���:��?T��<�2��ٹY�z�*��X��Xi��C4F?�L>+�-@��%�ӗ��B�Ǳ�� @�,`�@8vѳ��W���$��*"{�[��K����>�⋴��,��5ޗ��H�$��Q�P�ހe8��w�AO*f�lLL��K�f���(���:�pf��=��=1��ƥ\����A����WiffN�5��:}D,��6\��iV6�Z?�� 	P
��C� �@��;q&e3ڊ��c�{9��gqiARE�t�Zȑ��AW�ewo�A�T�e�ՊRg#)X��9�y������%��C�|}(�> յg��7_�g�S�єFׇ������ù'��]V�	���g��6UϞ�!�R��*�C��}�X����u���.��9��	o8[C�f�Y�1��4������R�T��_:�/�4J���j�$Ɛ"M�ӡZy���j��|�Fi��:��:�f&q��d�V�3�Ər)�����,��`�s��b�ߩ�-��-��c3 H�Rc��)l�������$�M����
��I&Q9��q�,��9�>Ǝ��J�L����,�VF��V��/��<l��u$h��٥��u�i��e �t�*]�vK�̟=}Jۼw��v�B�3��H�nݦ
JX��j���H����ԧFf�zG@&�$鞱��#��$mT�t����98�*�@��hQ	�ϲi�]�%�;B�R�M�l^���ya��jC�������R5;���#q���BZ�YfT�t��"ͬ̈�ݕ��]��s����dhrz^�<�Y�H[�=��߼C�6�N^ޥB����C����֕i��nP�<�S�zri�!�B�`-+�Xdy�: �m\�'���,�+j�@�Ll1A��n)xR��g�� ���[�q�$�Nנ)y��%k>V�f�fn^���P����"KNhw��F�,��Q	�������9�xQ��Ѡ�ÆI�AQ�A������m���Ȇ�@�W�����z*<e�ƴ&r�*\��~�󟡿|�;�}�K��)�Ԧ���"�%$%��s&����4GB[��Z�&�Mi����U���_��k4h��J�ҵ+4�
��+��.E�&�����FZ.�A��
�j�b����?��	8L�F�:����
�01�O����#yؼ���}85{!kB�9���!gq�4��pښ>���/<Fq��f�<+5��O�mBl��fm!�!)6i�2�#��<����΍o҉�	�W�*��T�J]�x�u>�(����3R��q�8!i���/2�^���� )i`�m�Pތ$Q6�)�y�H���CQ����gY��!Dd�M�yL~zZ������$$�B� j��֠���BPF��P�^^����iN<�Se96�3 �5�̳���?���^D�$��8e�:�����ܟ<���\�F�mꓗJ3=	Ezj4z&*��22�4� ���NҝPǂ��ʼ�nQ9�y {.�5+���F���G���\ �FD�x]U��m�P  vd 
w�ǃ�m���d R�\��
�*���)m��j	�x||@[;��FH�d#����,�[��*W�4�8O3�@���ݣ�O�P�`�m�V���;R	g�ء�2Q`R�4��5D�nܸ!l�{{;�� 1�������H�e��r�?��Ԍ���I���(\=��EA�$�;��q�v.p"R��M��uy��"�P06jo)D&����,�3�:���fC�5�>� "����rN�ހ�FƝ	��<x-< �;&%��
QqL&�Ht�f` W�������g�@���T_��?������\l�`���ћ-
Sc.T/�yf}�_D9j���1�7�;�kFaH�:'�	��}֗hB��eru�6Bdx�NN*@I�6M30
ԏ�$#����؞v��Gg�[��g�G���u��t��7�ZJ�g�y ;���m�)���`C���7t���~C=�SwG��%hh���!m5�\8�e��e��%��s�i��#�yT���5d�+UF�T�zc��5R3vkbWHMT`0��Fw}��쨋^�k��Ù?�xjF� ��vYO� F�٥�C����.4D��	�m�{�}Ԡ�6��`Of08�}0�|�� �
_}�N[k���o��	<'`B�t�*��u�#��D�8JlCce���&.�*��[f���m�2ɴ��b� ^�u���
�;>h;�ӑ�Jɞ��(:@L�&�"�� ��4Y.�'^|�>���RZt��mz�Gߥ��6�(`|�2��'���Ky��e���(���loQ!��r�0��=zL�GM�f0��z�h��и�p���,��o=�������K������e�aG�>�-��a�n+�+D:�,礇%B������R����	 T��@j�3�F�'�ތ�5�E��K�m(k@Q�b���s��3v��U��=`J�A��!'�ҹ�x�N������-愝��ߍk��c��#��t����)����MD�#u,��9Owo_�;7����ޠn��%i9ș�8i��3���;����Ѝ�p�T?l.�����:�W&�v�D�Z���s�� !^d�3sl�,��y�uYُ@f�s�K�y����J�W�P6�/As��� ��gj���x�)�4�:C���Q��cGO�mpy��(��������7�e�J����c�����v��)T8s2�x,Y2}�ڗMR� |ı`�#Ҝv"�rc� ��ڹ�t�_Tsf��Xı�'4�w� RLMB٫J[w�Ҥf�7I q��#7E�y�,OX�bHd@�ʆڣ�Szi�R���,�A��б�����'��|!6��ѹ���w�MuI������zZ����U)#���_���2�d�^?N@���I<�vO��C[¶��/g _��ן� �����7WN�t&F�X��*Ԯ�I��84�~"�СO���V/�g�g,iԣ!���Q_Pd �>�Î0��a�F����������M���J�,�H!D�;(k�	D���d�9! �ښF�c��w�>~B�j���0�VK51���ci,���񡐋�^�;[Ġ)[�P�u��"�BHE�8���a�]�t"�@�#��@P���ҏ_�1--\2Ѯm� = q�L�F  I��#�ʟE�����̊��硤S�I=X9і5oP���@Pڗ��*��r�qEҍ�}�]��٥��-Y�7� 0������0�u�|A��O��*��o|�K�~���W���W^yE���ْE��f�(L�bϖ��j�g@x���A��._�"Q���=1���0n<K��)��z��7L�X'G����2���
V���|��ԝ B�Z�>t#���?sxp@��S(��Z���-�z
!L�痨��?�3��i�����%���$��f�Q�?�3/�lStm�a���p��"#9<��vR�g�2+}�1=�k��NN�Z��4�D��Ɏ׎�̦ROe�m�k�N gX�*`г�`� /#�=;�8�ؒL��J���s�A�֋�����8���^L�%��ɵ�|���G�峟����X����cǜD��4T;;6ͤ�kfyf�x�tu�{����7�g��~ډ�|���$@d�7� ����D1�-[��[&8��w��@��Fj%���4�GySuz��޽G�n�~���5��ؤ�>��Ͷ��y��,{KS��qЃ�DI�H[����4��kcGDfc��\<ҼW��F�`�)��	�	-�O�'�R��1�3.���B|}�,�%à*W0"�F��vML������~��kYZ}���Cj7"�O�ȗ^�#�� ��2�ǸXy�=l��� 47������D?��߲��*�th{g��ֈ<��r�>��O�?��ߢ/��ѫ_ߤ�^��nvi�;oҭnSmf�uI��<y@�+�������,򵖾�鲬�XGX����vG+��ȓ�w�ڠד��� �����H#������m��H�L��H�fhϴp�L��ֵ�� )4�0�6�TAI7x~Օ�l<��[�J��.���&"(��4]�}42m tC��f&�t��-��߽!$5`B��j16�����)[�>c�< �����'#-(��
���M�"�'��
�p�����u�F-,^�:��]�S�h�n���*E���A����Sw0�c�H*�h��G�x��;/���G<��,y���8d.�{~��ή-�m6��?L�br�M��cl�"B�4�r7^L��5���U��ҁ�ߜ4�SJS��E'��Qόޮ�s ��I����K���z�6�</Փ���c�-�/[�T9��������$�=ؐ��� ߋ5}
��(0�=VoS��3	~�����yB��1�\�
%u�|LZ�f"���zwI�,�Ϻ���s���k���($��6�,^0��8�c	�L������f���>Wo�M���cMQOa�u2�jBqآ}�݀:�Π#u�e�� e�V�cd�l���B��^^��ׯ�����M�@�~��M�Q �BK�TED�<0��g�޻GD�z��Q8m ���s0�H�t㱗���0�	�Z���>�^�HIĹK�2U
U.96�;K]7��r�n��uc��I��"��9i�����I���Yò�g���H`` ��3�3;>���3��/	��������b��r�J��f��Y�(�^�ej�<э�3S����?c�X��ʍ�-z���%ݳ?�x󦖦H�|�A0�J�,L�a7�����%p��0�.8��is��o�N�b$`# ����?���ߧ���S��?�����yOMM3P����{G#� z���Š�X2/�%����=��[�~��_��?�����V�}6B1~}��#�) �����8L1�ݝ}I���KT��%��>� � ���� X�gK�V
��B�}�L���;[H����C/i�MR�I�2u�S�\�)�f�{^�+�����	g2L�\q���K���ߒl���A1��ieҭNޞD���&�I�5��
�}N�a��i�t�v�$��9���q�Hk|ϰO���I�hM����0��wP'k���*��b���K������LO�E��0P�&�Z߂��U�`u�U�v#��_{1F�,�D_���>��F3���rޡ����-j�Q�q@�vSz�^�s��ߺ)γ������z�Z�^\����)W���� <<�:,���}�Ǭ]��I�&C�(���qi/Qf�^j�<�g��=��eb�8u�eA���C9 ���[�tk�?��L�V���9�Y��s4����_?�^d�����;V� G�|�&"��o��b%�67�i&7A�Ks4}��w"������E�}e�fX`�)��R��Q}�2M�^��_���w���Ç�x�.�T��x}���k���~��R�g {�#Q�����[���7�%�10X�&��G�K�����x��d�Y��H���u7������u�v���0Z�=ṛ�M�7���7l�b��(���a�ix�(o��xR�ށj�B7o\�RN��b�����5c�i�12�C8��7Sf�~����w�T��bYW�����S�&%D�̄�H
"'pT8H��3JA,	��8˛����W'ir.F
j��Ӱ�q�A�T�.����"1���}�Q8�nP�h6(0��vm�{���3�P�b=N��6�N�Q2�Jnho挗�T����2�;��:
=���ee��VX�B�u4uc� 1�ʜ+���v��[��ݠ���eSc{��,!�4Ԥ/���62>v4g������}F�{f\^�3��/d��噍��Ka"I-CD'�ɚ��	��"�fU��=h��37�m�k�Y���@4vk6�f�&��3�L�:c JG�Ǝ���9�e��x�/P�����V�q�D���$��:���2��WO�]�D��(Q��̗�������$ED�[h zd>��q� }�}$������O�#d��o��\-��α�v��u����_3��>�������$2���m�i���T�����$�Q
�0x��o|��Ϳ��D��ƻ������Ƚ�y;������ ` �
G�m8���3�S����A��2mnl�w��]������C�k ��]��B�R���-��NO�P���{�9��?�}a���W�J����O.�P�����wW$}26D+�|�Y0h�����wo�o}�W�����:��O1@kS��egs�&���3/�~����g��q���� ��/_b0��45Y�ͭc��W�F���7\�R��sܽ{W����82NV�V<������C�Hd�Hm�ښ J�[����{��>u���U(樋�L������^�2����/Y� Mgf���魭uZ_{F�������Rw<�3`�ian��]]�L�^�E;�<��O���G�뤍	 ����Es�w�w~�����U��3��^�o��mY_]}�>Kg�"��K��l8�MEd���8� %�i�'��qbKjz��Q�{��3Ȍ;S�EI�f��=�Y������o[�� , /�4�l�X#��p�M�cƏ輳K�M/���ٿ�#}'o�4Қ-�{R���cl�g���'@��o��!�qt:�
$9%.}W���u�&�Y\eg�b�k'������ظ�	D�|ve
��	��Nk��J,���N�2 *ɝ&i�d�zG}�o�HtLJ��2���� Z����f��Z�Z���n���K���G�p=S������Y�,^�F�o,��1t�~��gbX�2dyғ���<�4˴hS� �e&,Q�R�>T�C����8���6�J��G[ ��~���~I��yn�6��� s�T*)SXbP�E���7)lnS�\�~Ź�/��l���m�@�S��E�D#�0�M|���?��0ĳ��ۤ�]q(�2��m>b�Y/!�ՍUZ�٤B�J!�10;���
i���3�|�e�Ǹ'��},��&�%d^�Rv������@ӴM�9 ��75h&P�?���!iJ0���"�J�/��J�e1�6��H8��GB���٪d�L��Z��}��#��(̸�D��2�rD�G��E�A� �`�u+�*�L͈�\SMmp��_yɢ���s��ҟ�m�@�cQ�R���g���8��&ϧA�G�A;�8vF>v���5��$��|�No(c-�'if����ݡJh���@5�t���._B��vQ�qآQ�G��u���unmBzc!�c��m6+0\!�8��w̤�z�K��|��������3}����E[p?~DTO���S�o��M�;s(��T$J	Ur��2���OT������9�=f���i�uΐQ�3G���O�Q'���K���U�d|�5.|��a��i�Hu-#��������Sh�,�5xB��<�fO��3Tr�4M��b��j�VM�ցH\,�ge�Yf��w�{��*8��#q����EƎ\#��CI�g�n�;��dS~lJ�e5G&v�{"�(2D���16}��I���2�J4	�����ld<�{r4 ��F-�l��HWNR9����P�aoHC8,3�C�q�
�牚�z}B��uE)mon�����gИ���$���?�HR��J�B���.���+t��5��@��Ezp���E�����8nnl�y�O�X*�E�/e��ud��Y�=��d]�Y��JD7�mĎ��Q�V<��J%�f���P��ln��`��������Q��r��2H���i��x��0b��T+PC�)5@�q��ss(颏?�-��F���ϳ����WD��Ҿ�#��o*��ޞ#��33��ܜ(q�E�������!�)W���;w��_����P�#�-���u�ﾻ@���B�>Q�k�(�����p }ˀ�P],)������H�>���3�k���!eX7#�2DFBQ��!^�ݾ}��z�6xͬ>}"��B���y٣��4hv�\�b0��)��0�k��έ��ǐ��?���gZ'�2l�&�����E��O�o�4D����3��A=d�^����LHw�������I��c�ڧe���ͦ��ĵ P]J�M�X*:*ΤHR�M�$9��<��a(Bc�IO���u#J�&�0޹��Y6P�ڬ�6v�ߋ�N(�L��B����S[2/�%`0�'�\z�tz{���q��l��R�N�;,y�F���S���ƪ�ɖ�`oK!ۊ\�m
�yZ�}}���%���#:��R��A�ݩ�%��t����Y�>�Qd�����7�G/YjE`�8� ���;Ų�痖f�����	�JQz�V�Y�1�˃\�0�����^��p �y`�n`]28���gԦO=�@9��XF���W�����z�`�y�e��^�{{�t܎);yEZh,,��?�� QZ�Wu�;�����c�:���Ǭ�4�4Ek�k��׆|������u�,SX�L�0��^���X@�q�:|H�P�I�I���$��4L6�F��ͽc�|�y�)�
��HOC�UI�*u��#�/��؀�V�>��|�y|�d�4��)������m߇e$���)OQ:l.�-�(DIrt�e�W�8�[43fp{�W�l�&UQ?9��3�K�6��ظ��0��m��^"P`Q25f5�N !��QzP�C+�X�Ld��<?���}D��]��i����,M-���+�<𤇼��ןH$ofi�J���a�rԌߦ��4���sd-b�����X��{�`'v��������y�Ϝ����hf� �.z~H�(�ʹ7=�d�Iȧ�2�L
�Ώo��o��;�X�t�dB����ŭHK�C|�f�!9%X���!v�æ�����R2��1}�*=���K��������[�3�8��
��6A!Qu��BV��Mxt�Bv������`�t-�����V�C�"�@AOd�5��睾�8?��u���׳��~�5��9~x]T*R!m|�t8��/4���O��$�X'V=�CM�p�5�,2)�����X�M���9�ߐ~F`%쵎YI��_,�^ �e.[��?h�~��=���{�g��`w��=~F>��à�*�ޡ�]�Z��`Ez����Q�l}��Y�"�}jw���+t�
�Xz��ghm}]�A
%��$�����H �%���#�6���0]�1ܺq�A���H�<��j�&2c�|�y�&�{��D�P���1��> ��G�W�\��|���|��k���2� ��ݼAˋRӊ(�C"2��D�Ld�* ���1��<�����6�-1fj|�0��n�=3(�</�wb��Ź��0�j6��W^a �����w{bvVgM�CD�������*��s\�ET�ez��u��p��@k"��PRB�����d�� P�*o�߃����o�ߧ�����՗�=���A�O4P��:�g��V:��0�P���"���%D��`��_�����mz��?�e�Sb�
^8aGx�Ķ��0H������^7٨�kMO�'5si�e�}��إ�S�s4���d���Y���� {�0�Ʉ���b�2�i���=��T���MC7��K��G����z5��`H&.KgL.Y0�i0��x�gm�ѧ��=�Cp��E�q�Dc 4� �d[��]�3��s���ӠORC��?�"�ASN�����ȩ�����&�?B_��u"���D�w�K��o��	j�Nl���ı
��wnK=���3��ޒ6W�vS�����
���%�����[`A��&��!��,��}��ޗ��3c@�����qj~�mf��޼B^J��m��vx.�.������=�:��l?g3p�.y!H���N���C�sp�"Ч�:��s�Sf���(;l� �2?p0�����% ^�P�4d*Z�z�&�,�]���K>-�LQ�����h�~�=���j�)����I��+�nOX���w����vif�N�<���� u�}Yc$}	Ņ 0O�
di�Ɍ��#�΁�ؚ�&=Xݦ;7V��T4��H�.`�Y�����H%�9=e���;�}�Go�{�1���-Ҡ3�:�	��dw�M�e�IF����s�5ڐ��ZP�9���� �4?,8k�R� 0���j8T��|gPBY5Y)��̄1�IO��Cf����fg%���W����$�M����VE2����?��N!W�S�}^ĭlH�V����wW�d�ML�Qmf�z���]��x�I��u�&��&������I�I�Mm�����V�K���gw�M=�O˱2����V�f�����k�ˮ&�6-T4�2J���	��4Q���z�1x���sf���_��7�y����&/���U>�cP�O���pLע�c����"�3^�����q�u�_%M��	��
�\h)�d��6!�У@�����
%�d	j�1a��L��m�ˬM>�I5�[�i<�4�Ga�W)����s|�x�����%�_�N��^�6������o���"��E�#�`�`D�e�5�WKP~GT*�.��ɺ�P�j\D������ۦr�(;�tx�������w���|�=� i�KC*4�d�v�� ��ld8������V �4���SIO
I�cO!�2�8�p��,5*��wH�7�gC�%u�[k2/h��'��:Q���y*(E��&�P�i��������w���l���E�CNC��/,(�B4��CV�!#/г'��������`��m�c�[�X�#6P��/|��V��2�`�Ra�a�A`VR:q�?���������67w�Q�Z�$
2(��ׯɼ"u���KKK���A-D�2?���7noo�D
+��������s��Y��/�%���d��P ����}�������D"C���ӳ�����W�L���ol�Q�Ցz�⌂�?�ʟ���_�g J�� ��T�O
�A}b�~��@KKW$������<��R,�F�#:  kk�vv���F��'Nv7\ߦ��uz��M0����F�9�� �#g$8�9{�dD {b��P���C�sb�#:��3�?N/��I(�Ƿ��Wډ�e�C�X
��(���5�ii�~Ei4�r'O��8H~�Sוa@�I�Rs����ϧo�h��y'���:�ԒϺ?�{��#˘���ܓw�;O�n�U�}����.�����T��-�8��2����hXw���|JHh��c��)74�Q<�Y���Abz�zf�=5(�k7̊|E/ԩ9W�eoml����0�"�%S�.��{T[X�>�}��@�,�T�1�"����۶_���j��o A,:	�'�/�,��5�u�
�Z�w��7�Y4��ē~��}i�����0k��,˵Jy��+eZa�7�����Nd)�?��Ă�XZ�R�P,����7��-ݼ&m��\@%�5�)�c�AoH� 5y�\�09K�ǢPj/��"��/P-_4̴��Ox��P6ij����)�	eYÁ�%J6�5X�(w���M��ʕ���d!s �:h�f}��Go?Y���kTg���%��q=4�G?KR��������?}����P'�Х�����y�+�	�����4H�p-/�3�F�6��4/4����,iʗ&�yl|�����h��K�m]NQʛB�h7���������W��-�<*zE��
+��o?C���W�4m �i�M�ȚT-����+R�����I�k�ʺ�π�'|��tfn�.]�!�ex��-�Et���%����/9J�t�;N�$߄��{�E��z��ճig}=���zF_��u��(e�Z�u�g�E�<��@���$�������U�����M'G��c:���Rf������?��8�L^��˿��4G��z��10���x6%�iǛR���SbL��cl]��(a��:W[L�{�a���c��������y�B�w?�]�3���m�qVu��R�[�b��gk���wʓ�y�����T���C�b�g|I��`P��0Gۛ��w�ԥv��2Xڦ;<��2a�$_��PC��ax��_xQ��{�'@p�`�����I_�Q-�.��K#r�nw�Ê�!-�� A3�� �
�j1�����+���])d��J(��tM\;`ez�c��|�*ݻw�����֛�����W��W��+_�:  [�o��cs�M/,
x���$r�ۿ��"W���ߧC��h��F��O���N�JT��3+���5*�+�wآ����t��/��o�͛��ۯ�%=��6뽢l�'|����<[����WQa��VW���_���.�e�싿�+��W^�*`��~x��4���6���-��￯L�<G/�%a1�f�u�~�<�R� �v�]I�M�s �	��o��ohg���x��f�%�x���Zͮ J0��o�д�8��r�KG�=���d �D�+�#�{k������+����}��ߣ�_{��lP��@�"�swnї��?���6����2�SP��6R=��y�Xyc�E��N9C�ڿ"c�pN\ِ�����HOV�Y�5����~Έ0���B��7uD�:�PKT,A\�����.e7�����I�l<�'E�ɾwN{�M��H+�k��2����^_(����ǳ�觝��z��ͧ	�9Ǿ����h�Ē�*KDx��F����}�;��lq��~1`��8L��܉ip�+#=3�+��Gl��s����ί����_�N c�J�Lsփ=�oN+ ĽU�5*�F����U:@D�٠�qC�_��GWnݥ	����HZ�xA趗�ёIO�=W�e�`lԵ��Ż����d�Ij�5��K2�e�������8�m�X�������y��^[��ty�����v[�W@0��`����4S��N�oQk�:�	�T� -`�Dj8_��k���5k�-�;�¶�X��=�	�'��G��;���ŲVK�P&�e��T/|�7�ߦ;w�Q�\b�����E���cv(�{�L��Ȅ���S���m�DV#�M���uNM�U��'4�/?�(.�Q�Co�s�O��+���1B�.)��Bg�����������|�����B��h��(�VD��Y��ju�9�^Nw{�@�,G�.��y
Z��7�^U08AS�|ZygE~�<����!�������m�76����x��Q���[�^�/�g��l�I�$�s媤�H���v@���l|'q˸0K�K��DW�vK�l�� l��ak�>�����P
�[��kpxL��f�/_�*��7���:��V�#�N�T�z*�"�����'�a�Xpv�gΓ4M,'�yj2O+��6M�Y��]p}k�O��ӌl���h
�y����Лi��3NN��TO�u��/�ݦ):Ϭ�|.}?�Jj��HgN�YJ9�2��/�ΛU���$}���Ⱦ�����M���Ή5G)U��Kh�������a��� Hy��z]t���M����|����_1nۚ�E'��4ݣ�#� �5�rk�(����Q��(�/�(�j��Λ+,0�]�9�Q�V6Q��_��/�V���w:f���Q6��BD�Xn#���ł(i{���6�>����˗��g��]�m(Fg��*��L�*�	mBe������:�g|���=G���_�9{���� �������R�:fВ�R�6)���iI-K��M���:d�3���x�
����^�	�#�'b(����qh�>�x��!W�v�G��7y�]!��dd�<�y��4B���҄*B�'�}���ˆT�F�~��7����E1��C7��<jQ�Ġ����(ԏ��T(���ý}>oI�K7�=�ݽ]Y����y���҆��J�.2�!<+�<�/yO<�ܿO=��������*���F2<��x�c��l�"��#3τ%�������牣���2�=><`�ٗ�C�,�n<D ��ge.'@�+�����,W�@
l$�k�S[�	���i�)�QO4ܝ�|�>�+�����g�����A������Q�Ć!�H�sn�gl��Uj�-�^ȵ}c�X����Q����ޞ��M'WY/��g���L�6Cs�zP!c�\�z������fp�xQB̑����F�f�zl��s����Q�|i�9e�N�O}���g���H�Ư��,=Z�����6K��v�q��H_/���"w�d��.m_{�-%en\O���LLU���e)��wbbJ��M~���u p *��ou>r� <��؀D�BC�Y�j�i�en��U����͙K+�p�&�g�����	��B�>��\,s*l��X�*��
 �<��v?i�LP���m������'J����b�J-s�:�*�S1y>J�GFTb�z�B��"]���1=a��,
���6��#�F�4Ä��_>����<ÀlZJ)�vYs	s5�a�i���0�uA�K8ŷ�~�i[���u�Q:95M9�ŨwL�L��8��ب�2)�=��5�,'s�>��0�()?U���L����-�dy�S:�1�g{G�w>����"U��,�y���RK�gitG����z�-��w��@��^�A��W��s^��Xf��_U��!K���s���95b硰}(�c��W��9��pY���� ���;ާ������������Y���}UW�� ��i��$(�D9�#�~h��r�j�j��tvW�ť~�(�r��Ha�F7�[���.�]�*M������""�2���s��*M�{/^�{�k�{��	���碣�T�`�m-`��PZz�q�TU�K�H�9��K��c���!�)�j�)Uڅ���L����� C�`�_-���#����YeDh#��PIrd�.|F���PZ]���-a�K�t�q�Js���0E�b�5M#���O�f(V��[8���JSl�41���^��7�}�/���_jt|�f��u����͂���~K5�llл�����
����<����o����{M�=�Oe!5*�o~F�����hX&2e��p�x��f��զ"k`Q5 ��l�ϛtd�o�G��Ԝ�7z����:@��g>��g5�\��@���S�N����� \g�4�d�w��Ky[��/�����-�o~���%zz��9�đ� �+���s��2�=w�ű�G�! P�5�-VT����q-[�(�ĕ�e� ��>�៺6%�)6D�=!��e;�� ����g�P)D��ў+J����G��f���>n����oJ����SNi�V�C�h��ud�9�"Gm����(.^�( �����~,=��XIe���3Q<)u�C)6�-���n��ccR3899%i�6)��>���t��E��K��YY�%}-H&��#ފ��^�v��҈�-��իW%��5�x[�N�@1����J��5)���ڶp]"(�{jǎصc�\7N�T���a�%���{�Fa��o*EI)��S�LCת�Ƽi�D�8�J(�������095�˗.K*h�C�A�!�{UIE+)�a+A[[R�� s��>���p�:;SH�<nL�о)H�5��}���@Wov޴S"�k���	�)ʍ������*�8zh�ܐ��|7m�,cZ`g(]�[n��=� �ܴ	˙]�)�{�`����`c'ۦ�_��{ϩ����]�����?@��bLWu:���/]���_��'h2<��C��/ki�8�R��h�em,��Oyl�ֺ�IҰmZ�7��!�w< �E��'�l�l<�>X~���������8��M>��9�@h�0=����ld<\��}t]��ԈP��� ȵ1\��C9��ώR Ϳ&��+`��o�6�]��7�qHn˟@Э�W:#��]�K�ϔK�zҪD��,wxe8���2��k9�߃B����]=�Μh8" �	�A���Z�r��:�*]��s���� ˝�cJ�4+k���*�9�#�?/�LS �I4�
�)npT��(�8�O��ʒ\�hY�Idri�+ �S@�ދ�EI�X��1$��]� z�:In�B#�ƺ�8�H,i&��֊-s�@ka��«s�Z':���f�m	���[��*�q���m4�����e\kt�2�;�"QA �r @쿱*��AG9�$��(}�$��'�׾"�7�0�{�!F�dl�����+��SȔ�"]�J"\U�"�}�g�L��̅x����-`h�MH�#� �#��6�g���D��2�d�� ��2�����)�)�uM��S��̜6�]F�6	�%�����f��w#�.L�O�*��9�P�J�	3�10�0yc�xS��&!����p��2u�kP�����κg���p��A��2}������8�J�YF�P�L�y�?�.�\D�KW�o^�F���a���L+�MS5�Ui���jZ�|ʲ��&}���� ��t��`i�hoX��2�h��\�1k=�����#^��{ \�]]������uxJ>Оa���;CBT�V��w-l�p6~���Ȼ�j�������Rƍ!�;Ns��,������r?�s�>Yf-߳Q�<Xq��f���WN�vϸe�Q��~Ϻ_9Y�Qr�S��\����Xkl�ȁ����D�>���� Z�Z�vvfW=&O��Q�@N�+`m-M
�Hy��H�W0;� la����[n��#Gp��E$	�q�g:�*��!G��G���]7݄;��K��S��q�]4&i;�B	}t�Ϝ�����Y��r���@�����u!=ٽg/�y�Y�c��`ɽU��e��9����Y�����f>�0`ضm;|�!P�tV�O8��2��o��#G#O�߱m���,�J(��2S\���<�(��ݧ���R����nհu�q\�>��׮JMa["�?�dr_EC�C`���=�)�|-�L�k�Ν�����L/-�HˆDK�/K���M�@{�=]�R��Y�`x|�5�V�W&�10�S���Z\Z�ϥ$H�ָ���~:%{&	�������ۓ�%�g�t��)iq���y�޸1Kǎ�8�d��p�E^���*��":�1�f�I[	@�98� ��)Yt���99�����¤����XL����uK�P�����ض};�;.v�U�h�Lq�Z�홏/M����!ea��,��{P(;�,��f���|pdǆ�uz��,�\߶U��T��J�W�j�����B�X����/��s���_����)̚��t�d����r�U�#;�M���kf��� �!���k�}:ۯ\��+�[*�j�c�k|��c����6ҝ�6"\g��u�v�k�u�א���8N��][ǔO�K��S�����ZZ��9�S��5�S\�۱��8v�&
���P��x#8�V���{8Y]-������\���ӏ�����i�\�J+��
9;��#�d��j�U_<@�T�@q]� ��y�����v@K�ʒ~��Xɚ0
����H��dz:��8�B���U�*e!����8T+9��ҹ�:���H�ng�'�>�2�6���j�A2D�����9t_ˣ%F��Ul�U�5. �й�u(jo���S7�!�������7VFzm���-X�h��0�޷��d�S�9�f��Y�vzN���5!����l�b�>�!;��^tƏ��\��b	�T���"W����\����d�RH�#�f$�i�����K�6=��l��B��/c��+�l�%���FH��+�dy�nd2Jv������{�����.@Օ�aP�x�J��0#V�EV������������+�⋟{�ˬt$�IiEt}��$��HU	�Zy�~x�<�]�D��8��HB6CEz
i�ԻI�6~�b�7��nC0������t�*��%�&J�.N�3�(�|e~%R�L�B%J7p7)��D6m*��V��,ZA�0��y�M��G���簪�@P����ּ�F��u`�ͽoz~uTJ:�� w(��g���:��:�������ST�R�0�!�1��Z�#���+�ƛ�h�
е��]\����V �v��)ɪN�Qko�+�����Av��؂o|u#��g���z�S�}��� �)6V]�_w
U��K�4��]���L�P]2j��ߪz� �w�����X�omȱ��?>S!�VJ;�%$�tETđ�B��j��{�2����@P�Au][H�f�ːnl��h$��_�_|��O@�`_�?.o����f��J�139�}�k;._����**�?L>�Q���.RBQZ��&:��I�1��Vit�Z�Z��j	�����~"O���7Q� ��r)K�$�&7)7榐��I��k������W����?�!���a1Cg��	2����uKj��J��
�:'L�/�?y�w���_q�p-���q��f![Dy1�L���礖-)���B�|��:pX���B����8-�:!�m�$�a��� .m!�9%�<3\��ƾFrN�\S��v�5d�c`@�G������z�R}��$�SI鯵�� ��׌�0-Z�H���HHE��wt����:��%;r��R�L��#�L�ú7C�ӊ�,i���%�jf�^�
� 3_j�O�SV��ֲB��l�Ւ%l���N��Q@}2q�����Y����`ג��Q2f��Ê�,B��V�+;(�NQ�W/{�UX�������5�Z�h�73B�G��Z+�D����'�w�k���8��-7��8]=�i{�i�\�-n.��j$�Q�C�(�L2h��i���j��?���8^2�e�!@Q����j�ܴf�~�ׯ��E`��{j ����s<��_�*���u=w��W���O�RTT�x���I!�1J��l�rJ���pk)&2��H��s�s'����>�s�~� Բ�+G�9C �i}��z�zjTFJx�T���)R��:�$Q�X��-�w���0 ɶ�Ә����ܼ��`���� p�9�s��� %��ޖ��ζX�}�R��,�m�$Z#ݒ�RX+ O�(_��-na�&8Ox���$�o�Z!��.��m1�'��-L6;�#}�s{���/���^������[Y �ӰR�5�L]E&X��� l�צh=�H�rZ�-�*%��C�t�|!��<�8��^��x��$�%N�W��jOK꭭K�td��h� GOm�R/��/c9���W���������EZ�P�0���Қ�	r7؈%RH�z	'�˄S��܆���Fv��Ay�<$��l�G�b�QD#�%�*�o!n�iM��M�a��*���;z1?s?���Й������@g�4h���)�fÖ~X!EC���G?�?��&�]G���D;)�VI*W�P�)*�*>?�kʹN��W�r����>p!��c3a`9�XU�kN�C��ˀ�J��=^f�I�����"X���M�'�<<,�49��x[9�t���/�V�խ~@f@�c<�V��<T���m6ph姿�Ek�E]���|�n���1���/[�z�hEᮻ���t���7�\��6 O��	Wٻ�/��Ds�|���׎��JO�y�|Ə��:���F����4*q��ͣ�>��Wj���wi���	V������X����6�s�"�&��1�<M�Kl������Mv�i���U�&Jkz��yq湪���V��9��;�%��,��-d��Hq�7��*��,�._�I(GeoH?+a4,���� ;�Ae0�u�/GŤ/�!���ÊԿ�)0�k0;��D� V��-��X�%R���֜\V4"`�8��|xf%�WՑK,��	[����s+��K�z��]c)H���({��5\ El�/� ^�z��e�l$�!đ&T�R��/��Fȫ�
rW����tuRj�xάhC���׏#�����
�3������>vZv3����8]���{irFt�,�ZF�"LP������,��0�2�ktmצ��Z�`+92dH����=:���	�ZВ���S��dlT���(	s�n;���G8�Ŵ���t���!�
���WYt;;��ՉI�*�����%�a��3���J�P%��p�H	�Y2Ȗ�VeOs=�80�9D��3�*�G��ڄ!����p��'�N1�m�Te�e��מB��LՍ�h�F�:�za���lj��i�}�Sm,bl��G�4��#.I\'g�X�\Q?V�9���q�A<�/��]ag�|���Q{|��� >�u=F�-�V�ƮO_5�p�n#0h�,1�]R��
o���P,�%���#�մ;�|�#�ˡu��6�B9B��#��%W=�F�Uq�?MU9j�mTzӱU^&�8�)��g-��Wu��!���cB���8���*�0k帺M��Q�^��X'ޚ꾇�����rT�)R��0�2<��;F�<7Kr�Ag���X�/��2%��/J��
��8Z%���ߋ��1LNO
�G8o޾.^���}7!D\ǥ'k�@Q=]�[[]����mqtu&���o�2$k����d�ֲ��b1��x_�$�JQ���G�q��q�'ضu;B���}+X����kg��3֋��Y��X$=E__l���d�OLN!��#ٻ	�`�n�����LA|�I7��e)vp��^9d=j�K&׼I�G*�'�z�4.��[joE�V�L9�T9�#�����;��eL�<9E�iaHoȮ��V�$�,�*ׁ8:��SE�$vETEm�/G���ʒ%D2���L�����4�������۷����oW�ʈcC��gc������+o⣓gQ�#t�R�P��{���*	r6�~��=�,%��߮B�	�F���,6]�+y&ap�g��R�N���2#jy	%B����!r�7�Ꜥ>kC,堡,v���L�D h��<��`������1�������}��v3e��_�Իn=�2�O�AT͔��U���'��S
�4�-f,~���>(�TKH- �w~ud�ivv�'�Mj.=D����hN��'Zp|�j��^�����~���4���S;κg����m�fi��h��*��Υ�ZT׈بf�`�~n�9��F�e<�M������?���6��;n��>���)5�R��체Z��2�ˎ �2;������ei��EP"� ̟�y6N�z[���k�r{��.��H/.�#������B� �$S0�tA�,�=���N����6H�q�&��8-'E������D�c�K�-����xX�*	+f��D�U5������(�8SiiA{6*Df��tv!�'��Iʜ#qRo���x�8E<F$��jN�a�ˀ��8ݣ���*(��aI��B۴U����uZ�I�J��K�
��2�bC"��֭��' �`lfj�˫������\��! ��Cc��� ̓a%��}�r��%�ܤ:z$͓���sHvvcddL ��ܜ��y�i��*Z�Xka��#�\/؞l�T2Ne�p�4��`ۭ7�އ��I�t_S2���tc�+�ud�0J ��;��m��*�����G!J�r��7�����0O�P�|��N�<yZ�̎X���Z��ݢ8���O�=��R/Xd�G0h"�|�پ{��������b:�@K���j�/Y�; ���3�-���ɧ_ߘ�s��E�l�9`)Ԝ���(,o�>]j�l|TwxK��\���̼k߳|�~��TE�k��}��_�)�&cɵ%��L�4�L��d��	hL��!���;q��I�rSx}>�F�+a28|x�u�JXŁNU)�¤�� �)��nV���a��JU�4-�QI�,�K�·V�=Ñ(#$�x5���Jʶ�����F�`j5�e����0u����Er>H?I��;6������{����$�Z�6nٹ=���;̑~Y^\ٓ"�2:<H�%���rX�^��|#��J��dG�Z����ʞhGoO� Bf"��x^d���[�u۸�\�>wS�H��$����EZ��<PX^�<ɝ^Z�i����^AK4���Q$ڹ��T��j8���J9�B(���14�Gc��	ydғX)E0�B��V,�U#Sn����$Ji�P�L�2,c鵷�f�~�����̒�g1[��r�뽲��8�m��"��"� ���;�NEے���eYL2�A8w(�.���@�n�`2�����(�в���r�+��M�!J���6���L���$���@����.\�C|
;��^K	RA2 ��Ә���G���7�ƱS�-�Ht�L�ҏ��J��l�D^7E�\m�S7�i��_ߺƈl�pR��Gz2�@`�.�1�x����H�3��*��z��b��H���?!��idH����q�Ƕ,wM\��*G~���<����_1 ���7�C�ś]y����g��r����gԌ�6���w�ߺ����ѩ����O���i������Ɔ�aB�R�P_��T{���R�c�g�q#����k$��[N��р�_�7/}\? u���D�1*=#�����5DM����*CQG�e������o�P����[�w�)��n�O=�0�o�$͆�}�<�I
]������U�	�HF�e�J�~��Ȭfq}z
�=��~��R+���?&�UOLI�F��G����1\���5�>�y�f<�ЃH��������S*���c��"�����o�����Fpaa	��#GH���s�.<���%|��%u�A^�$I�xR�ǰR�4&���߶G ���G���kd�{�}����'�\a"R����5�ĤW�j�E`n߾�05=�c��	��M7߂/������o��K4��rU���Ԡ��<��gp뭷���ia\�������(��o�%�*|�O_��177KIA���h��Q��rۋ�w��'������ǎ����8>��_��?�>.]�,T�\K4��ՒԄ���a`����^Dc�Ul�ڃ�}�M|��C[G'^����kW&���X�������]=���h��[��c����%��f��>y����c���_���4��;�Fr��k_��+8q��� �qG[�d!J����bC��d���Z��v!��M����X��N���/6�9��9�or;R��J>���a�!XVj>�x�^;�N��q���]�An#����g�{�Z?\#ڡ����l퀶ܱ�.�u�����k���(�,�`� \�]U�}3�0h��{�f��l����U1�\�5��!\�{j-Ԝ+�-�^�8G�+�7b	�Ίz9�kdT�:��E��l�ڒ�����JEW��Q�-�8���l���a�K��ZD�L��N]>^Xe�tD��饀�ΩQv5�A�Q�~�]�3jcz�C1��u �)t�|6�V�������HJ��޾~�;zp��E�t�-����9!����9����N��|^�Sa��p���>~t�(��>ߞ���:qU��ѭ�C���4[XZD��_͖�.TT����B=L�f�& ��Za�+���e,�e��%�W��P�D
a��k�@�����>���wF�IKj#[v�µ�8r�tD�e���
��.�t�0H��!�`T�%�"��'5����L�-Hc��c�ku����C1�3��NI@9Gy�����8��F��l������d��`!g�2U&�6����B#͓���e{po���4
t��:�98�Ź����y���Ħ�1B�����c��5�9	s���`Ivu �� A6��8���n"N�/�x��l��Xp�|^}�<- 6��7t�q�"{��ev�rȟɂ�"����.:F!GFP&��Z�.ZQ.6��\*��6Ѻ�x����|�(��#��5jJ���&}���҃�_��K�1T!��-V�y�g�����}����i5)�2}��@�g����0�:�y=�bnN��� ��yÇ�R��������F�� ��4)!.PrLZ�%d�*c�ҊZ�7�3\��hRL��/�����qkc��QA��.��[I���S=�Y���N��C���t���S���ox�T7ȕ����M'��t^af�!���_>O��T?1
��8@�Y�P{-��⋿��?�)�y��nBWw}.���HoA&���,���ca���Lua|�8��Aa�|��:�����}����>@I� ���HD��WӒ���#���g��K/}��G�#�����$�"x���cavI�
7��c�O!)Y�-��>Rڣ����M����=�Ξ.�����Kf�5)���w8�2I�XZ���/HT��cƷ�c˶�8s�D:w߾iZ����'���F�3)�j7�OK5�߇�dLf��h�@4G7���O��O<��������wd1#3~����d��͠��]]�4:f[�+t����H�������X9c��9���1\�xQzo�:~���N���ґ� w��%\�t�>_Į�;�Ѓ�#E�u��ՙ�091!��PHQӕ��0w�:��}�v$�ۄH����ȸ����`j�Ɯ^���~ã�����^��9�j���1rzhG{
{n�[7o ���?*�{��'�?�˯�·�ǯ�7p���}��}Ѿj�L!�֢�pɠ�1=�ܳغu�� p�-BΞ?���y;v�p9qm��r�h+�b�<Yo��,r̍�N9�
����4��询��6�Qk4]�u��R�Hc�zg���2ʵ��'��b~�#��ev�56�'�l_
����T)���ǁ��ˠ2M����Z������V���oIʺ�k~�,����`�gF}��>�Q%�m�C��R�6�	��Zf�V�.i�>�Y`�2w��!�:B:��a�c��6��Um?�.���
ሔ"Y�Y�H"��	z��'`�%X��\w�HbT�Pt�.��|���u��0��tk#˻��S�F[X3�'�=��*�)���R �5�ӓ����Al߱�G��έ[	��47�Ç���=�N9&G�����3�� ȞTA��-���8�w���������Ŧ�Q�DC8|�,>�x��=�~����3�!�It1X�s��hK!�NUJ���L����*�/˙U�͸s�-���F�滺�Aow�Vp��5dE��b8��9�-ar���5��~��FZ�k!����T�M�\-��������g+���i���D��z��7 m�J��pm�N!ut�o�7P9GK[��<a�����a���q�.��0�R	����t�LS�����xh�90ކV�r�L�/�ɹ���=�<s�1/�,bj1#FRa����E����q�]h��т�"` X���2�8���5'L���d���A�"�\ך�P���wYn�Y3`AR�d�!�V|������̮��	�̉�6TR��	:�����4x�i%�Ri��Vd�U�L��l����h��ePujAPCJ}K甛�]}�O����*�� F��	0	c�((G��M#4Ma�y_� ����7p�ƀY+��Ǜ�ҵ�*3󾗆�)Q�f9�����L+?�W�ׇs<����aiS��=����� �u��Hp��Bʷ~5�k�V����Rj>X?���������Y�{�m��ș#�k����l�޵|��(݈�|��}R?���F�h��'D7�	��$�U`Ed_����IF߼{/^��/��o�G��ֻ�a5���0:�Q��l�;vR�o-�6<B`������lي��x+�Wp��Y���a�<}˫d̏��o�N%}��R��������^Ǚ�g���& C�t ���sgq��q���ܙ���\��w>�18<���%9z���O9{�o�
g�|۷m��������c��o>���<�Q�4R�v���	<��gH�0}}��s� ��p���f�p�ob�w�;DQ�_�_�e�XD�tZ{_/��Խ��g_�h!�+:t?��+r�y�!<��~i��5�)6<H��ri��88gqy��x����ß��e����a|�;�ɫ��Sw��$E�<�������z+���Sӈ�$�O/�opwܹ���n�8���u;�����b4ϯ~�ص����K�����nl�5*3��D7:�J���x�3�`�WjA9�x�������N\�µ+�$���'��<�_��6�����yo1c*S����y�Q�c�
�`����K���O�����_�
G�d}9�l���%#��,G/�\SH���8vߺ��̓Btp��E��u���ǽ�݃GPZH�.����G�ƱH�<���i���7���c��F�[?;���D�-�}�&���Q�'��}�8Ś�p������Nͱ4��I��`��_��؍�"�5ӫ��7#kԋ��jÚA��-�Л��	;�ܴtm:tGgǵ@���hf>?��#�D�\�!�R%ۺ�[�8^$���9�������CX�Z_����Gg��R�Y�@��5��F��d@t�^V�2ݖ��AU�7���:�,���lcr���濅O�r�>���T!��c2��B�=�y���^c�JOn��!���9$)H��q&���:I�p=2G�
�y�Y�=S� �{	4#PY��-[�O@��#����!�Zf��!c��g������;���H��"�5���ba�oށTG;�`�t�9��Y�Dq����l� OJ�	��s�*�+��w;R�$�;�p��d�o���w˸���4�}���g��|�>	�dredI���h۷�%Ս2�{!���<����d��VJ�4��eխ�VjIOT��%v[E�zI�� G�R�aU�.�
�d8C8����L+��~��*�?G����`)C`�@�Na�7��}�޺c���7$���_�L�I2*Z�"��jH_��pKk��Y��`1��Bǖ�~����)>�d8Q�?M��	uǤ��E?U��(�S����A/T�*���(�<Y\T�M�lՐ54���7(���7�=����d~�Fċ�I5r?�[1iU���>�Z	S��6Ƶ���������KeI�
j�a�S���Ћ��D+��ĵ7Z�.��Cܢ��r��u�0�4�����8bB������U��v."��}����j��/���U���g�Y�~v/~�@�wǯ�������zfY�a�l9��$��F;�:��f�����Xc �Ǥ�s~Ϸ�H$j���Rk�[}��~��	J/�1�]C�Ձ�k~8�՚V��a~���֞�m�2ǵ��j���Wf�rl����^�U�{��/�-�<9<;��:`��M���e��B�#feX�8v�4��t~㋟��q3���3�c��߿�:6�o�s�vane�@G7�x��9s�[a�;i�������1��\�M:��$��Ӓvǅ��K���~� �$&���yY����'UJ<�bH��V��{;xp/^����~��Ǆ����@"E#�v��/~Q�4><�K!��q�itX̗
�Gv߼�tG	o�����>��a�Z|������<�y��x����<z	�/�cr?@�;����e3�j1���=p���S�aN�<�{�[�T*e��C{p�����/���% �kً��AK��W����O�c�N��ܳ���øx����8{�,BSx���������?#�&N��Kj1#�t�ڹ��K���!�y�}�)��ɻe�[�������o�&�~�I��a��x�B���JJ�R�}��������Ͽ��?�~�?�g<L��W��7�������D�R�V٬��Cel4$�;�i�6\����?�#�ڱ��[�[����E|u|ݝ(3�?T�&�Ռ�W064����{a�<֋���_�c$xKa5��S�q������ ����O�HŒ���sU%��U�f[�Fs*�d�V7F��9j�]�h��
�d���n�/������W(Ͽ�����,�nM�{&�h�=�7�)eN+Ѣ�>��5{f��ɹ(JE�L����g��50�>�)���Q���n����I
ZF�{,�5z����^[א�u?<��i����"O��aU�֢��P/������QJ�V�j��\��vO��p ��4�ZO���
4x,�ڎ�XT@�P'o�6ǲt�X4L�8
h��8*����%@s���<�� x���FU]\b����S�V����.q����[q��{��dIG-c��42���7�1̝8q���T{+��q߽��񊘙���}r�S'�UM��~V���{���=yێm���[�f���pm�
ɱVa�֭XXY���X^R(�t�rw
�H����;���kҀ��M$���rW�{g�B:s5��ё^I�?uzB�st�ᡔ�R��V09}���{��0�i���ϥi�ƫ!��19�okZ^��\o�2�Mų��{e��^"�X��bn� �hXİͬ�����*��C@�쌞d�Ѹ��Sh'��6҅��	�7f��_"݆	F&��۵A�䘐�#��e6��`J�h"NF�*t!�x2�0�0�S��X�^-�r�q��-{rJ�چҌ��@Zx� c���h��1lnr�NY՜�5A߳�|HH���o7_�ڨ�M↴�(+y�]U�(lGj/y�B���48M^w�'6 �~��у���?���jPW5}���M"[����M���N�;��Տ_ ��ץ\�'���d�#5�^֧�y`���b�rL�ʩQN�5Me��515	ވ�?<���?�'���-��&�z��Q�_��=a �Q��TEa�>T��F�0����n<Z���x`p1���c�aX����r�ƌ~6N�J�]'�8std���W`5�r=k#�p��!lqB`�a�u�Hd�ϣ{C)�V��l���62a�})�M�����o�׊=�}N� r�w�GR�%,%R.���%�K�}�Z���qO�~X�(]���'���~�eL��������6vߺ_����ϼ𬀫#'N����1�݋���=��B�BJ������іV����o���s�ſ�v߱�<p ��q�[[���ROx�&[$�*��������������Q����? څ��毥|�K_������>:t	L�]����Ӌ�y�ٓ���o�)F�0�J��5�&���A,҂��ܴǏ�Z:+T�ein�F+܋���)��?���Ԙp+��g��k����k��"��;q��)�'��{N� []^A�g@���i?L\��`5���L(���#'q��א��$`4���?F��C����J�̚Ծ0p�ƢRW�����K�$Cg��O��1" ���+�O��?`��-������ēO����R����4Ì��<�2��J ��L���1����������k��'?~�TmHzDr�R�VuyL5�[�He���;��A�Әn���o݂?:�����������Oؽ�6\��J�9�K�����l~p�C�y���ԍ����9��'���ь�,�"C['��4���TV2�%k
�(���"�!�ݯ�V��1%n�*��3 �Њ�@�_~x �d�(g����.i�'�>�4
���@�h2b�ϝh�g�p�F�@�g�������L)�>ߧ��S� ��дj�����
���� j�W�Q�"��^���cH��/2Z��e�d��!ױY�/��]C�ӌuP���DO���l�u�F M������
o�x��0�*��Z��y�D�:�oi�3P�d���d�e��l K�[X�Y��t��b�@_��e#�Xv��l^���$�,p��1\�x�}	�������&�2�P��B6u��S�z"c|�ft����%�����c9�������s�Eܠc�Dn\��C�zIO�$%j���q���	��E�V�XɮIy���nL\D".nĵ�Ki�8vV�,�jr��rv��׼6��B������C�y��sA6�A�PI�q���X\��#�V�c@3��N|��W�V�P��ݛ�R�g�-����G�s�kc:�ln<���8c�	/����b3Q����F{;�m��	$�H�;E��8��{&o\ǫ!�\A�%E�fMz2�Cq�Ln�jF�xeI5)i�Ǔa�5f�����6Is�x��BRt�@�&�_��)�u���M(��W��6|ͽ)w	���:�j�P������w���~��Ȕ7�t�GϮxF)�SpN8�������ȕ}�a����}��A`&M��{*j����t?U{��~Z�r�1�MjfӇǐ�,O��j���\`}M�G&�>�`�O��`��s�F�*����|��솘|cp�/6{4��Zٗ��)��,��:z���8�&$	ͻЮ��`�?o�� ��Z��<����F���w�ep�1U;����9�y�e�t����c�F�����7Fn������2� �mI�mM����l���s�;3���ф�����
)�����}�JY����u��g �eb�<��',�m��q��30�<�U!����:��Bخ"Wʠ��h�HGF�0=1A��o���Eē�Ҝ�ȩ�d�.-�#]� �ъ|ږ����K0J
:75�b.�P$��T�̃�:0�iMu�rk��²g��ū��Ƣ!��N8������J>��r�tFB�B��4�A�>�?0���� �V����w�~WHR��m8!PX��ʬ�z�r-\����&p���q;3\ކ�~�>>�1�h~�o/��c#��������>�W1�+�hKF�4�+W����C�bf2�1s��N�ݹ��A��vI;%nyd1�_[�$�R	a�֛p�}����ҥK�L�12���114<���oF�����~��Z �:0P���ނ�SS���_��W��C,'��j�n�C��Fʼ��wރ���d��08���g�t6������	�E��/>��^Z�Lё�#��C�+��;vIm�jf�
�i_t#N�r�Ʋ���;������Hݩ	`a��B�<���|�����\������������g?�(���?��i���;R3�̳���M���_��_�����i��$CH���;�1>r�_��l����wy� ��xf��a�8ql)cW���ad�-`h4ry=˰>�"�&�2���U�崳�g�y�-Q-�����wŜ�Ql�ڤ�� ��e��k&��b�8Z�K�я�������>@giW�O6��7ru���IjS&����c�: �T㲗��_�ze4\bP�wo��j�M����k�zo�04��sPh���z�qj��=Z��q%�
����f�<7�?U��m����p�\vuV�ö1@���	�Լ&ǯJ��U�L_;+��5��rIZ�XvD�v��b�d0����"�|>')����W��-d�ϮJ	V�t`�d!��r�;��`�&=Ƚ��Q�|3kX�>%@�"}�E$��H1�H2N�[l�p�����i,�LI�I�Q)����ce3s�<�D��!Z���~��5*��Ԭ����ʁA��i {%P`fKZ�-�l�R_�@0v���ӄ�%�!�`:k�{�K����r��qAK�`H���&�o� �Gg2����H	��u�+Ȕ�[�����w���g��f��B]А#-8�Ņ���{+��9��d#�
e��@'��9.�p�����D�a6�]��B$-|8���祥K����mA�{j(!�7j���h�1����Ư�np)�B.�+�X@s1'�����~����wS���n�gcZ7~�P0�?�fV�5�����q*-�d��<�j����m"#F�Փ�غ�Y�g��L�#�oƣ��킖_�j=���0�wy_�4�w��>N����;�ﮇ��I?�<e_1�]��JԤ"�vs�� }��jF�i�⟿��h�6����&�l�wj.�I�24��ƔN�b/X8��O�^+f2��l��{Pn�
�&������	U�,�S�P`ҽ7��*�W��X>᭥�
�|�]_o��o���q*�RV �5S� 7����HfG�	]7��������w���g���bW����c;Pp"Hv�!��A "�kW'�[M�/��?��T��˕?���۰��0�e3�;ѷe;r��Ϟ�@��qO��m���ϸ�Ju�Jۂ�-;���	�����p��ydsE����^�pqB��{���F<JF�s��}�>�7�|G��s�=���އ���N�������R��I �����N	��g����C���3O!�-�W�����6�O�M�%p��í����053/���;LN\�&���$F�c����J:���E�o�t��:���v�N����,�/���)��7m����G�欗ѱq��20�8x�"���j����}��Y���&,/.��ߓ����fw��i�<��������O�5-���>�?��*�tv�!��(�Jש�S�?�T� �����H���C�č�y�m�t�]���~}!��h����x�w���M��'?<z�ϝ��	tww�ݷ`�������G���?��O	�͊s���ߑ��?}��<=�;��C__���,-����\������{�Y-���^�� {ӵ}`�E���9/�k��Էy�4���Cd���(�e��	������t$��j���G�HW7����7?��І���yn��ζ�:�Q6�'wjO�2�\�eҞ�Tr��<�sj�ޔ�pE�/����H��e�N^;?} �.��=%���3q5'��oZ��@����#������f��~5eBn��mŤ��S*ykfyc3��v�f�~�+N��ϙh��Pa��,��[&z�ng眥_�C��`���F䎏A��7u�y5��=��Sl��L���N�V����+��0�aB|�(}	�������P*�ݲ2�_��#�Bw�S�P;(��%P _�R[�Q��3X�:K&��6XqK!K��`vM�}��a vTVXU�u��1���o�1���¢	�]�뢃��_�Γ@Bn/��<f�I���~�vd{Aq���f"���>�K�w3m�,E�����W���~���5a�q�$�G1��O�Q�*��_a�DJ��J    IEND�B`�PK   �i;YF��-$  ($  /   images/d88a5b0e-66b3-4edb-b452-47f46dd40326.png($�ۉPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  #�IDATx��}y���/+�ξ�o��[-��I�,�as�k�k{b����Ĭ���X�ځ=�����zc<�'^cds�!�!	��VK�-�}TwuY���<��ZjI�T���̪���z�|��}��p�����>on���,?�aW���Gy瓜{��گg��ש}�w����7@�tvT��2 ]��|j룰dO�f�>�}[)uP)�{���B����ත����0ۂ���G"�[�UEoUѡ
:#N���@l��Ӵ?�(��d6��F"t�"W�� ��b�rR���.(@޼~��`BS��i��b-'N�$�^G���L�&�m#���X�%O;��e��"�>��$<��v']g��/9��ou���	S��;/��!~ d*0I42q�C1q�b)��Jb�:%&�2�J�#=�N )q�Ɖ���]H��U�Oeo}s�����؂�8�ca$2!�>tp� ��.6l�`d��i�,��b��L���dSv%���ޭ�<�[�ʲ��߲JBj
A����c���cy��<����f\C�`MC$&�SI�B�{M�W����}�o*�Q;�й\������u.\�3��f΀V�1?����rȆM>������� �K"��f�⿧8t�R�<[:��ZjtN�H�'�P�N�0�C(�A/��M�6u`�z<'��.jF��R�4R{��8"P���F*�h��R��w�]\G7AO+���rC$�r��;�)��� �q����wl 9���iʠ����0��ފޗ�";���N߃��/C��Q�(�-y/�N=��ڊ��6$��3�f�C_K5�,E��-��Ș�5I���������9C�5���
����)ddK��@(.0����bٗ��Cli=�<�i�������М�pB�B0��;g,��`dd���+uZE��Ɇ���/�=�܃E�!�a6��+���v�F�2�B� #�����l{�3�$�1嘪�H�QT��	WR�@���b��4h�-�|~�, c�0ad0��1Z�@J�Ĥ���0���*!�?���� d�-alղfԮhE�D���C�X\�ٜ0J*���͛��s�!�N��c�Nk�o��F|�K_B�|yfh>��v���}��R�����8Z?N�������]�1����%Ʒ�ёhFk��^W�� �B��r���e�H��5h�$���z�C����L��.�1��O����l`X���9��Ha�PV�ԡ"������J�q�X�|9�|�I������S�r�J|�+_��^t,
A�4y
���0=��a�X��oB*�'a3�t��4P�����XVَ%��D�S#"):�`��I��҇�e� ���J�W��0�8�@�����V"g�W�ƞ�c�=މ��0g���
��3����2X�]�yÕ����y���_��9o�<|�k_�O<����3$�s��8�&����Aqm��݋��QX��.���o܌�<�l���0�e��Oh�ê�K�&�X$��ּ���3�"1�\��LW����A	a�z�P���0�H(���z,�h�����L���Ǯ�Q��aE�*���8�2LDt���>�0�g����P�!444�z���6�7�,,��ߎ_��gȲe����^tQ����_��ub��M�/@�|Ri����`�s-@�D�$���~	��,����#U�0\�pU�H@��[]�� ��baK����*��h�8�f,�h�p�������J��a��}}"�?84g#������O�{<����a�?~����k��/��&&&�Fz�t�k��@����������x�w;j��9�(dl��>�6 �>3����+��v�HG��E_~��H! F�Ĝ�J��n$�¶> aEP�!��v2�`��h�J���wJ�(dD�B����1�t���+�������7����G��v�څC����ڵk=PX}%�I�T���wf�TWW�pVSo�����"��/~��5�nˡm�'ȵ-@0L�=u�`&�^]��hX�d�R~(��,�s���$!�խ�
�3�S���H�-3�� j �WJ@��Q�φ�*�(�l�W%����-�:v@���p
�<��	��_�Ǟ��z6��<ۍ�����7�)��}�Y���<�0����3�<#^ß|�OP���I^��y@��yCGC��5]������dq��h��9�
ny� ���X.(��*O	=�+�5�A0lU�����4r���*ɵ�Ӷ۰���3�o���s�{̠u�i*.{�������-ro�\��c����sp�+=#@�����Ν;1<<�U�yU��8�0����v�G�0�"0\�}y�"|�i�0�??�4��'0E�x�Q��#n�0��3�;��WB�I�FĴ��[1$O[�uqUǥU�yh���%6�>�cAàW��Gn�B�����<����cŊ�<�3d*�7Ŵ���6��a�Z�9W2�@ gmf��WaUr!�I=�D:X%�De�gC�*��|=9�E฀ؒ� ��{�dDD:t�W�ለ-㇤R��+m�`���7���d�\P�.���M0���w�?�B̆f�A_444$�s�Z�䟮��gUe���w����-ע�\���� �f0� J^�q���\Ȏl�-g�*͕���+�tn1+,@��QS}o����VH���/�'Ɵ�.�.����$��,N<�'N�Άf�}2��5���[��E� �i8@����^ppw��� �m�8��D�i�t��������F��)��OM��CgUE@��߆�ߪ�[9�������v���� ��:���C"�\N���Ff0=cw�T� ����~)���<
8�������L��x����'s��dLP�5A�-�XE��.�(�NݿxyF��P�,4�j2\��u܃�s��<9]�iX�������N���K���+�_���Ӌ��-ۀ��z�=�Z�[�RHQ�́���
�D̆l`���U%�����T�׫�*��w�GǞ�Q a���M�����~ؐ��贀�t��u�U��� ��au�6���;Z�̏a���ƀ0X��'q�3���4ޚ�tx�n����I�λOvn�	�
v	GZ�wL�汫uk����销0��k���4J�e�)�Nus
��s���'?}D���p��B#H,%�az�S���T�P��fP�w;���g�!L��`wJ:=�Ćͣh�cA:y��90�+f��k��3�@�QW+�pK�:D԰dL���'Ĉ�b&b5�^�Lh����)��H���[D}��80epD�jߠ��1�p�)�dF@�wmO���Y���p�aUuC�*��jě�S!@X�ݛ�(��խ�S9=KL�p�3��������o@���$}?�OG�5��{gd 1���r����{���K��I:a�����^�ǍX-�������I$;`��Oԯ�k��A��÷'�%>ܘ�Puι��thF@N�PPE���
V[qԺ�~�H����Xe��hy���d����M�s�-7�s�O�@q���5~�B�����`*	H�MKP������n�*k]�R�J�s����V�E93G2ܤ�jؠ4�kpϜk��]/�t��K��J���������= <�u�c���~�?�����X��K4an�A\���<P@�}/��ڙeڎ)i�o=�]�������t,z�l:h6r)V�3� p_B�ĕ߹��]GQ���~�ignY,W&/!�v��k�/&b���?���%CR���Y��tv5_��n��X��n�Q0P�����w]G ��M�������"Z�/Y2���p�y��%��jQ�����XSx���%C2ʦ�Q�TQ{������N�Ԑ��آ��!����}������0^��om@b2'�bZt-��b��C�6N�Z1�c�Q�3>�Ĥk34�����t~�q箆����>v@��cM��n%0���v#��
 �R�Ib��@y�1�:=���(fR"��E���g���n�F�{fM�Z��^��Fv�"E��
���3z�=�u�[yK6K�G�!���n����l�l&7%��b�%6��k��*��"NcЮ�[�w��;���'%��|F	)���S���]˲�.��M��ڽ�q�'P'��K��dGܱer(�0=bp���awK�"%<�rab.���U�SAi�<}|#�V�`�4���>k���=��rs�n�U�t2%ŒG֑[]�wh�îH.�މ�"%��(,WF,|����y/��������@Ϙ�{�"��0��e0J���H_2���&/�l�A�,1�'tM�3q�PH�"��5>@�b�iY�f0g���$t��q
r���w��/[�Շ��(ъm�q�C߸{jk]�M�y*��52u[�t�2�����!�2�̲%$�-6˫:	׽�Y�U��v��r�<��k]C�\pF��1�h�S�H�3����Ɇ���<�I���$�rVY��V$	����<n0�#Gx��L�,�i�`9�@�}�}VcI�!ܑՕ���&��d����I�%D�i��n�9E�R�fG���c; ܑ���T}{���>?��H��w	���"�0P߰��rg��ivda���-�sj�v����r6���i�Aol��Z���*�8�a��r@��G>6E������9R��&@��A�p�?��0E�e<Ό$��p��w�Wk2 �՚�a10�`��,!��l'���g��9sr�(8�܉G,5q5"�VV�;\l�ن4��9,φDH]��P�� �R��?-ϝa̳ȸ�����V��k���~�7�D��}�Ό��?�����߸�IX���VY	ob��gze��Rr`D�NC�����͏4�Z<�> �g�%Xe���`f���#�ʈ�)�c���&��ޔ�}Γ�z�j9�3-��pY4΍�y�E��ס�t��^RgVh�Q/G��F. ţ��Y똚��"����v��t��	.j�,.��%`)���p�p���ʲ�u�dyF�'[Q�}'J�ޥ�5!j\Qrc�K��v�����	�REj���i��H����G�eX΍���݁�3�/�T�:�r~�,�7��R���e��ȭ0��B7W���ኢx.o �n�^V���� ��<��Xٖ��p�p�$��e,�]^#�l�k���P ��UR�I�����(ә�W�v���6�$#���Cp�� QvS3	1A�/�
�rtfs9X?�+��Eq���rE��l���ha5|���6]�Nˎ�,����%C^�M���#;�E_uҫ�ڋ�}���[�~�>$�x�'�dGr���e��®�ŵU҅�r#8J��S;01��ծ��?1��!��PQ':���Dٰ�!KѺ���ftge^M�)�f���ߒ�'�*��{m
��o��Z���a�T5�L�'~��^9(��#Wx8ȳ��!��P[���C~5F1�E�h�6BRR[T팣��Q�
����Rrz�G��%�bi�x���t����i}�`���:5���w����q3�x{h
 r}G2)4U֗��,���I)Zg&5��؝�׮��%t�6����4�;Z��V�g#2u 'R�H�NO�ީ��H��N��WYv@�lH
�������>�p�ŨI�~q$H ;�&IIDbe)9�x�@QMaµ�Lt�e�=�p�@�^�h9sF��^�n��_p`���!Q�rL�|>XA�O*t�����q��R	�D"�T����w��JB�K��PW/����q��W|Ǟ��y���:����p��rQ�1�p�X/:�sexPYJJ�7������T�{o젷�� �����d�a@X�"Z�,��_���5��`N�OG*���;����RR����#'#΅xI��1���C��r8�2�@�� ��+�����<��U=���2���$E�EA	}���	�V7�#�Ĭb0�f�+.�̩�wG�I<�����pq�PH�A׀u��ֈ�*zy?�>����u㪦U�6����waE�b��#�DX��I���g���!��x�����*�����o{���-w���������Mc�
�߆�T`�<Vt��R�ވ�D�<2�!�H��C�V)9+��&	���j*:����ޑ'���Tr���P{C�CRk1Hُ}Gpe�j�{���$.l78���{^���HGXCj_/�~��?>�'w: t
/9�xo�m���(��06����X�Dn�E��g��@$��iU�:�]�~�(��I�izz��>ˊr����[lRާ��D鷺ؖ�ƫ�\U/�.FbV�7�s>�f����,cׅW<��`��ƹc�QpP.0ˊrL8�5���G0n��LYg�.�;(E*"�Ҟp?׹�V���l��m5.�9@H9������kv�W�������*���V�u)6ѳ�qr�h[	�'�_d�0מ���u�*Ĕ^�}GJ��v��Kwb���Zԥ��\r�urn7dcgE7v*��O�/������|��|��o��~��je��<����c�
�R�X�W#|j�������&����G1l�c�r�dO�RإjXټ�c
�6� 6�l3X:~?��&�K��E�ƌbݱᥥ� L<�Ū��7T���<�X��Y(=�'�˚�89��!; �PK`4Fj�-C{�s����;��dQ��s�I�\�]1���-�Z����~� phxpW�,aSB�9!y.���2?F��/ḋ�Ԝh��<��%c���T�Y�ʗ���F������bs
�>1�b��4�]x�C�R�R	���J$	����:V�,�������"��z	7�>�O�ْ��J�!���?oA�Ϸc�ųV��E�[����0�a�����;];��@���H!��*�.,�
���%sۻ�[��]�+��D'���xE�Q������f�^�~�֭�?����f��t.�-];��qړ-�~�T��6���;5��FI #䃡:j�������~~�yw���4s`� g}/��rlܸQL�U�n�m�oh.
ݠa�����\a`8���H������7v%Li3���������U����;gޝ�`A��͙37�|3��y�MN:��> C_t[W�,<r��o�#�,j�@[��p�Զ���x}��F��ؖ�'�llOJ���z`�:
��������/��b�1�k���^:(%�(�wމcǎ�Z�B��?:�Ј����)�l����C�rb��硱�N~��d���Y*x���C�0�O���P����@�v�0lKˑ����E���$�g�%�E�g�9p�@��Č*����C�g?�6o����G��fa�	̸b/�7�i͌a[�.�'j�����I�E6�5�d��uHx=�#c=΍�=ˊ����+q��a�������w��W��_����UW��===3��Lx5�Ç˪�.�|a։_��W�~�zlڴ	������o��1�@��+p<:�ɰ��-����C�aj#Hƫі����zĴ�S�����Z���¸>)����,�7��W��oƉ��,�}�7�ݐ����ר߶m��I���O?��~�e׶�Y��W��������b�вQ�=�W��1I?N�����p��ch��Ese�T%*��.�� r���J�\��A��g�>3��efs��UG�**$�E*�=jq+����3`��I�G^��W���{�`����jۧ�S��,!?��Op���˗���ª�*�	&9F�������W��^�G�i�r
`xe��ѓ�zeKN�05�*�Ǫ#�����a
�(�s�ŒM��Wd�,���[F�᪶j
M5؎�
q�c���yM=�h��g-��F�R��~YY" $}}}��������i������ǽ�ދ�˗#��ʧ^�����F������'7�t:���ڥ)�>��+@������K�;\j0A���iG� �t�	f�((�V�+8�3�lb��Z����.��9��lB@-y��h�0*��$��/��N^b���A�S�b����oK���m��fvww��'��m޼y"-�!^OZ:ɠfm7�EZ�c"=w���ʔg�����fn<����������?�U��^���x��=Ԁ+������.�6� ���=Ś��.E{����Jr�/u2�@ngE/�x���_X���[������d����3p`�l.�ܐ�@_u0�'�E�W'��5M�=��l#x���")��.Y�;{d�=b�b�0^ӂ��s��zժU��v��I�r*L���6���QV�e��Q(��7P��&_��&D9sp<�+S@��P�}E�_WeØ;��5���5X��VX�1��k�=:00�36g��=��r�#S���2z�\�qÆx���H\�zL�
GM\�A_2���8Y�FZɋ�/�2}��ſF������VU	�<$�k����?����9��ʍ���S�ܷ�����{F��݋�I��!gCw�u{�O��L���'�>�@:n�|�ʾ�n���^Gx�1կP�כb�Qϣ
�o�l0��C�dy�	�֦�h�n4�xV�������u�[R�(��y�Gp>�2b�h8]����孧���TkSs|4�ZL��% �Q[APt���=
˗�q f��	��+J'�M�mz[��V�ns���A0CF&�C$H���7� K!�k�b����O�'�qi�%dk�&����S�8 HP;�!���c�" �	�~-��Gҕ�����q��Fs�Y,p�G�&V1R�]�=|��Ge@7�☗l�D>�&�H�`�sK��� /v�W�^�0�� �}��*�q���$H/�������G� ��[w�������B����l �(�G�������&��@�b�    IEND�B`�PK   �i;Y�H�izN  �g  /   images/e9a9c672-7031-4851-9c94-029b4a1edcac.png�y8���<IJD�Tv=��%�Ĕ%���JvBD��3T�RTDdkAkֱ� �l�m�X�l#acx�����������q|��:������s^s���ޖ�{7�P�-g�蘠Pz��6q�+�O����pzi���	�nr���<c�B�V�����v�\��{���㪷��-'�����5w7/{O'y�[ίh'��P⨳:�.�'LPî�⺦G.���ۋk��:�`���zr�K|����T�<��:<���zU%{W�.�K�F�P��t�ݙ*	�I!�K�[/G��0ؑ0�-#����H���'c,ےAII�a���S4FH���X��[�؄�������������������U�n��� ��؛�++M���Ә"��x�}��ݡ�&��Wә���q���%�l<��TT�P����sk�7�W���xt1�W���x�h���\�%�nxs����#e+��!m���r��$�� &��~�2ּ=@B��kq���5��w��R�� \�]+~g�T��J��Du?Zi,_<k�6p�\�׈��>�P�cT0)S9��Mc�#ɹX�m�?��]�eD��P��j�J��?7�+ˌ�ς���LR�u8?���)10᭲�3W{	����-jﱨ�Ti|�����������~�����$����;��Q�p�:諳w��^�h�x������]������F���j����(������'�f�|�u�~������<�MՉ~[��k?�����bf.٥]&�g�?�9":(ᶺn�N?;���!�Ӣ�vۻ���xU�5��	��gj��ZU�w�$�+ǜ�-+A�r�h�V��9�U!HZ�ޓ�1G�8��pl�~}�c���x���x?���:$!��-�{�J@�]���]L-��p���#�� �t2x+���M�w�̻B٨~�n�)�ӯ_+��3�� ��'�ors�����p'��M���|�	Ydc���h��)�4Cf}r�Uśh'wv�!��[Mؗ�c��(����_-�R�-��zdwۤ�D^�O�m�����1��,+�	^w�M��̿A7��b�BN��m�+`��wMd���IL��q���8Y	��o������cYX���-�U6�¹�ˋԠ����o���`�~�X��Te%�0�L�z!��l)p��D��W �V �_�>&.����/O����C'7�	���9�����z�����o�ݟ��Ba�o/ݝ�ť7$}�2(�b�UωW��ʶ,��\r�t@yzz<v1:K�w~�97ց�������]Y$�U?�t�����zQ�(�1q-O�G�_��roֱ��(�������sVC�q���<��ఛ�q�:�xdK�ޯ�[]��f�9��Y]O���k�x��'�K�{zZcۈ
���=��'���O��/쿋�1()�d�)M�z������c���L�<wS�����?o�O��N{�D1�1�(f�M���� !���|z��2I���#}�m��1�${����x����� ��lpە��o)h����5@<��S'r�	fQ��+��p�T��X��l���qC�/7O,�U
 ���a���{�_�e50�o)�IנV�X���¨-�ѡ�z�ꅒЕ��K���a���M �O����_��[�
�r���v�I�{ʹP�ն*�ͦ>:IvN��r�9p2����J�� �1�5[Ŗ���9���{3�IE�M^?�,�� mB����k����?Sb{�`,7�Fj�&�[�P�� |3�D�ؓ���>ܴ�/�_pw���T�y��Y5g.S��5˨U���xgP�w�c�R/�W�����KN|�c���nW�|�q��DXQ���,,gp�&�оxS} z�>c�����tź���I�G}^ '��%�yϭ�m�
4�}c�5`?^�6J�tR_p?Q���\�*���xhr������t?� ֔��"�,b�S���z��D��A�[���7��ƕ���מ�fM�X�"�]�@��9�
� Pܹ̩{n���� Jy�9��9������1	-dD�5��X��JZ�m�FÓn����n)�دR�H�[Ҿ�f�v��2��|�4��h��y?Q"���Fv�:;�.��D���BI����K�"�"�Nn��< �����D��G��%<�c@�?b��AD�ےT��Z��G�'�����,�����6��CN�������>j�}O��P`P-vx�E� ;M)R��aP. �s�����o��T{�Ұ�{a10��f���XH. J��¾n�;��!��Y�B�����J��7����]c�J��$���$����%���ݕ֏ ��~�������)e��uX>����q��Z m=mm]�\���_��}���{WE�'�S��Gq�#�j59����؉�h���_�� n�+��K�ߝ����ooo��=	��~� ',��4��E`����/3�UeY�累�
��o;�gk�@`��ץ�XDQ$�e�v�N�Bq�Tr��~�a&�x�^9c��ܧ�E���9�:)�IB�a�<�j���	��­#I5�:H$hF�Tk�r��{����~�`>����7�g������3���aϛqC��#�T���Y�G6U��m۾D����"V�=�:X�bd��U���!N����m�|6h�]�>��� ��l�À	{29�{�C��������+*���q��^��V�r�oY2^0�\�����,��tL4`�q�$��O�n���K��۶)���J��n�x�[�+�|�S���%n�7��~p����5�i-�%��}�``�ns�Y�e��f��?�a\nm?� ��7pΑ�Y@���lAhU;9�6���(eEݖf�'�~��{����8���ԁ�����D�z���q-+�4�z�d����D�_�1n�{j?�*����^u�HS�c�y�U;� p�4;[���A�-Ue�Am�oz�>��ɲ���i=�����~ў�a�\���Ts��D����%N #�D��l	�I�Pn�5\|�^�~�h�5��)�����hn���y=�ߧ�,���'�#z����JŇ��̀By��b]�y��[�+�uS�6׺˱���mM�V�����"DK�Դ�bؼ)�ݦ�q5��"��R���k�>��܄��Ǘ������z��S���N�l\?�
,\O�+�,B���@��'==d�������~���w��@����l���Ϟ��H�J(fv{�� �Kܒ����p��1I��Ju_�Ԍ��~�t:��3p���!�*w��Q׍g�	\v5���E��b�?��S�x4��! �I#T�?��v��=�i$��q`���N}��߿�f�Y��
l���yq$fi~�����\�s ���V�YLE�װDa����K�ȡ5WH25�b�+����iJ׎�;L�sEƮ�6�ҋY�_7%h�"`a�1�-IƨNl��Ɛ�c�1���'_u\��(�'�:q��M��?�=���R&�H�(D�/�(�^ア��������6�	�w���ig����[���Z_���m87#�0ęg�S N;�m(9�n
���K9D1��]�]D�#^2,�[rT I�]�;n[��[ӏ�qX��-i;-�����x>�ex�|£R�_�
Op��pG�aI���-Y�)��BM�I�zg�ch��Fc�� �S��`�x�!�CZ'B0�`Et����S�7���1���T���Ľ�#�1����Wz̩����c㎝��� �Buvt�`�oZ*;�Y�#J��g�!��
seZ���HͨP�����xgH
���:1R�6�uט>!��	\�w�F��ݒ���0z壆��*��.����4`��R"�iE��f�vr׉{��M&��j�E�Ӷ*��~��М���`�Y)����������I ��	��f�`�qd ��@�O������P�� �:K�Fn�+�Oa�s�w���]M�%m��!&�� g�q3b %^��~ᴭ���W���@\��Bj?��̪�n�+��l�=����;��i���9�	����F9?e�>t�S�+O�b�glK���'�T����@�����c��4�K���ւb�u�C��!��n$i���6��?��n�F����_�R|@�T`EwJ�l^m�Zg�1�,�ƭu����Iޜ�L1�v���Ƙ����eA5!5X�D`���K'���_y|�@�Iծ&�?дKH���v��e[��4P�#M�G&R60JJ���+�n��;�t�Yo�h8���b��n�B�������� Uf�x�- ��am�O�?��>��J���(�o�3,�?���X#�;��p������U����&���Ϲ�!���F�5�h�.��s�S�T��3���WNT���#�D�x�sG�@�;�iTH��}.����M�@��Q
�m�Շ��(����q��5CWWU.5��} �G�s�>l�MaA,hC��N����,�&�U4J�a�@���xh^E;@�Ҷ��'�5�˭�Fs�m�!�n9����㳳w�U�Y9 �&ߐ�TcA|vOt�T��hw��a5r�"��6�u�>0MkV0Oi��?/G�.�o=�ݖ��5�X��ۃ����|��$��P�U�h2ғjc����F	�5䜇�o���L5V�m�w1{�*���?|�V�a�+?W�y;�8�uĳNV�VS`d�8vs�X��R� m�	�n��)`e��Pܚ`��_4��.o>����_���jP�B,�MN)=0�lU�԰xԓ�c����gp{p*`zP����Nn7�S���6���
?�0_���Qj#ս����4����y=���qο��Q������ǌ�L�+E��`���f���}�uD��$���N�^�:�TQ$(��w���ع�Say�{R�7k��]5�S���_�;�,;+Jm�b�vȩxW�����#�2Dǂ�ӳ�wZ숴�$o^3Z%(��E�[�Vo�x�� �!vFk	4O�k�*j@ʩR�����I��)/�;SJ
��<e��=5�=�4�W��s±NO�c�&��>Y� ��s���<�{\nчK�/�,��HBm����fz���'��m���_L�5v�xP���y�}���k�h����5[lt��f3�y�m������[��?�������T�p"�)Sݗޏ ]�PXL��{0�UeTox������~Im����W�������6�&&F����Z$|K�q�h������VwW&+J f|@�k���Ho���`��KM�1a-P�N��w�=J�Ǵ����e}	���}��5�k[ ���}4~���=�����~V�U��2"MA9�ʐ��]0y)4�!k�	(���r����fU7?*�`��㨦S�cc�ӳ���z�?���*�ZM2���q|��IE�uA!��:�o&�}�:��v})���ʮ��1H�u��R�1��{Sz�XN�p�V���^z*���
�U{7���x�&�d��I���6Q#�� �y���{��*���)�.r��Q(h�h�LN��u�6���h顤��tI:4vdh�Յ�j�������5�>�U�^uy�F��gڪ�91�:ø��l����;�]�W>�{@��U�d�z0��o~�X��f�`��sz-J��:c˜ۇ5�h��7���;�H�S�i8����7u�����x���o"[�#�+��r=�;��v��7���e�J������֝����iq(Ӯ����id%(�S0DY��T����gl�3y����eS��֌7l��CDK�͊��@� ��J'�)�z6?Զ�|�O}Z�S���r&�f�bP�n�x9w��y���p
��� �b�~�d��0}{�!�~s0(�ExJ��%f�JRa��px���&�p;�����ϝ6�ٵ��[��ٟ'cp���$'=Nxp�*AZ,)�56
g�o�(�@����+�Ƃ�]Ml_���T�)�W����e@�D�f�����E���I-���]ޯiV|�T5�a�%�l�T0���'����*!�P�@%|������:j��N>v,�Gɉ
T�ݵ���!n�͐�kԋ*��w�=�p��B�		��F6������h8�?�:�R�*ٌH��6}7�����w�"��4[�t��y�:�у`�k�5Z��bU{�w@Fas��+R��eȼyN�L|4/'�?�]���/����arB���+ L*�����la���62L���C8���MX����G#�]���Fn���QY>��E���N�x6Yg�i����Y�
��[g�dRD؊���n�m��}&�(��̼5R�-��e���qC_��O�;�l��l�4�)e;s+��;���
�����<̣P�6�0�~~�X�aX��)�O+q�����lOV��䩍��e�s�>�F���f�hk?բ��1}�����X�/�y� �%�����H��䕥�J1�ʕa�z� ����p��ԡ�����g���m��k{K��T���7jʽ{��*&�g~�l���(�x�X��h���aa?cm#��n�O�=7?�4_b���@G��Xѐ$��>V�W���H4����m�gOO$%�����,�w[��h��8ih T,B!p����-���wb�{$n֏�[:�uSx��r�<G�I	 M�s�FW+��A�� �]��*�͞J�;q�Ll���P+�^���$�) �_�93�4�� 2���h�ɏ���s��~�jy�~wM<G"�^��Q7úm��>���XG�����_�5g�6��O�����,9hy����X�м�䠱��%r��ljx?";�u#�;5��xY\G/O���0�u_�t4kt�N:��G�g�����J�"p-�!�e~
]�i�G*�,]��dg�uخ2^+�@"ǶR4y�=��t��d���C*ˤ��U���Xɝ7޶��z&�w�wX�mh��0������7��l��š��f�<�R3pܒ�Hle�6H���*T;=��)Hf�4$-q��������ɼ>}�v0^��	/aV���TɾM4�Jk�����iL����_�MV���%.�$�z���6j��?צj���R9=M.d�}�3�jyG��{���PJ7�O^Z�����������G��Аq�b[�.��ӟ�@��1�ӽա�˨C4���Yu���8�)��E^�r���P�3�I��:�c��p8T�՗����(͔:�C�_`C��
�}L��[R�+͵z����ê�U�r�J����}�
��	�� �X�������:C�����b�Jl���[��\�70���%e|��yVb����EW��S��� ѲĝER�|9t`y]0h��1sQ�U�El�xj4~�&/�'�(I���ő�	��.��-S`"~`��X�rW�.oU�3d>�[����D�i~�'��<��
F8h�ڕ���"���Z~�bGnD%�/�^�OAg��UV��`�k��"|�r�xk+�IR�t.��H7̜�w���a��/��
�Фw9���X�5w,�O�mF���N;��e��'��Z8O4���3�7������oz��Qc�{������6hվx3q��M�t��!'�p�m.rR�!�t(���p�N%=[ٹ���*+}'-G�m��E�?FnWy��ڌ�Ds��⽪�"�w��ݻ�E~[-���8ottG�e)#�ޛ	׸�}���c�}u���a�Hht�Y�g�祆�ڏp秞��~H���χ�"��#�K4ɲ������هɞ[Z����Ơtڌ�,+sE��>�
f��Ga�	sWN����_���G:�ꚯ�t-
�#-ʈL�j�#W���'�d��ؼ����TdX�ާ�� ���w�i�׏2�!����o��ߝіXz9E̟���].���{�F@@�aX�ӥf�ϣW�5jB�9|��q|y"E��t���/��Fb29�R��H���MP�kѣZQ�l�V:���Ga��R���J��J�f�~ܽ2kc5{:~��g�26�>�X��Kk�x�����hfA&�]�E6NER��E�s˛2�i���p�?�,�NxE���Ęz�k���"Q�@d�M�+[[�\�qw���R/�����P{)�蓰�A�i�����#~���|��lQ����6��%�S���0sfX���������$����n<�ݻF��j� :Q��Q正/a���)
_����4��j�]���4\/����:�IA�}��(\΋bbFe?�Zg_
�0�J=7�4�����	`l�}0	�9��FP��|���X[��,��+>:KC��ۣ��U���IŤ�Jm�����^�ԗ$���x�HY�v���3�*�u
��W"��^�����S���ƩI�$Mm>E��1��ç$�5�"V �G�?`f��'��S���G�ؗ	�,;l>��J�������>�u �`��x�F/�٠;)D\�Kt#q�F�bhFl�%t�������ퟕ"�����n�x�����sn�뱸ё2�� ���/Jz�	��8[��,�]cZ�P�[��L<|RK7(}��Y^���/�6�OP<�p�^���^�t��p�W6�b 0I.qs=n*��4�W�`
c|��]���~ 4��unF`�$�r���ͻ4_����^88X�k���!��F��.X�gM�T����<-2C�Z��)����g���2�}��[6��b�Эjwƛt�"l|���De��@=kʼ��^�AW�5��I۔~y���ԭ��+�������?��.-3l�;��_�Q�p~+���\�\��Y��T�+]�?��`�~�,�8��l�9��Mr>��S$�u⍈�d��{��'j;�s��_����� ���,���x���H���0�H=o:�s2���z�a��Q��%5{f7��������~�����k5%��I��h��S�>'�'Qd��'?׺����u[4����A@Q�c<��A�H�n��q*�)��a�K��|�n���r)���W�K���M�&�#ѿ���T�i,�6���JJS���i�)�q7a�OU�@|F�����ͱ.�%��W�'�.��t_���g��E�|��Z�x>:m=��Ů�f�S�ox4�71B�䯌���X�^��wߕ�qj_>�����O���gܣ)�#E����z��'����m��^G�!�٣�ޠw�*�Wd�U����F��w:�Je�JR��=�&u>9�0�*��V�!�3;T*%J��_���զc)��y�#YTe�s{f���r͈0`� ��[�S���6k�fQw0�^��|-���@>~-�=7��6^��2�#�T�������J�"U�Ћ�ގ�Fs�Fg�U�����9��c���f`L��/&#��jqn���Uc鐃/v򙞨y�E��j��^7���l��������E7j�k��s��#���'�m�&�U�[O=
p=GqU���N����KNy��n�#AX0����h����<�Li�P�GP��[�?_��mW�y�i�NZ���N�i|���*�E>�xn�V"{4:�IM"㌺��iv���C����^�f��$QU��v���}m��Ǝ�"I�V ���鸚e��ǟ)��z������my&������F�['����Y�1Z�F�6���k=�o|�DG�[��oz{��ة_���qa��+��S�"�GM�^ݙX�ǟ��˹g,���n?��s���¾���9��Jc0�H�Z��(C-���Q�2z����zF�֌�[��U������#�o��~%��5�)�f��-�V�_@[��"�WV�!�	 ��[R[+��v:���F+x��n��ݣr��a�q�+"W7�3��	)���U��1p鏽�cw��S^a*=�A�0ǟ�{���!��:���Cq�s$[[t����u
�`�J�����_�P�M�����0s���UDl���F���Q��;L	9�焤M�<Ɋ�+S�?��J��e�_N�m��4�-qN������甔2�bT��ne�8�H���n��a�gk3��S�\�^޵b�I�)��)��JU�}���\�(�����o�k,��<��A�H��1ǙI=є�\�{q�D����Z�x�F�����-Dl fZ�$sJ=
K)�t�	�۫�h�hj�"�����
�/�ˬ"��T���!%��T�w�7qaF�T9�1���F�׶l��Ȱ�}�s����lϑ^�T���뿉�2���"�>�|��)1���P�G�*B!�<5�3B�����4��j�܂y:*{S�tgqq�l�Y�v�a�߱\ӯl�o�/�q��}7����hyٟ0e��]N�d\oOm�˱׊��o�f�A?��}A��A��<��t�m,�)&��lE�a�O��4�
�io��ǝ�Z��I�Ml��󧓝Iɸ[�L.�QIO� �bRꜢ�i�%etU��q}_�G�����6��Qo��}���"7�)L��.�E�K�����\�{���G�����H1��H3�0��\c��$4f[�\�f�[;�3B�ݤϣ-u|ͺg`��g���a�v����C�ÄTݳ*�v�z�e��c"��c);��'�:�,�6y����Q���}WD���0�&�@�8���M@?�O+�=7!����=x�t�ۣ랁�׻�EV�5��Z���S�Q{����O���b�5��ghK7��n����ٌ��6�s X�S0���x�%ԴM��Y��>��'u�?��pMɓD��j���e5؂a�;̗��#FzR�A������@��"����%�d7"Q�3cG�D���vޚ≅�֏e>���ͼ��(h>�sB�K]�k�ʹ�N	����K�8Q(;n�B���'���V,���Ô���f+<h"�\K�;��!S�+�Thȱ��2��m��"��3>��JcL����=�%�G/�q-ZT�Q\�M�nn���II�@��I��Ι
��X�V���X].q�5��)�zy� DJ~����5�Zd�ӥ���z����L�>��3����-�H�ӱ�8ګ&��i����Qs��`B�o͊��]-����X�7��q<��1V؎��@L����]�e����JD�8[3ߗ�l^����֚���ŏ��u-/��֦k�e`2;�~N�ܼ�T��-�S�JFW��Z�W|-�7�z�t�>��.�� s��	�ʥ?X�i��w"��s�En�.� �����:oM\�A�a}��:�uُ��7ka$�_y�K�>�������v���d��ٚ�=��Uą�r��/C�hQP�$�t?	�[�u�r��7��y��o�8frufh���1�C^�L+���ð�԰��p+�VmH���G��# ,n��V
�9O��!���Z�)�����Z1�K�< �p+��'A�Y��GJ>�ux��|�U/p���Ǡ��sSO�5`m�@5���]�sK{�:	�Ի������,X���q�
�hiO�����I������_��O��\�[C�|�t,N�T��]�d�K���>f8P�4zS���|J�?��,N�,�t��lw��M�DY�����Z��G��L��|��T�q�B��\��P�<��P� z9y�>\�I��6?5���mc<�!�t��(���Ϣ6��{IDz�|�-��~������
�.��dw�"��]�L�k ��m[j����,�V�>��i�����ё�ڝq]y��A�)�,/L�Dx��l�������u�:��͘4�8Z�)^TX$��bU$��aͲ7ER.mZ��}�=����/T�c1x�	e���!S�����?
+~w����,%����FB�v��c����Rn�zW8���7N��A�����X��*XWa�A��E���J|Dr0Y�ֺ�[�k�;��JXï{zy>?��eX���a�U���-@Zh��i��ý �/�w��o^��Z�	�9�F������{����Gz�'{�j�B9�~�OSKߦ>��S�3H�/��+�,�r��jM���s5�1��� ���%�}��A
�A+��JuhHle���Ls��`@�����B����Q$�+������"����e��Ǡ��D݉�k�1wa�Ӄ��	�/!�6?��!JOE�d���y~��d��ȵΘ��OYd"������Zez~(�� ���M�z,��d��l2��e�7^J4����i���^V����#�A5�%��\bBf��MGk��];��~BNW�!�٪�E����!��z����`�}h�˗_�`g��=�r������$�+�%�"��K���*����o���O��lY�i�cڄ���������Ș 	�]%�ѓX�+����yM�͇���:��AnP%]��7`AE�+l��S/:l4��P�
rK��b��Y�"bbc��~�0�HOb�H���k�������9s`��{^;��ĕt�������Pb���Z	��	�����i<o����.+�Yƨ㤋@h�&�)���E�t(3��\�|�͡/O�7�N���v�	��0@�L�߭) �ۄ>�㌰���C���1{���s���|�������>Tg`.��p"�Tm� l�E'��$Q����A2��3q��0�ݚ��ϱ�)%��(�5/O4��$�$N}JT��/M�e�~�W �P ������ݖ��*�r',,��M�����rP�oɯ�X��I:?dyT��~�1�@�HJw4�|��7h����g�1���p(��<e���w��?-zF�		L�u>�Pj�V�h�m��=\�Eď����Nк��(s�v[x6_s�� sauּw|�=u���.�����ײ��~�j7�@����R-�9��h�=�Gs��y��,|���3x0��)w�p��^}�<��ڂĝ�{/�����\�
V��<�T$ę3A��+q�R7t�u�`-6�"�s^�k�x��J{��]�T὇nA��$KF�=�K�gP[����A�<	�7�7!~�\���^F��m���,�����`jw��֌����j	�A�[ ��r��)�@�vjͤF��{۽�k$\��r�O�u���#����`E9�	���@>Z�4�jʳ��#�,��,�gl�ea�jY )W���6�I��{[ �%���	c�����S�_���w�@�hlB�� �M������������Ĳ�As��bar�}�u~
}�U����__��P�$*��}.��L�H[ۉSiC��=��������?�:a��(p�F�9�l��W,�׿y#�I��]�����A
^��d` �OÎ�-�X΂�[����g�?��5	9v�b�s@7\��7^�|dgNt�@jx���r�V�6�gl�l��T톅��ޮ}(���� ��W0+b�1˄����d��믙ʞ��?�
S?b72��um��t��".�	�c�o�����k��w�]#���������}�Z@���ej;(F�}5�1I@"�FJ��l�2��.G=�:~Lu�ujzON�%�#?X�T�2��W~v�=�����+M=�w��_-AX%Ky{�#"�m�ߖ��R�-�Ip��?ů�x����?�^a�Iq��1�Y�����R�_�>{���0:���mU�ꚩ�/���E�!~�Հ`d�ר{�mPF�;U��/�rX��{!�O�)i�ٮ��]��?�Db�e������_��ɚ�X��}����o�
��"ܸC���z7��Y��a���I��m�g��f���u��Sܾ����c�+��1h�Ǡ�D
����V�&|B�J$�g���6̍�n����\��ϊ~����&_��Ő�-�|r����W������6�����Gy����X}>��R�o�K�Gz�)SuSjM�٬�t
� ���&��G}v��ޔ[�|1C>��#:�Z1�Yj��B���ҹeS�[+��&*xqԓ�2��ߨFE�b�#Zy�M7��zA�C��y`2��b�@N����j�VYM����dߋ�;�]�jUB�������u����A,/�*�W�2`��BO�h���&lT���J�פxB�>DZX��eg��'	�O
����/�`�>{��L��;�if���f��wJ�P��q�b���P�Ǉ�(�~��qΥ�ΒQ.�]�����6��}?�vq�M~h��gN@�\;E��c����W�F�&_�c/��5m��>!S����
 N�2����3X�eq�e�}N E�֢�:*�N�����Zr����U  K��{ /v4��g���E4r�G�5ʰ�/P&=�L@�@���vR��SW[-��<"�#�˩oj�-����L���=tA*�,k����&e��J�I�a�d��,y�����"��DBʑW�]	ou'�e�����j&h���}Jj���U��U���ˊ�*��(�1UU6kXB#|@�_����
6�9lrڏ9[{�p���� ��?�S[��j#����q�B�LDA+�V�h�eh�[n�x�E\3sY��f�w�.�Z������<��mmx�_Ξv�ltX�>A�O�n�@��OF��|\�k@��V���� 
�cWsx9�)�x������a�9HhX��6�~N�l�1�lk c�TC� �u-ͷ�_͌{�'m���LP��s��H-D݀BCXcJ�[g3EnFp^Jٸ{�#�l7v�D9���55N-I��ak�7y��/��`'�� "cQX[|,;p���2y���H(\�ZY�N�|��Ծ��jNʁ�
 � Ҵ��׆@�0�dN��Ʋ�ݚ+�+�,������(?�iZM�&.����SL��V���$*pc��#�ru_T�@~�}1N�����lx�����j&L�=?G^�~�ޑ� �r�*�Ѥ ��&�5bd���Q1����CF��2Ƣ���ܷI����4��/��%0ғI�hf�f�]�P������ޛgǬ�5�De=��� �$�n�w�i�/m�{�	�"/��l�P��ch ύ�u�BR����9�?�)y��z�.g�U(9�̏����%���Bd��M��(.��2���	�d_�M�u�IAl��M��S7��"އE��W����xb-dϗ�K8�����i��1�%۝���{t3_�ɓSK	�*���v���l�7��E;���0��';|��/=P)��O��z� i��E)V-�Ni���]g曂���Ř���f|ǽa�a����8�Dkw��J�9�_{7�����s�B�ӊ���n�=�;�+P�D�B�='��O�[��m��
���U�س��F�5�)Q��vG�,�w>�&���E�m���:�~�`�|�H&��7�Y\'����e�S�C��i��6lɃ���؏{��*+�J�7�p��R>��� �i_v�M��H�V �H~s���T��C��Fnp ��.�R 4���o :�g�y�U8�B��'��:bJb
=���uv�Gz���V�w���oH�ѥ&��/Sz���Ʈ�k�(�Q���j�J@��S�;sЫ!3?~Aѵ���{u���3����S4�a�,ր�z�=��%}��h�J�N׀8ݿ�}���c�t~@�:�f-�X����}7��D!�����.c��A�:u2��ֻk��M�\4�_0g�<+�!5��/��?�0#~�)�$f)<�"4up{M>�2�u�,+�Ɓ!�HVI�����e�$cr�d�.
�N�?��)��Sg�&3�[�����/�� i@2�KP\2E��q4�����܈�Iz��X��}#G�Je�G�l=N�Gv;�Ԭc���j^F7q���l:q*p��PΥ��ٗ�W�}E<��z��5~PȨ�Ȗ_V�R��W�{��C��8�R>�8�[9�2���x&`��H�ߘ��>H�"�=o�G��[뛽d����⾈��H��IE�FC=�PF�-��+����6w���L�ٸ����0"��o��?2��㇘6��&�آr{ w��H�xWId�]��o���#���lS��	u�\A�|͝�$HD���5ښdӖ���2nG��'Y�ł�b$`��n���j��ec��e��ۡ<�͇%r0Y���%U�Z��W7(w�Wu�ρ@��f�̑�w����e߭f&��b�4ɒa�K���'TzVh�Oiyq���W�|�%:�9k	�{����rl��)_�� ��K�t8�� ȍ���~N��䔷�=|�k�@�>QX���#d;���K��A_�nG�@�Av�^af]��z�;婚Sn�Fj��b@�r`#�+P�$ov����&ʂ%2�Up*��S;��D�ܚ����a�T�%L0�4��<�!S�4�[��z6��w�����ƞ<^�X�e�8��E����箛y��e�D�Ub)�_H?
��"��k��E�~E��ɯ�a{�
f*�hH���&l� n+(B#��:�r����z���&�������O�a�X�$�����)�SyOKs�'��z���`�B�b;*�4�O3�B[��\�*�?����Y�
r58�\ <H�cLl�y�+}.��8Q�Wk�O
���'M�X���%{�~����9��t1��m�(�UayW3�t��zƆ���7�5��Crd۷;�a�h�?� �ТN��K�,a�,�e�lr����#>�r��v��1��TǬ~��6�d���1D��`�:k�s
&w��h|I�c��ډ�ou_V@�A*u
%��
�T!��u>���!�<pa}���	���Os�����p��^<e|٣�K?,xv0ED"l
�����*��I��	},E
)�Gj�<k���jcLۂ���ϵ��qr>�au�i�U������ɋN��l��/-��VZ�Ë�e�K�2/�^�
��î�?@��=#t�#�P�n(��Rx��\3�[܀ճJx��v��y@#��q��[��z�������[> �}O��(>*y<o����{��h�J'��w3io59bl�_�t�?�1I�P��W�|���E_&�9�����)�w�r'쁡����;�`N�|���]z�L.�2q�(��2��-���.p�V���d��B�s���'���)��uOsA��F�w�l�;#c�R�Q��b�ؽ-���R�qe6}�xo�G���C�31��^�;DJ�����]�=(�]t��ܮ�ق��qX����IO��6��B>)����T�_6q0�i$�`��40�<h�2;�;C1	4_�(�%vK[��	�����j���P�����j7�䙫q2��tM�~|�������M��@�2��'m+*�c#��8N�>��[�t��W�=x��c�FP 7�M{ ���6堇_�4��H�
�x�ޱ~�2�r�'�]f5A���ݸ{�Q��a�e��ӓ��~?5 3��Q:EA%��?�d��������I9R�W��)�<���)��a�z?8���d��!iu�`��&�\(��0Ƚ�A0��x��)���aK�ۘ46Mq^;�QQ7Ik�j�N�jSӉ�&�>,`�Է�f�y>׶�p[=0c�s� =8�)�cb1��WᏢ�"j�D����u��)A3�놂����+g}�?���<�����a��أLeTY� m����xPΐ6!U聄M���6ԯs%`�����ϥ�}���Z���	�2iN>�?1�׫6�|=p�ѝ�8���w-��X�����T20Q�Ҷ��g蚴�,�uc-��g��/9��=�D��ͯ1[)��>��}��|f�b�$a��|���u9�#ǍT:C ';�����4�<��1�3���3V�_���Gm%'*����M����#/�-��&��④ �Y88��U�|�.�JK��X�	$W��Y��bD������Rk�-I`nX �](�1

���e)�;�"����[fH����>#p�Y�%*�C*=I"�7���iѱ����h��jļ���N�Ճ:�mٸA�t��u��kRה BT�^NMB���5v�/��R��V��iQ7�r��T�0�`+���V��&�����aw�>)����5	�4�C�<	z��o�.C�@#��#[�Vd�1����%b����9`R���u�ֵ96��C27���E9r�)g�����u�x�̸؉���O��`p_�m�j�-y���9��L�l����M|K��2F���>O�X��4p���rj��Q�Pcv&dֽ]�����v�<��w�Pm�������=n�/�z�J�Ld3�ŗ���� FZ���s���x-:e�����H�{J8��V*�D�r0n�1�S�o0��l�H} ��Z莸W� �	1���x�鰪5~Ko�W>NdO�,�F��U�=���g��Y���3�K)���,���F/�zH��K����&�f��l�R��ۯ�ݶ:����೶󯧂
��E�5S��OB���/�
��1���?�\����gP��� �2ͯr �| Q�v�Bכ߇v� Q%�F`��Z�|\ˌ s`�5�&����po�	,��& �T
Z�S�-����\�'�Z-�Y@���T�	9p��5x9J�_�����-��X����[�˭��y��M�[�G!��޼�K�_�}�=�wrc�K�g���!)��y�����U�r7�4%ÁB_�w[�ۯ��+�(u#V;��C�,f�:�-�=8�N\�f���'<K����ɋ�\ F�V����}k�I�鿀�������tpZ��u;rx-�A��[ L^��2A�mq���^�R���2P��Z�������m���_N������V[޿z������:������I����������{>�]�	�g{�7N��{;���V���h����׶�kÖ���_�r~a\��3ooo����c%O�;:����)�2��.�����Ӟ��o.�� �F��W����0)xs�y����>��q\_G�&�������u�����U+lǸ����������k�����ɷ����G��^NWR�w��GƧ�g��vT��Vi(�z�a���?��*�ς��"N��� /�>�ܟ2���!h����4�ݏ!�����D���__[��5�����Щo�����+h����Z�P��n����O� 4��|}}|������,�d*gh����-S.`�|�P95�
.u�!�e���� _��+��w@��Т�%;� � *e`�*���+h��f�Y
p�d��6Z7 m�뛉ۨ�W��~�04�Ad/~t��y�A�������P
�m,�K %�z;�g������ɐ�
�H3�����=������7+�}�7���l~��ҿ�o;d��f����&�꠵ &\�J�V��m;�AW�dg��&��\��+��c���lp8^ �A���ա���W���A�3N�C�"(��^�o�+��(�d�!2C�l���F���!a|�Q��R��峺�xKb0��!2J��<�S�4;����'#�g��-���1T�TU�"� �;ȁ����"`�?u�NX�7\nm�����H�"dxQ��������2:�>����w+	M�jk݀Z-�F�ϊb�jr�N�	�;��ӡL�`y'*ѦL�3!�	��m|������@�%�������7d��I��'����u�&�\~���>�f`aJ�wr�-5������	Vu� +��L�_}r�x�l����=� b8\����@;g��a�3�H�[�<������)�	 PK   �i;YB4��  �_     jsons/user_defined.json�\[o��+��"���/~S��pˮ�:
#���D(R�EN��쒒,��p(	-�R/&�����9߹��x��U���q�c��d��h|��|�7�,׮��r��_�ݼ9��ݽǋ������Q!1|��U�8_�
_������g��|:���^��V���N��h<��c�M+���Ȑ� �Z�|�m�#�n5�q����f�w��N<����C"*��&9��10i�Z��j��kv��<�K{�xy	O�\Mf�f�|���l}y:Y^M�'�)lĘ�F�W�?w�)�ܸ٬�l���4{ޭ���}a��t+=���>"��`�<��O��2~�Z�ao����[�ޜ�����4*��4�v��`�VT���,,��*X��eA�TU���YL1��U�=;͂�!�y2��R\���YTAi�1�b�!f��b���IE�����A���u��7R2d�3�c��֙��ȃ�D�l�X�A���u���CB1R��CB�J�7y�!�X���E��b��O�CN�J�'yR�!�X���<��U�� $O+:��d ��y�� �;aO)y���<��]�ʪ��w��y��x%41/�(Z�i�Z��(A'�Fk������a�cN������ �ĵ�V�'K�6S�a��D�S��xt�C�ϱD��e]�����8��ȉ�W�VF2��҆���d-kD9�P�F��ie-WT�'
6m�u9Q��JdSFN�m���2t�v�Ф���x-t��<QȱZ�2y���uХz�IHH�q���C
\�[������ЈD��{�֊Dڡ�
����"��v��5�D"�Pe���7"��v��5_܉D�١�
�|.�g�j*P�J$��Bt7lA]�����]3�����fK+`�
�z���:ey���H�X^e2C0R�0�W��0�TP��U&3#��e8F*HF*ː�T��T�aYEX(4e�d?9*�!�zԚ����Ԑb=jMT�׵jȰ�&*�SjH��&*�sjȯ�&*�(jH��&*�5dǵQ���!�6�5Q���!�6�5Q������BAc~UE���t�`UQ!�2�aXUTȫLg(V�*��UE���t�dUQ����*�~�z�^�,b I���*.V��z;�^nd�g�y����\�麟^�@��(X�j�#�~3;�_^�
�&��'ˉ���k����Oi�'�I��uk�j���/Eo��� �c������7aBZ�m Ȇ�"�c�ͬ�ν=ș��l��f�O ��~��ͽ��է�r����S��y���QFF�'��c�²G7C���>�aj�ƈ{��: b�ǭ�u�6��{�6s�s ؆@�(H�#�}��U��Y��v?�6�KB0E	���䌓Hν�*Mnn*�W� �Ѵw3�C���lJ��NH�P�(?��5��>S*�)`��{�(�E�������~��Rm�yn�{t����sT���yx*e����=������n���0�����y�qr�{���v�Җ;��!�Ң�H�F�&4<7���F84�x���i���.ʨ�V���K��$q���+�̳V&���k"y_Tx��g{��_�1%�Hi�h��&V�ڧ�y�M4��Ȝ�=8�� *<�����>�dg�8[�2�V�sPB�}h��#)o����s� .���el����u!\�r`�A	��s�<QMvQ��Z��
��Ɇ,qC%�O,O�����G2�4�1E�L�d���`ȥ�=1ŔL5Z!<������	��� y(@	v�hWgi�"�v(�x�`��|+@(b�N����F�F1F`�i��C����f ��x�*$њ��4S�@ �T#��CY@���:@U#Io�����Y�<
 ��`�:0����'�7�a�pc�� @4<�.+*���;J� �6��}��$�mX��R�N k8�j�
��|<��v�3�D�]fz�f�3x�{ H0L' t`�ޥ��%�����X?��f�P�(a�����(1*��"�	B44��	�MJLM��l )Ԫ^BA@�1|�G(lR�$�](�]u�������8�G%� �M�h���-)qȏj���{K�}��&����H�u��QJ�'XR��ǸakzK��]�  uR�u�S!@��N�QؤԬ��F���XR��M p
{ө�4�r�MJ��� T,��Bi��n	,V�;KҴ�Z�]�Ji���.Ǔ�n6��V���Z����J-6)q\�wY$7{���CBIpj���C>ͺ��3������cKҷ��'�^����+���]ϊ?���E��C�р�����Ԗ��<��9�b��(Ql�C<*�4��|���q[>�
D�tT�d}(:�m|��}p�@�ђ�?��K��/8
�� ١�N�>�!�4	� H���P8N����D���%�眛�=�@�[��09����z���N��V8���+�C���j��cF��N��`)-TQ)U��lQ�EZ�`�B��Zo@��X{x�H4☀7��"è��dc9x��7����I���z��:�l<"��rXE�,y>o�P�.F���ռj�B�6�K���A�*�]i�4�VX�����7�x�삌-␴"mZ�L�R�X<4���D	摆{7��Ҙ��-��?�2MUX�����E4D��$�w��b�fG�2JI�](������`��ޢ�&��:����u0��q��`\�:������E���k�Z�Eձ�(5o�Hh�7xr��ȷ�����Gk���d�#�<J���`]��qZ�5I-�sD.*0���$D4�P����7ݩo�4����4,�u#���H�h!�`Rq߲���T7TfJ����W�5����%�����.AA��$�J�(����t͐$���)Iq[ې4�Z�C1*��f�4���.�ֻV�!ِ|��l���]LV���m����v-��V�݆�t�V�����9�׀��t���&���kDe�[���ŕ��n�Ş�}��q;�\�ܰ�������ۍ�o�b	w���?}\�׳ ��]�ӷ�_�3� �\Y�ȞP�nV�oX�T;���M��X~�9���g�si1���I�(�`�<��x:�9x���τ��X�����@�X,�t�7��r�.ְ�����YƑ�N#l����"�U�>ž���X㥢Ha�A��7aj�$x������q�X7���o�~KzRp��ϓ����/�HN�_���x����x ��E.f�ٮ����z$��m�,
�Sh��h����#	������X[�^�º���,ӄg��!�;�z�T��R�C��#T�|���X>��?PK   �i;Y�K�e�5  E�            ��    cirkitFile.jsonPK   �i;Y��(� � /           ���5  images/0add2520-d67e-4490-80cf-da78ad043e6f.pngPK   �i;Y�R�� $� /           ���Q images/179c08ce-6e18-4019-8002-932a24469ad1.pngPK   �i;Y=���C; �; /           ��2) images/21a1dd99-e68d-47c5-b9b6-5144ca492781.pngPK   �i;Y����7  �  /           ���d images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   �i;YF@vw'� � /           ��Fv images/36b3ed9c-16ef-4839-89fb-9e068aa5b597.pngPK   �i;Y'(�5W �@ /           ���. images/4737cce6-ef6b-4e79-82eb-dab57378d86e.pngPK   �i;Yh`Pҷ!  �!  /           ��^K images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.pngPK   �i;Ym_D�� �� /           ��bm images/51bdce1f-f35a-4993-9bab-5f201461b496.pngPK   �i;YM�f�  �  /           ��p= images/54318eec-5d24-4037-8f7a-d01382cfeac9.pngPK   �i;Y��N  +Q  /           ���F images/55dfa5c9-aad1-4e65-bbd0-3dabf009b856.pngPK   �i;Y/��<  �>  /           ���� images/686a6ed9-be7d-4d85-81e9-18457125bd85.pngPK   �i;Y5��s� � /           ���� images/7b4f3c61-861a-43c5-a680-e3c3f7136b2c.pngPK   �i;Y�IM��  � /           ����! images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK   �i;Y�&�}[  y`  /           ��N�" images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   �i;Y�i{J�� � /           ��+# images/bbc1753c-83ed-490f-889e-b8df35028df1.pngPK   �i;Yp>r�  �  /           ��B* images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK   �i;Y�ɯP� ȉ /           ��{0* images/d509810e-83a7-410e-8a4f-883955ebe6e7.pngPK   �i;Y��<���
 ��
 /           ����, images/d75681bb-bbce-4690-8af0-fbed32c25461.pngPK   �i;YF��-$  ($  /           ���w7 images/d88a5b0e-66b3-4edb-b452-47f46dd40326.pngPK   �i;Y�H�izN  �g  /           ���7 images/e9a9c672-7031-4851-9c94-029b4a1edcac.pngPK   �i;YB4��  �_             ����7 jsons/user_defined.jsonPK      �  ��7   